module real_aes_2444_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g192 ( .A(n_0), .B(n_139), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_1), .B(n_769), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_2), .B(n_123), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_3), .B(n_141), .Y(n_520) );
INVx1_ASAP7_75t_L g130 ( .A(n_4), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_5), .B(n_123), .Y(n_122) );
NAND2xp33_ASAP7_75t_SL g236 ( .A(n_6), .B(n_129), .Y(n_236) );
INVx1_ASAP7_75t_L g228 ( .A(n_7), .Y(n_228) );
CKINVDCx16_ASAP7_75t_R g769 ( .A(n_8), .Y(n_769) );
AND2x2_ASAP7_75t_L g117 ( .A(n_9), .B(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g458 ( .A(n_10), .B(n_234), .Y(n_458) );
AND2x2_ASAP7_75t_L g522 ( .A(n_11), .B(n_168), .Y(n_522) );
INVx2_ASAP7_75t_L g119 ( .A(n_12), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_13), .B(n_141), .Y(n_504) );
CKINVDCx16_ASAP7_75t_R g429 ( .A(n_14), .Y(n_429) );
AOI221x1_ASAP7_75t_L g231 ( .A1(n_15), .A2(n_132), .B1(n_232), .B2(n_234), .C(n_235), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_16), .B(n_123), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_17), .B(n_123), .Y(n_477) );
INVx1_ASAP7_75t_L g432 ( .A(n_18), .Y(n_432) );
OAI22xp33_ASAP7_75t_L g760 ( .A1(n_19), .A2(n_110), .B1(n_111), .B2(n_761), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_19), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_20), .A2(n_88), .B1(n_123), .B2(n_172), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_21), .A2(n_132), .B(n_137), .Y(n_131) );
AOI221xp5_ASAP7_75t_SL g202 ( .A1(n_22), .A2(n_35), .B1(n_123), .B2(n_132), .C(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_23), .B(n_139), .Y(n_138) );
OR2x2_ASAP7_75t_L g120 ( .A(n_24), .B(n_87), .Y(n_120) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_24), .A2(n_87), .B(n_119), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_25), .B(n_141), .Y(n_219) );
INVxp67_ASAP7_75t_L g230 ( .A(n_26), .Y(n_230) );
AND2x2_ASAP7_75t_L g163 ( .A(n_27), .B(n_153), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_28), .A2(n_132), .B(n_191), .Y(n_190) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_29), .A2(n_234), .B(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_30), .B(n_141), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_31), .A2(n_132), .B(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_32), .B(n_141), .Y(n_493) );
AND2x2_ASAP7_75t_L g129 ( .A(n_33), .B(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g133 ( .A(n_33), .B(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g180 ( .A(n_33), .Y(n_180) );
OR2x6_ASAP7_75t_L g430 ( .A(n_34), .B(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_36), .B(n_123), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_37), .A2(n_79), .B1(n_132), .B2(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_38), .B(n_141), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_39), .B(n_123), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_40), .B(n_139), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_41), .A2(n_132), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g107 ( .A(n_42), .Y(n_107) );
AND2x2_ASAP7_75t_L g195 ( .A(n_43), .B(n_153), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_44), .B(n_139), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_45), .B(n_153), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_46), .B(n_123), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_47), .Y(n_752) );
INVx1_ASAP7_75t_L g126 ( .A(n_48), .Y(n_126) );
INVx1_ASAP7_75t_L g136 ( .A(n_48), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_49), .B(n_141), .Y(n_456) );
AND2x2_ASAP7_75t_L g468 ( .A(n_50), .B(n_153), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_51), .B(n_123), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_52), .B(n_139), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_53), .B(n_139), .Y(n_492) );
AND2x2_ASAP7_75t_L g154 ( .A(n_54), .B(n_153), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_55), .B(n_123), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_56), .B(n_141), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_57), .B(n_123), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_58), .A2(n_132), .B(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_59), .B(n_139), .Y(n_150) );
AND2x2_ASAP7_75t_SL g220 ( .A(n_60), .B(n_118), .Y(n_220) );
AND2x2_ASAP7_75t_L g483 ( .A(n_61), .B(n_118), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_62), .A2(n_132), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_63), .B(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_SL g183 ( .A(n_64), .B(n_168), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_65), .B(n_139), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_66), .B(n_139), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_67), .A2(n_90), .B1(n_132), .B2(n_178), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_68), .B(n_141), .Y(n_480) );
INVx1_ASAP7_75t_L g128 ( .A(n_69), .Y(n_128) );
INVx1_ASAP7_75t_L g134 ( .A(n_69), .Y(n_134) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_70), .A2(n_100), .B1(n_762), .B2(n_770), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_71), .B(n_139), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_72), .A2(n_132), .B(n_472), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_73), .A2(n_132), .B(n_446), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_74), .A2(n_132), .B(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g495 ( .A(n_75), .B(n_118), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_76), .B(n_153), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_77), .B(n_123), .Y(n_151) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_78), .A2(n_81), .B1(n_123), .B2(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g433 ( .A(n_80), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_82), .B(n_139), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_83), .B(n_139), .Y(n_205) );
AND2x2_ASAP7_75t_L g449 ( .A(n_84), .B(n_168), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_85), .A2(n_107), .B1(n_745), .B2(n_747), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_86), .A2(n_132), .B(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_89), .B(n_141), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_91), .A2(n_132), .B(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_92), .B(n_141), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_93), .B(n_123), .Y(n_194) );
INVxp67_ASAP7_75t_L g233 ( .A(n_94), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_95), .B(n_141), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_96), .A2(n_132), .B(n_217), .Y(n_216) );
BUFx2_ASAP7_75t_L g482 ( .A(n_97), .Y(n_482) );
BUFx2_ASAP7_75t_SL g105 ( .A(n_98), .Y(n_105) );
AO21x2_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_106), .B(n_758), .Y(n_100) );
INVx1_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_103), .B(n_759), .Y(n_758) );
CKINVDCx11_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
CKINVDCx8_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
OAI211xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_108), .B(n_744), .C(n_750), .Y(n_106) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OAI22x1_ASAP7_75t_SL g109 ( .A1(n_110), .A2(n_427), .B1(n_434), .B2(n_740), .Y(n_109) );
INVx3_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OAI22xp5_ASAP7_75t_SL g747 ( .A1(n_111), .A2(n_435), .B1(n_748), .B2(n_749), .Y(n_747) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_357), .Y(n_111) );
NOR4xp25_ASAP7_75t_SL g112 ( .A(n_113), .B(n_250), .C(n_294), .D(n_321), .Y(n_112) );
OAI221xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_211), .B1(n_221), .B2(n_238), .C(n_240), .Y(n_113) );
AOI32xp33_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_164), .A3(n_184), .B1(n_196), .B2(n_207), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_115), .B(n_393), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_115), .A2(n_363), .B1(n_421), .B2(n_424), .Y(n_420) );
AND2x4_ASAP7_75t_SL g115 ( .A(n_116), .B(n_144), .Y(n_115) );
INVx5_ASAP7_75t_L g210 ( .A(n_116), .Y(n_210) );
OR2x2_ASAP7_75t_L g239 ( .A(n_116), .B(n_209), .Y(n_239) );
AND2x4_ASAP7_75t_L g241 ( .A(n_116), .B(n_156), .Y(n_241) );
INVx2_ASAP7_75t_L g256 ( .A(n_116), .Y(n_256) );
OR2x2_ASAP7_75t_L g268 ( .A(n_116), .B(n_165), .Y(n_268) );
AND2x2_ASAP7_75t_L g275 ( .A(n_116), .B(n_155), .Y(n_275) );
AND2x2_ASAP7_75t_SL g317 ( .A(n_116), .B(n_198), .Y(n_317) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_116), .Y(n_374) );
OR2x6_ASAP7_75t_L g116 ( .A(n_117), .B(n_121), .Y(n_116) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_118), .Y(n_153) );
AND2x2_ASAP7_75t_SL g118 ( .A(n_119), .B(n_120), .Y(n_118) );
AND2x4_ASAP7_75t_L g143 ( .A(n_119), .B(n_120), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_131), .B(n_143), .Y(n_121) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_129), .Y(n_123) );
INVx1_ASAP7_75t_L g237 ( .A(n_124), .Y(n_237) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_127), .Y(n_124) );
AND2x6_ASAP7_75t_L g139 ( .A(n_125), .B(n_134), .Y(n_139) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x4_ASAP7_75t_L g141 ( .A(n_127), .B(n_136), .Y(n_141) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx5_ASAP7_75t_L g142 ( .A(n_129), .Y(n_142) );
AND2x2_ASAP7_75t_L g135 ( .A(n_130), .B(n_136), .Y(n_135) );
HB1xp67_ASAP7_75t_L g175 ( .A(n_130), .Y(n_175) );
AND2x6_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
BUFx3_ASAP7_75t_L g176 ( .A(n_133), .Y(n_176) );
INVx2_ASAP7_75t_L g182 ( .A(n_134), .Y(n_182) );
AND2x4_ASAP7_75t_L g178 ( .A(n_135), .B(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g174 ( .A(n_136), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_140), .B(n_142), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_139), .B(n_482), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_142), .A2(n_149), .B(n_150), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_142), .A2(n_160), .B(n_161), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_142), .A2(n_192), .B(n_193), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_142), .A2(n_204), .B(n_205), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_142), .A2(n_218), .B(n_219), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_142), .A2(n_447), .B(n_448), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_142), .A2(n_455), .B(n_456), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_142), .A2(n_473), .B(n_474), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_142), .A2(n_480), .B(n_481), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_142), .A2(n_492), .B(n_493), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_142), .A2(n_504), .B(n_505), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_142), .A2(n_519), .B(n_520), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_143), .B(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_143), .B(n_230), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_143), .B(n_233), .Y(n_232) );
NOR3xp33_ASAP7_75t_L g235 ( .A(n_143), .B(n_236), .C(n_237), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_143), .A2(n_470), .B(n_471), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_143), .A2(n_501), .B(n_502), .Y(n_500) );
INVx3_ASAP7_75t_SL g269 ( .A(n_144), .Y(n_269) );
AND2x2_ASAP7_75t_L g288 ( .A(n_144), .B(n_210), .Y(n_288) );
AOI32xp33_ASAP7_75t_L g403 ( .A1(n_144), .A2(n_274), .A3(n_304), .B1(n_334), .B2(n_369), .Y(n_403) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_155), .Y(n_144) );
AND2x2_ASAP7_75t_L g243 ( .A(n_145), .B(n_165), .Y(n_243) );
OR2x2_ASAP7_75t_L g259 ( .A(n_145), .B(n_156), .Y(n_259) );
INVx1_ASAP7_75t_L g282 ( .A(n_145), .Y(n_282) );
INVx2_ASAP7_75t_L g298 ( .A(n_145), .Y(n_298) );
AND2x2_ASAP7_75t_L g335 ( .A(n_145), .B(n_198), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_145), .B(n_156), .Y(n_354) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_145), .Y(n_423) );
AO21x2_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_152), .B(n_154), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_151), .Y(n_146) );
AO21x2_ASAP7_75t_L g156 ( .A1(n_152), .A2(n_157), .B(n_163), .Y(n_156) );
AO21x2_ASAP7_75t_L g209 ( .A1(n_152), .A2(n_157), .B(n_163), .Y(n_209) );
AOI21x1_ASAP7_75t_L g515 ( .A1(n_152), .A2(n_516), .B(n_522), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_153), .Y(n_152) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_153), .A2(n_202), .B(n_206), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_153), .A2(n_444), .B(n_445), .Y(n_443) );
AO21x2_ASAP7_75t_L g461 ( .A1(n_153), .A2(n_462), .B(n_463), .Y(n_461) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g390 ( .A(n_156), .B(n_165), .Y(n_390) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_156), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_162), .Y(n_157) );
OR2x2_ASAP7_75t_L g238 ( .A(n_164), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g244 ( .A(n_164), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g257 ( .A(n_164), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g419 ( .A(n_164), .B(n_288), .Y(n_419) );
BUFx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g348 ( .A(n_165), .B(n_298), .Y(n_348) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_166), .Y(n_198) );
AOI21x1_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_170), .B(n_183), .Y(n_166) );
INVx2_ASAP7_75t_SL g167 ( .A(n_168), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_168), .A2(n_215), .B(n_216), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_168), .A2(n_477), .B(n_478), .Y(n_476) );
BUFx4f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx3_ASAP7_75t_L g188 ( .A(n_169), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_171), .B(n_177), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_172), .A2(n_178), .B1(n_227), .B2(n_229), .Y(n_226) );
AND2x4_ASAP7_75t_L g172 ( .A(n_173), .B(n_176), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
NOR2x1p5_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
INVx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_184), .B(n_315), .Y(n_417) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_185), .B(n_365), .Y(n_364) );
HB1xp67_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g200 ( .A(n_186), .B(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g222 ( .A(n_186), .Y(n_222) );
AND2x2_ASAP7_75t_L g248 ( .A(n_186), .B(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_186), .B(n_224), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_186), .B(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g306 ( .A(n_186), .Y(n_306) );
OR2x2_ASAP7_75t_L g325 ( .A(n_186), .B(n_252), .Y(n_325) );
INVx1_ASAP7_75t_L g332 ( .A(n_186), .Y(n_332) );
NOR2xp33_ASAP7_75t_R g384 ( .A(n_186), .B(n_213), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_186), .B(n_225), .Y(n_388) );
INVx3_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AOI21x1_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_195), .Y(n_187) );
INVx4_ASAP7_75t_L g234 ( .A(n_188), .Y(n_234) );
AO21x2_ASAP7_75t_L g451 ( .A1(n_188), .A2(n_452), .B(n_458), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_190), .B(n_194), .Y(n_189) );
AOI32xp33_ASAP7_75t_L g411 ( .A1(n_196), .A2(n_247), .A3(n_412), .B1(n_413), .B2(n_414), .Y(n_411) );
INVx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
OR2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
INVx2_ASAP7_75t_L g278 ( .A(n_198), .Y(n_278) );
AND2x4_ASAP7_75t_L g297 ( .A(n_198), .B(n_298), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_198), .B(n_269), .Y(n_326) );
OR2x2_ASAP7_75t_L g380 ( .A(n_198), .B(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g338 ( .A(n_199), .B(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g396 ( .A(n_199), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_200), .B(n_213), .Y(n_362) );
AND2x2_ASAP7_75t_L g399 ( .A(n_200), .B(n_365), .Y(n_399) );
INVx2_ASAP7_75t_L g249 ( .A(n_201), .Y(n_249) );
INVx2_ASAP7_75t_L g252 ( .A(n_201), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_201), .B(n_213), .Y(n_272) );
INVx1_ASAP7_75t_L g303 ( .A(n_201), .Y(n_303) );
OR2x2_ASAP7_75t_L g329 ( .A(n_201), .B(n_213), .Y(n_329) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_201), .Y(n_381) );
BUFx3_ASAP7_75t_L g410 ( .A(n_201), .Y(n_410) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g279 ( .A(n_208), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_208), .B(n_297), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_208), .B(n_368), .Y(n_367) );
AND2x4_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_209), .B(n_282), .Y(n_281) );
OAI21xp33_ASAP7_75t_L g311 ( .A1(n_209), .A2(n_278), .B(n_296), .Y(n_311) );
OAI32xp33_ASAP7_75t_L g333 ( .A1(n_210), .A2(n_334), .A3(n_336), .B1(n_338), .B2(n_340), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_210), .B(n_297), .Y(n_406) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g339 ( .A(n_212), .Y(n_339) );
NOR2x1p5_ASAP7_75t_L g409 ( .A(n_212), .B(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x4_ASAP7_75t_L g223 ( .A(n_213), .B(n_224), .Y(n_223) );
AND2x4_ASAP7_75t_SL g247 ( .A(n_213), .B(n_225), .Y(n_247) );
OR2x2_ASAP7_75t_L g251 ( .A(n_213), .B(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g286 ( .A(n_213), .Y(n_286) );
AND2x2_ASAP7_75t_L g304 ( .A(n_213), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g315 ( .A(n_213), .B(n_225), .Y(n_315) );
OR2x2_ASAP7_75t_L g377 ( .A(n_213), .B(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g394 ( .A(n_213), .B(n_325), .Y(n_394) );
INVx1_ASAP7_75t_L g426 ( .A(n_213), .Y(n_426) );
OR2x6_ASAP7_75t_L g213 ( .A(n_214), .B(n_220), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_222), .B(n_223), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_222), .B(n_303), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_223), .B(n_337), .Y(n_336) );
AOI222xp33_ASAP7_75t_L g341 ( .A1(n_223), .A2(n_342), .B1(n_347), .B2(n_349), .C1(n_352), .C2(n_355), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_223), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g369 ( .A(n_223), .B(n_248), .Y(n_369) );
AND2x2_ASAP7_75t_L g331 ( .A(n_224), .B(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g346 ( .A(n_224), .B(n_251), .Y(n_346) );
INVx3_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_225), .B(n_252), .Y(n_284) );
AND2x4_ASAP7_75t_L g305 ( .A(n_225), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g365 ( .A(n_225), .B(n_286), .Y(n_365) );
AND2x4_ASAP7_75t_L g225 ( .A(n_226), .B(n_231), .Y(n_225) );
INVx3_ASAP7_75t_L g488 ( .A(n_234), .Y(n_488) );
INVx1_ASAP7_75t_SL g245 ( .A(n_239), .Y(n_245) );
NAND2xp33_ASAP7_75t_SL g414 ( .A(n_239), .B(n_269), .Y(n_414) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_244), .C(n_246), .Y(n_240) );
INVx2_ASAP7_75t_SL g291 ( .A(n_241), .Y(n_291) );
AND2x2_ASAP7_75t_L g295 ( .A(n_242), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_243), .B(n_291), .Y(n_290) );
O2A1O1Ixp33_ASAP7_75t_L g316 ( .A1(n_243), .A2(n_281), .B(n_317), .C(n_318), .Y(n_316) );
AND2x2_ASAP7_75t_L g393 ( .A(n_243), .B(n_374), .Y(n_393) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
AND2x4_ASAP7_75t_L g292 ( .A(n_247), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_SL g397 ( .A(n_247), .Y(n_397) );
OAI211xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_253), .B(n_260), .C(n_287), .Y(n_250) );
INVx2_ASAP7_75t_L g262 ( .A(n_251), .Y(n_262) );
OR2x2_ASAP7_75t_L g309 ( .A(n_251), .B(n_310), .Y(n_309) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_252), .Y(n_293) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_255), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g347 ( .A(n_255), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_255), .B(n_335), .Y(n_401) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AOI222xp33_ASAP7_75t_L g359 ( .A1(n_257), .A2(n_360), .B1(n_361), .B2(n_363), .C1(n_366), .C2(n_369), .Y(n_359) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_258), .A2(n_323), .B1(n_326), .B2(n_327), .C(n_333), .Y(n_322) );
AND2x2_ASAP7_75t_L g360 ( .A(n_258), .B(n_317), .Y(n_360) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp33_ASAP7_75t_SL g273 ( .A(n_259), .B(n_274), .Y(n_273) );
AOI221x1_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_265), .B1(n_270), .B2(n_273), .C(n_276), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
AND2x2_ASAP7_75t_L g413 ( .A(n_263), .B(n_351), .Y(n_413) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g271 ( .A(n_264), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
INVx1_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
OAI32xp33_ASAP7_75t_L g379 ( .A1(n_269), .A2(n_310), .A3(n_380), .B1(n_382), .B2(n_386), .Y(n_379) );
OAI21xp33_ASAP7_75t_SL g398 ( .A1(n_270), .A2(n_399), .B(n_400), .Y(n_398) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AOI21xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_280), .B(n_283), .Y(n_276) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
OR2x2_ASAP7_75t_L g280 ( .A(n_278), .B(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g353 ( .A(n_278), .B(n_354), .Y(n_353) );
AOI221xp5_ASAP7_75t_L g307 ( .A1(n_282), .A2(n_308), .B1(n_311), .B2(n_312), .C(n_316), .Y(n_307) );
INVx1_ASAP7_75t_L g383 ( .A(n_282), .Y(n_383) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_282), .Y(n_389) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
OAI21xp33_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_289), .B(n_292), .Y(n_287) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_291), .B(n_356), .Y(n_355) );
OAI21xp5_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_299), .B(n_307), .Y(n_294) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_298), .Y(n_368) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_304), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_301), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVxp67_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g320 ( .A(n_303), .Y(n_320) );
INVx1_ASAP7_75t_L g310 ( .A(n_305), .Y(n_310) );
AND2x2_ASAP7_75t_SL g319 ( .A(n_305), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_305), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_305), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g324 ( .A(n_315), .B(n_325), .Y(n_324) );
INVx2_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_320), .Y(n_385) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_322), .B(n_341), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g337 ( .A(n_325), .Y(n_337) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_SL g351 ( .A(n_329), .Y(n_351) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_331), .B(n_409), .Y(n_408) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_332), .Y(n_345) );
BUFx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_SL g342 ( .A(n_343), .B(n_346), .Y(n_342) );
INVxp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g356 ( .A(n_348), .Y(n_356) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g375 ( .A(n_354), .Y(n_375) );
NOR4xp25_ASAP7_75t_L g357 ( .A(n_358), .B(n_391), .C(n_402), .D(n_415), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_370), .Y(n_358) );
O2A1O1Ixp33_ASAP7_75t_L g370 ( .A1(n_360), .A2(n_371), .B(n_376), .C(n_379), .Y(n_370) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g372 ( .A(n_373), .B(n_375), .Y(n_372) );
OAI211xp5_ASAP7_75t_L g382 ( .A1(n_373), .A2(n_383), .B(n_384), .C(n_385), .Y(n_382) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
OAI21xp33_ASAP7_75t_SL g386 ( .A1(n_387), .A2(n_389), .B(n_390), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_SL g421 ( .A(n_390), .B(n_422), .Y(n_421) );
OAI221xp5_ASAP7_75t_SL g391 ( .A1(n_392), .A2(n_394), .B1(n_395), .B2(n_396), .C(n_398), .Y(n_391) );
INVx1_ASAP7_75t_SL g395 ( .A(n_393), .Y(n_395) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NAND3xp33_ASAP7_75t_SL g402 ( .A(n_403), .B(n_404), .C(n_411), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_407), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI21xp33_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_418), .B(n_420), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVxp33_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_428), .Y(n_427) );
CKINVDCx11_ASAP7_75t_R g748 ( .A(n_428), .Y(n_748) );
AND2x6_ASAP7_75t_SL g428 ( .A(n_429), .B(n_430), .Y(n_428) );
OR2x6_ASAP7_75t_SL g742 ( .A(n_429), .B(n_743), .Y(n_742) );
OR2x2_ASAP7_75t_L g746 ( .A(n_429), .B(n_430), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_429), .B(n_743), .Y(n_757) );
CKINVDCx5p33_ASAP7_75t_R g743 ( .A(n_430), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx2_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_436), .B(n_665), .Y(n_435) );
NOR2xp67_ASAP7_75t_L g436 ( .A(n_437), .B(n_584), .Y(n_436) );
NAND5xp2_ASAP7_75t_L g437 ( .A(n_438), .B(n_528), .C(n_538), .D(n_555), .E(n_571), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_464), .B1(n_506), .B2(n_510), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_450), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x4_ASAP7_75t_L g512 ( .A(n_442), .B(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g530 ( .A(n_442), .B(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g551 ( .A(n_442), .B(n_552), .Y(n_551) );
INVx4_ASAP7_75t_L g565 ( .A(n_442), .Y(n_565) );
AND2x2_ASAP7_75t_L g574 ( .A(n_442), .B(n_575), .Y(n_574) );
AND2x4_ASAP7_75t_SL g596 ( .A(n_442), .B(n_514), .Y(n_596) );
BUFx2_ASAP7_75t_L g639 ( .A(n_442), .Y(n_639) );
AND2x2_ASAP7_75t_L g654 ( .A(n_442), .B(n_451), .Y(n_654) );
OR2x2_ASAP7_75t_L g686 ( .A(n_442), .B(n_687), .Y(n_686) );
NOR4xp25_ASAP7_75t_L g735 ( .A(n_442), .B(n_736), .C(n_737), .D(n_738), .Y(n_735) );
OR2x6_ASAP7_75t_L g442 ( .A(n_443), .B(n_449), .Y(n_442) );
AOI31xp33_ASAP7_75t_L g603 ( .A1(n_450), .A2(n_604), .A3(n_606), .B(n_608), .Y(n_603) );
INVx2_ASAP7_75t_SL g720 ( .A(n_450), .Y(n_720) );
OR2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_459), .Y(n_450) );
INVx2_ASAP7_75t_L g527 ( .A(n_451), .Y(n_527) );
AND2x2_ASAP7_75t_L g531 ( .A(n_451), .B(n_515), .Y(n_531) );
INVx2_ASAP7_75t_L g554 ( .A(n_451), .Y(n_554) );
AND2x2_ASAP7_75t_L g573 ( .A(n_451), .B(n_514), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_457), .Y(n_452) );
AND2x2_ASAP7_75t_L g525 ( .A(n_459), .B(n_526), .Y(n_525) );
BUFx3_ASAP7_75t_L g532 ( .A(n_459), .Y(n_532) );
INVx2_ASAP7_75t_L g550 ( .A(n_459), .Y(n_550) );
AND2x2_ASAP7_75t_L g605 ( .A(n_459), .B(n_565), .Y(n_605) );
AND2x4_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
AND2x4_ASAP7_75t_L g576 ( .A(n_460), .B(n_461), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_496), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_484), .Y(n_465) );
OR2x2_ASAP7_75t_L g506 ( .A(n_466), .B(n_507), .Y(n_506) );
INVx3_ASAP7_75t_L g657 ( .A(n_466), .Y(n_657) );
OR2x2_ASAP7_75t_L g705 ( .A(n_466), .B(n_706), .Y(n_705) );
NAND2x1_ASAP7_75t_L g466 ( .A(n_467), .B(n_475), .Y(n_466) );
OR2x2_ASAP7_75t_SL g497 ( .A(n_467), .B(n_498), .Y(n_497) );
INVx4_ASAP7_75t_L g535 ( .A(n_467), .Y(n_535) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_467), .Y(n_579) );
INVx2_ASAP7_75t_L g587 ( .A(n_467), .Y(n_587) );
OR2x2_ASAP7_75t_L g622 ( .A(n_467), .B(n_486), .Y(n_622) );
AND2x2_ASAP7_75t_L g734 ( .A(n_467), .B(n_589), .Y(n_734) );
AND2x2_ASAP7_75t_L g739 ( .A(n_467), .B(n_499), .Y(n_739) );
OR2x6_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
OR2x2_ASAP7_75t_L g498 ( .A(n_475), .B(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g563 ( .A(n_475), .B(n_485), .Y(n_563) );
OR2x2_ASAP7_75t_L g570 ( .A(n_475), .B(n_535), .Y(n_570) );
NOR2x1_ASAP7_75t_SL g589 ( .A(n_475), .B(n_509), .Y(n_589) );
BUFx2_ASAP7_75t_L g621 ( .A(n_475), .Y(n_621) );
AND2x2_ASAP7_75t_L g630 ( .A(n_475), .B(n_535), .Y(n_630) );
AND2x2_ASAP7_75t_L g663 ( .A(n_475), .B(n_583), .Y(n_663) );
INVx2_ASAP7_75t_SL g672 ( .A(n_475), .Y(n_672) );
AND2x2_ASAP7_75t_L g675 ( .A(n_475), .B(n_486), .Y(n_675) );
OR2x6_ASAP7_75t_L g475 ( .A(n_476), .B(n_483), .Y(n_475) );
NAND3xp33_ASAP7_75t_L g670 ( .A(n_484), .B(n_540), .C(n_625), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_484), .B(n_587), .Y(n_690) );
INVxp67_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_485), .B(n_672), .Y(n_693) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_486), .Y(n_537) );
AND2x2_ASAP7_75t_L g581 ( .A(n_486), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g646 ( .A(n_486), .B(n_647), .Y(n_646) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_489), .B(n_495), .Y(n_487) );
AO21x1_ASAP7_75t_SL g509 ( .A1(n_488), .A2(n_489), .B(n_495), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_494), .Y(n_489) );
AND2x4_ASAP7_75t_L g541 ( .A(n_496), .B(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OR2x2_ASAP7_75t_L g677 ( .A(n_498), .B(n_622), .Y(n_677) );
AND2x2_ASAP7_75t_L g508 ( .A(n_499), .B(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g545 ( .A(n_499), .Y(n_545) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_499), .Y(n_562) );
INVx2_ASAP7_75t_L g583 ( .A(n_499), .Y(n_583) );
INVx1_ASAP7_75t_L g647 ( .A(n_499), .Y(n_647) );
INVx2_ASAP7_75t_L g729 ( .A(n_506), .Y(n_729) );
OR2x2_ASAP7_75t_L g593 ( .A(n_507), .B(n_570), .Y(n_593) );
INVx2_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g733 ( .A(n_508), .B(n_630), .Y(n_733) );
AND2x2_ASAP7_75t_L g626 ( .A(n_509), .B(n_583), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_523), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_512), .A2(n_640), .B1(n_657), .B2(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g553 ( .A(n_514), .Y(n_553) );
AND2x2_ASAP7_75t_L g607 ( .A(n_514), .B(n_527), .Y(n_607) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_514), .Y(n_634) );
INVx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_515), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_521), .Y(n_516) );
INVxp67_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_525), .B(n_639), .Y(n_638) );
OAI32xp33_ASAP7_75t_L g655 ( .A1(n_525), .A2(n_656), .A3(n_658), .B1(n_659), .B2(n_661), .Y(n_655) );
BUFx2_ASAP7_75t_L g540 ( .A(n_526), .Y(n_540) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g682 ( .A(n_527), .B(n_576), .Y(n_682) );
OR4x1_ASAP7_75t_L g528 ( .A(n_529), .B(n_532), .C(n_533), .D(n_536), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_529), .A2(n_620), .B1(n_714), .B2(n_715), .Y(n_713) );
INVx2_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_530), .Y(n_722) );
AND2x2_ASAP7_75t_L g564 ( .A(n_531), .B(n_565), .Y(n_564) );
BUFx2_ASAP7_75t_L g644 ( .A(n_531), .Y(n_644) );
INVx1_ASAP7_75t_L g660 ( .A(n_531), .Y(n_660) );
INVx1_ASAP7_75t_L g695 ( .A(n_531), .Y(n_695) );
OR2x2_ASAP7_75t_L g652 ( .A(n_532), .B(n_653), .Y(n_652) );
OR2x2_ASAP7_75t_L g696 ( .A(n_532), .B(n_697), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_533), .A2(n_570), .B1(n_614), .B2(n_633), .Y(n_635) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g679 ( .A(n_534), .B(n_588), .Y(n_679) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx2_ASAP7_75t_L g546 ( .A(n_535), .Y(n_546) );
NOR2xp67_ASAP7_75t_L g561 ( .A(n_535), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g542 ( .A(n_536), .Y(n_542) );
NAND4xp25_ASAP7_75t_L g669 ( .A(n_536), .B(n_540), .C(n_621), .D(n_633), .Y(n_669) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g706 ( .A(n_537), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_541), .B1(n_543), .B2(n_547), .Y(n_538) );
OAI22xp33_ASAP7_75t_L g689 ( .A1(n_539), .A2(n_540), .B1(n_690), .B2(n_691), .Y(n_689) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVxp67_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
INVx3_ASAP7_75t_L g568 ( .A(n_545), .Y(n_568) );
AOI32xp33_ASAP7_75t_L g684 ( .A1(n_545), .A2(n_685), .A3(n_689), .B1(n_694), .B2(n_698), .Y(n_684) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_551), .Y(n_547) );
NOR2xp67_ASAP7_75t_L g590 ( .A(n_548), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g643 ( .A(n_548), .B(n_644), .Y(n_643) );
AOI221xp5_ASAP7_75t_L g667 ( .A1(n_548), .A2(n_556), .B1(n_668), .B2(n_673), .C(n_676), .Y(n_667) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g600 ( .A(n_549), .B(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g715 ( .A(n_549), .B(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_550), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g557 ( .A(n_552), .Y(n_557) );
AND2x2_ASAP7_75t_L g575 ( .A(n_552), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
INVx1_ASAP7_75t_SL g615 ( .A(n_553), .Y(n_615) );
INVx1_ASAP7_75t_L g599 ( .A(n_554), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_558), .B1(n_564), .B2(n_566), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OR2x2_ASAP7_75t_L g701 ( .A(n_557), .B(n_631), .Y(n_701) );
INVx1_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g641 ( .A(n_560), .Y(n_641) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
AND2x2_ASAP7_75t_L g572 ( .A(n_565), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_565), .B(n_602), .Y(n_601) );
NAND2x1p5_ASAP7_75t_L g614 ( .A(n_565), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_565), .B(n_607), .Y(n_728) );
AOI22xp33_ASAP7_75t_SL g725 ( .A1(n_566), .A2(n_726), .B1(n_727), .B2(n_729), .Y(n_725) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
OR2x2_ASAP7_75t_L g608 ( .A(n_568), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g618 ( .A(n_568), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_568), .B(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_568), .B(n_672), .Y(n_671) );
AND2x4_ASAP7_75t_SL g673 ( .A(n_568), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g649 ( .A(n_570), .B(n_650), .Y(n_649) );
OAI21xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_574), .B(n_577), .Y(n_571) );
INVx1_ASAP7_75t_L g591 ( .A(n_573), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_574), .A2(n_611), .B1(n_618), .B2(n_623), .Y(n_610) );
INVx3_ASAP7_75t_L g613 ( .A(n_576), .Y(n_613) );
INVx2_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
OAI32xp33_ASAP7_75t_SL g668 ( .A1(n_579), .A2(n_639), .A3(n_669), .B1(n_670), .B2(n_671), .Y(n_668) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g588 ( .A(n_582), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND4xp25_ASAP7_75t_SL g584 ( .A(n_585), .B(n_610), .C(n_627), .D(n_642), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_590), .B1(n_592), .B2(n_594), .C(n_603), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx2_ASAP7_75t_L g625 ( .A(n_587), .Y(n_625) );
AND2x2_ASAP7_75t_L g674 ( .A(n_587), .B(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_587), .B(n_626), .Y(n_712) );
AND2x2_ASAP7_75t_L g723 ( .A(n_587), .B(n_646), .Y(n_723) );
INVx2_ASAP7_75t_L g609 ( .A(n_589), .Y(n_609) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OAI21xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_597), .B(n_600), .Y(n_594) );
AND2x2_ASAP7_75t_L g726 ( .A(n_595), .B(n_597), .Y(n_726) );
INVx2_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_596), .B(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g703 ( .A(n_601), .Y(n_703) );
INVx1_ASAP7_75t_L g688 ( .A(n_602), .Y(n_688) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_605), .B(n_660), .Y(n_659) );
NOR2x1_ASAP7_75t_L g617 ( .A(n_606), .B(n_613), .Y(n_617) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_SL g716 ( .A(n_607), .Y(n_716) );
INVx1_ASAP7_75t_L g698 ( .A(n_609), .Y(n_698) );
OR2x2_ASAP7_75t_L g714 ( .A(n_609), .B(n_625), .Y(n_714) );
NAND2xp33_ASAP7_75t_SL g611 ( .A(n_612), .B(n_616), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx2_ASAP7_75t_L g631 ( .A(n_613), .Y(n_631) );
AND2x2_ASAP7_75t_L g636 ( .A(n_613), .B(n_626), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_613), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g710 ( .A(n_614), .Y(n_710) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_619), .A2(n_700), .B1(n_702), .B2(n_704), .Y(n_699) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
INVx1_ASAP7_75t_L g664 ( .A(n_622), .Y(n_664) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
INVx1_ASAP7_75t_L g650 ( .A(n_626), .Y(n_650) );
AOI322xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_631), .A3(n_632), .B1(n_635), .B2(n_636), .C1(n_637), .C2(n_640), .Y(n_627) );
OAI21xp5_ASAP7_75t_SL g678 ( .A1(n_628), .A2(n_679), .B(n_680), .Y(n_678) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g645 ( .A(n_630), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g702 ( .A(n_631), .B(n_703), .Y(n_702) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_638), .B(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g658 ( .A(n_639), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_639), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_645), .B1(n_648), .B2(n_651), .C(n_655), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g730 ( .A1(n_644), .A2(n_731), .B1(n_733), .B2(n_734), .C(n_735), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_646), .B(n_657), .Y(n_656) );
BUFx2_ASAP7_75t_L g697 ( .A(n_647), .Y(n_697) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OAI21xp5_ASAP7_75t_L g721 ( .A1(n_651), .A2(n_722), .B(n_723), .Y(n_721) );
INVx1_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND2xp33_ASAP7_75t_SL g731 ( .A(n_660), .B(n_732), .Y(n_731) );
INVx3_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x4_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
NOR4xp75_ASAP7_75t_L g665 ( .A(n_666), .B(n_683), .C(n_707), .D(n_724), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_678), .Y(n_666) );
INVx1_ASAP7_75t_L g737 ( .A(n_675), .Y(n_737) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g709 ( .A(n_682), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g736 ( .A(n_682), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_684), .B(n_699), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_SL g732 ( .A(n_703), .Y(n_732) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NAND3x1_ASAP7_75t_L g707 ( .A(n_708), .B(n_717), .C(n_721), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_711), .B(n_713), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVxp67_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_730), .Y(n_724) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
CKINVDCx5p33_ASAP7_75t_R g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_SL g749 ( .A(n_741), .Y(n_749) );
CKINVDCx11_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVxp67_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
AOI21xp5_ASAP7_75t_L g759 ( .A1(n_751), .A2(n_756), .B(n_760), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
BUFx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_756), .Y(n_755) );
BUFx3_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
BUFx2_ASAP7_75t_L g766 ( .A(n_757), .Y(n_766) );
BUFx3_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
CKINVDCx5p33_ASAP7_75t_R g770 ( .A(n_763), .Y(n_770) );
INVx2_ASAP7_75t_SL g763 ( .A(n_764), .Y(n_763) );
NAND2xp5_ASAP7_75t_SL g764 ( .A(n_765), .B(n_767), .Y(n_764) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
endmodule