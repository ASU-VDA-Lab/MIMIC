module fake_jpeg_2490_n_590 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_590);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_590;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_4),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_57),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_58),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_64),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_17),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_65),
.B(n_74),
.Y(n_128)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_66),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_67),
.Y(n_175)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_70),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_71),
.Y(n_212)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_72),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_73),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_38),
.B(n_34),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_76),
.Y(n_147)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_17),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_79),
.B(n_84),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_80),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_81),
.Y(n_184)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_83),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_25),
.B(n_18),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_86),
.Y(n_201)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx5_ASAP7_75t_SL g156 ( 
.A(n_87),
.Y(n_156)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_88),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_89),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_18),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_90),
.B(n_122),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_91),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_93),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_19),
.Y(n_94)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_96),
.Y(n_139)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_100),
.Y(n_164)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_103),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_24),
.Y(n_105)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_105),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_20),
.Y(n_106)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_106),
.Y(n_180)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_32),
.Y(n_107)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_107),
.Y(n_185)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_108),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_32),
.Y(n_109)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_109),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_32),
.Y(n_110)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_110),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_111),
.Y(n_194)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_36),
.Y(n_112)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_112),
.Y(n_199)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_36),
.Y(n_114)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_114),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_39),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_43),
.Y(n_144)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_24),
.Y(n_116)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_39),
.Y(n_117)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_117),
.Y(n_202)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_34),
.Y(n_118)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_118),
.Y(n_182)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_23),
.Y(n_119)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_27),
.Y(n_120)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_37),
.Y(n_121)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_121),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_38),
.B(n_18),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_38),
.Y(n_123)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_123),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_37),
.Y(n_124)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_124),
.Y(n_203)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_42),
.Y(n_125)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_125),
.Y(n_205)
);

INVx3_ASAP7_75t_SL g126 ( 
.A(n_23),
.Y(n_126)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_126),
.Y(n_213)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_42),
.Y(n_127)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_127),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_65),
.B(n_43),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_133),
.B(n_149),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_84),
.A2(n_26),
.B1(n_55),
.B2(n_54),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_135),
.B(n_220),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_79),
.A2(n_120),
.B1(n_90),
.B2(n_47),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_143),
.A2(n_28),
.B1(n_27),
.B2(n_100),
.Y(n_224)
);

INVx3_ASAP7_75t_SL g289 ( 
.A(n_144),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_56),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_145),
.B(n_159),
.Y(n_221)
);

INVx6_ASAP7_75t_SL g146 ( 
.A(n_57),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_146),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_26),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_123),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_157),
.B(n_12),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_59),
.B(n_54),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_117),
.B(n_56),
.C(n_55),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_163),
.B(n_23),
.C(n_52),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_81),
.B(n_48),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_165),
.B(n_170),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_86),
.B(n_53),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_92),
.B(n_53),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_176),
.B(n_177),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_61),
.B(n_49),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_63),
.B(n_49),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_178),
.B(n_15),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_67),
.B(n_48),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_183),
.B(n_191),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_94),
.B(n_41),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_70),
.A2(n_110),
.B1(n_109),
.B2(n_103),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_193),
.A2(n_214),
.B1(n_28),
.B2(n_99),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_71),
.B(n_41),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_196),
.B(n_198),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_73),
.B(n_35),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_78),
.B(n_35),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_204),
.B(n_207),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_80),
.B(n_47),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_89),
.B(n_47),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_210),
.B(n_216),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_91),
.A2(n_29),
.B1(n_28),
.B2(n_27),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_93),
.B(n_29),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_96),
.B(n_29),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_151),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_222),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_161),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_223),
.Y(n_327)
);

OAI21xp33_ASAP7_75t_SL g324 ( 
.A1(n_224),
.A2(n_262),
.B(n_286),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_161),
.Y(n_226)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_226),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_228),
.A2(n_277),
.B1(n_284),
.B2(n_285),
.Y(n_346)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_152),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_230),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_143),
.A2(n_23),
.B1(n_52),
.B2(n_4),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_231),
.A2(n_260),
.B1(n_278),
.B2(n_204),
.Y(n_305)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_132),
.Y(n_232)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_232),
.Y(n_336)
);

AO22x2_ASAP7_75t_L g233 ( 
.A1(n_219),
.A2(n_52),
.B1(n_23),
.B2(n_4),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_233),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_156),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_234),
.B(n_255),
.Y(n_308)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_130),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_235),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_128),
.B(n_2),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_236),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_237),
.B(n_250),
.Y(n_301)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_168),
.Y(n_238)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_238),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_192),
.Y(n_239)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_239),
.Y(n_318)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_154),
.Y(n_240)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_240),
.Y(n_313)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_182),
.Y(n_241)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_241),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_136),
.A2(n_23),
.B1(n_52),
.B2(n_5),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_242),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_159),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_243),
.Y(n_331)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_148),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_244),
.Y(n_307)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_155),
.Y(n_245)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_245),
.Y(n_314)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_173),
.Y(n_246)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_246),
.Y(n_325)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_190),
.Y(n_247)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_247),
.Y(n_340)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_211),
.Y(n_249)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_249),
.Y(n_352)
);

AOI32xp33_ASAP7_75t_L g250 ( 
.A1(n_136),
.A2(n_52),
.A3(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_203),
.Y(n_252)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_252),
.Y(n_338)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_190),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_254),
.Y(n_354)
);

A2O1A1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_142),
.A2(n_52),
.B(n_6),
.C(n_8),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_172),
.Y(n_256)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_256),
.Y(n_348)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_199),
.Y(n_257)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_257),
.Y(n_350)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_130),
.Y(n_258)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_258),
.Y(n_302)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_218),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_259),
.B(n_264),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_L g260 ( 
.A1(n_194),
.A2(n_3),
.B1(n_6),
.B2(n_8),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_213),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_261),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_179),
.A2(n_3),
.B1(n_8),
.B2(n_9),
.Y(n_262)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_208),
.Y(n_263)
);

INVx5_ASAP7_75t_L g341 ( 
.A(n_263),
.Y(n_341)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_200),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_141),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_267),
.B(n_274),
.Y(n_315)
);

INVx8_ASAP7_75t_L g268 ( 
.A(n_139),
.Y(n_268)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_268),
.Y(n_310)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_184),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_269),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_141),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_270),
.Y(n_345)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_164),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_271),
.B(n_272),
.Y(n_337)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_195),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_205),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_273),
.B(n_275),
.Y(n_343)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_207),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_185),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_276),
.B(n_279),
.Y(n_353)
);

INVx8_ASAP7_75t_L g277 ( 
.A(n_139),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_193),
.A2(n_3),
.B1(n_9),
.B2(n_10),
.Y(n_278)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_150),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_188),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_280),
.B(n_282),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_128),
.B(n_3),
.Y(n_281)
);

NAND2x1_ASAP7_75t_SL g321 ( 
.A(n_281),
.B(n_283),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_180),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_210),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_216),
.Y(n_284)
);

BUFx8_ASAP7_75t_L g285 ( 
.A(n_201),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_144),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_142),
.B(n_11),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_287),
.B(n_292),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_220),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_288),
.A2(n_291),
.B1(n_293),
.B2(n_294),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_137),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_149),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_174),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_150),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_165),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_296),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_196),
.B(n_15),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_298),
.Y(n_317)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_187),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_140),
.A2(n_14),
.B1(n_147),
.B2(n_215),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_299),
.A2(n_214),
.B1(n_191),
.B2(n_153),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_305),
.A2(n_312),
.B1(n_320),
.B2(n_344),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_266),
.A2(n_198),
.B1(n_186),
.B2(n_197),
.Y(n_312)
);

NOR2x1_ASAP7_75t_R g316 ( 
.A(n_237),
.B(n_176),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_316),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_253),
.B(n_129),
.C(n_170),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_319),
.B(n_333),
.C(n_335),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_227),
.A2(n_202),
.B1(n_209),
.B2(n_217),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_322),
.Y(n_380)
);

OAI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_251),
.A2(n_243),
.B1(n_224),
.B2(n_229),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_329),
.A2(n_255),
.B1(n_233),
.B2(n_265),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_248),
.B(n_160),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_330),
.B(n_288),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_221),
.B(n_138),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_225),
.B(n_166),
.C(n_158),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_227),
.A2(n_217),
.B1(n_212),
.B2(n_181),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_289),
.A2(n_171),
.B1(n_206),
.B2(n_162),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_349),
.A2(n_289),
.B1(n_226),
.B2(n_223),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_331),
.B(n_290),
.Y(n_356)
);

INVxp33_ASAP7_75t_L g408 ( 
.A(n_356),
.Y(n_408)
);

XNOR2x1_ASAP7_75t_L g357 ( 
.A(n_333),
.B(n_319),
.Y(n_357)
);

MAJx2_ASAP7_75t_L g411 ( 
.A(n_357),
.B(n_303),
.C(n_311),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_358),
.B(n_362),
.Y(n_401)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_307),
.Y(n_359)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_359),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_316),
.B(n_239),
.C(n_236),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_361),
.B(n_390),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_320),
.B(n_312),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_364),
.A2(n_385),
.B(n_387),
.Y(n_404)
);

INVx5_ASAP7_75t_L g365 ( 
.A(n_342),
.Y(n_365)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_365),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_366),
.B(n_374),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_300),
.A2(n_233),
.B1(n_260),
.B2(n_276),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_367),
.A2(n_370),
.B1(n_373),
.B2(n_394),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_300),
.A2(n_233),
.B1(n_299),
.B2(n_281),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_368),
.A2(n_381),
.B1(n_383),
.B2(n_345),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_331),
.B(n_282),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_369),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_308),
.A2(n_244),
.B1(n_263),
.B2(n_267),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_304),
.Y(n_371)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_371),
.Y(n_406)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_304),
.Y(n_372)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_372),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_305),
.A2(n_212),
.B1(n_181),
.B2(n_175),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_317),
.B(n_286),
.Y(n_374)
);

INVx6_ASAP7_75t_L g375 ( 
.A(n_342),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_375),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_317),
.B(n_249),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_376),
.B(n_386),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_334),
.B(n_291),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_377),
.B(n_398),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_346),
.A2(n_285),
.B(n_262),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_378),
.A2(n_347),
.B(n_353),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_301),
.A2(n_167),
.B1(n_169),
.B2(n_131),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_326),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_382),
.B(n_384),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_330),
.A2(n_258),
.B1(n_235),
.B2(n_175),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_337),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_324),
.A2(n_285),
.B(n_270),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_309),
.B(n_272),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_328),
.A2(n_268),
.B(n_277),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_326),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_388),
.B(n_391),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_321),
.A2(n_294),
.B(n_134),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_389),
.A2(n_341),
.B(n_354),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_344),
.B(n_232),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_338),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_338),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_392),
.B(n_393),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_332),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_309),
.A2(n_323),
.B1(n_335),
.B2(n_349),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_343),
.B(n_315),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_395),
.B(n_340),
.Y(n_434)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_318),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_396),
.B(n_397),
.Y(n_428)
);

INVx8_ASAP7_75t_L g397 ( 
.A(n_310),
.Y(n_397)
);

BUFx24_ASAP7_75t_SL g398 ( 
.A(n_321),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_400),
.A2(n_418),
.B(n_423),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_385),
.A2(n_339),
.B(n_351),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_403),
.A2(n_407),
.B(n_424),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_378),
.A2(n_303),
.B(n_336),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_380),
.A2(n_318),
.B1(n_302),
.B2(n_131),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_410),
.A2(n_412),
.B1(n_422),
.B2(n_390),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_411),
.B(n_413),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_380),
.A2(n_302),
.B1(n_307),
.B2(n_352),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_414),
.A2(n_421),
.B1(n_426),
.B2(n_427),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_363),
.A2(n_336),
.B(n_327),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_368),
.A2(n_352),
.B1(n_306),
.B2(n_350),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_367),
.A2(n_189),
.B1(n_350),
.B2(n_348),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_387),
.A2(n_310),
.B(n_354),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_363),
.A2(n_340),
.B(n_355),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_425),
.A2(n_430),
.B(n_389),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_379),
.A2(n_348),
.B1(n_341),
.B2(n_313),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_373),
.A2(n_313),
.B1(n_314),
.B2(n_325),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_394),
.A2(n_360),
.B1(n_386),
.B2(n_362),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_429),
.A2(n_383),
.B1(n_391),
.B2(n_397),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_366),
.A2(n_269),
.B(n_314),
.Y(n_430)
);

NAND3xp33_ASAP7_75t_L g437 ( 
.A(n_434),
.B(n_395),
.C(n_374),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_435),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_432),
.B(n_376),
.Y(n_436)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_436),
.Y(n_494)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_437),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_409),
.A2(n_360),
.B(n_396),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_438),
.A2(n_425),
.B(n_403),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_411),
.B(n_357),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_439),
.B(n_451),
.C(n_453),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_412),
.A2(n_362),
.B1(n_390),
.B2(n_358),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_442),
.A2(n_447),
.B1(n_456),
.B2(n_440),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_402),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_443),
.B(n_446),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_417),
.Y(n_444)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_444),
.Y(n_478)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_416),
.Y(n_445)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_445),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_416),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_412),
.A2(n_409),
.B1(n_421),
.B2(n_401),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_447),
.A2(n_457),
.B1(n_405),
.B2(n_422),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_432),
.B(n_393),
.Y(n_448)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_448),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_408),
.B(n_372),
.Y(n_449)
);

NAND3xp33_ASAP7_75t_L g486 ( 
.A(n_449),
.B(n_450),
.C(n_463),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_431),
.B(n_392),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_413),
.B(n_361),
.C(n_381),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_406),
.Y(n_452)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_452),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_413),
.B(n_371),
.C(n_382),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_434),
.B(n_388),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_454),
.B(n_456),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_455),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_421),
.A2(n_375),
.B1(n_365),
.B2(n_359),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_417),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_458),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_418),
.Y(n_459)
);

CKINVDCx14_ASAP7_75t_R g490 ( 
.A(n_459),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_405),
.A2(n_327),
.B1(n_325),
.B2(n_279),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_461),
.A2(n_427),
.B1(n_414),
.B2(n_424),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_462),
.B(n_404),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_415),
.B(n_428),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_411),
.B(n_429),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_464),
.B(n_466),
.C(n_462),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_428),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_465),
.B(n_467),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_401),
.B(n_404),
.C(n_418),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_415),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_469),
.B(n_479),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_470),
.B(n_458),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_472),
.B(n_484),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_474),
.A2(n_497),
.B1(n_440),
.B2(n_448),
.Y(n_511)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_475),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_451),
.B(n_401),
.C(n_430),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_476),
.B(n_488),
.C(n_495),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_455),
.A2(n_401),
.B1(n_407),
.B2(n_426),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_477),
.A2(n_480),
.B1(n_442),
.B2(n_457),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_464),
.B(n_423),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_460),
.A2(n_426),
.B1(n_400),
.B2(n_414),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_439),
.B(n_433),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_460),
.A2(n_441),
.B(n_466),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_485),
.A2(n_491),
.B(n_435),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_438),
.B(n_433),
.C(n_406),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_441),
.A2(n_410),
.B(n_420),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_453),
.B(n_399),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_489),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_500),
.B(n_504),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_483),
.B(n_446),
.Y(n_503)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_503),
.Y(n_527)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_489),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_481),
.B(n_445),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_505),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_506),
.B(n_515),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_SL g533 ( 
.A(n_507),
.B(n_509),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_496),
.B(n_465),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_508),
.B(n_519),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_SL g509 ( 
.A(n_470),
.B(n_436),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_468),
.B(n_467),
.C(n_444),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_510),
.B(n_520),
.C(n_472),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_511),
.A2(n_512),
.B1(n_517),
.B2(n_518),
.Y(n_523)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_493),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_513),
.A2(n_493),
.B1(n_490),
.B2(n_491),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_486),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_514),
.B(n_469),
.Y(n_530)
);

NAND2x1_ASAP7_75t_L g515 ( 
.A(n_471),
.B(n_454),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_SL g516 ( 
.A(n_484),
.B(n_463),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_516),
.B(n_488),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_487),
.A2(n_449),
.B1(n_450),
.B2(n_452),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_473),
.A2(n_427),
.B1(n_443),
.B2(n_419),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_496),
.B(n_419),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_468),
.B(n_402),
.C(n_420),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_482),
.B(n_399),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_521),
.B(n_478),
.Y(n_534)
);

XOR2x1_ASAP7_75t_SL g525 ( 
.A(n_502),
.B(n_515),
.Y(n_525)
);

A2O1A1Ixp33_ASAP7_75t_L g541 ( 
.A1(n_525),
.A2(n_485),
.B(n_506),
.C(n_508),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_510),
.B(n_495),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_526),
.B(n_531),
.Y(n_547)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_530),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_512),
.A2(n_497),
.B1(n_474),
.B2(n_487),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_532),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_534),
.B(n_505),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_499),
.A2(n_471),
.B1(n_477),
.B2(n_480),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_535),
.A2(n_517),
.B1(n_519),
.B2(n_494),
.Y(n_553)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_536),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_498),
.B(n_476),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_537),
.B(n_538),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_498),
.B(n_479),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_539),
.B(n_520),
.C(n_502),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_523),
.A2(n_499),
.B1(n_513),
.B2(n_504),
.Y(n_540)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_540),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_541),
.B(n_545),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_529),
.B(n_503),
.Y(n_544)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_544),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_538),
.B(n_501),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_546),
.B(n_537),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_539),
.B(n_501),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_548),
.B(n_516),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_550),
.B(n_551),
.Y(n_560)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_527),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_553),
.B(n_522),
.Y(n_558)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_524),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_554),
.B(n_522),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_555),
.B(n_557),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_556),
.A2(n_558),
.B1(n_562),
.B2(n_565),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_546),
.B(n_526),
.C(n_531),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_542),
.B(n_494),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_559),
.B(n_563),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_541),
.A2(n_528),
.B(n_515),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_562),
.B(n_540),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_549),
.B(n_535),
.C(n_525),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_566),
.B(n_547),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_564),
.B(n_560),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_567),
.B(n_568),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_569),
.B(n_558),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_565),
.B(n_547),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_570),
.B(n_572),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_L g571 ( 
.A1(n_557),
.A2(n_563),
.B(n_543),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_571),
.A2(n_566),
.B1(n_549),
.B2(n_548),
.Y(n_576)
);

NOR2x1_ASAP7_75t_L g575 ( 
.A(n_570),
.B(n_561),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g583 ( 
.A1(n_575),
.A2(n_576),
.B(n_572),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_578),
.B(n_579),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_573),
.B(n_552),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_577),
.B(n_574),
.C(n_569),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_582),
.B(n_575),
.Y(n_584)
);

OAI31xp33_ASAP7_75t_SL g585 ( 
.A1(n_583),
.A2(n_580),
.A3(n_533),
.B(n_545),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_584),
.B(n_585),
.C(n_581),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_586),
.B(n_580),
.Y(n_587)
);

NOR3xp33_ASAP7_75t_SL g588 ( 
.A(n_587),
.B(n_492),
.C(n_507),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_588),
.B(n_475),
.Y(n_589)
);

NOR3xp33_ASAP7_75t_SL g590 ( 
.A(n_589),
.B(n_533),
.C(n_509),
.Y(n_590)
);


endmodule