module fake_netlist_5_2265_n_3830 (n_137, n_676, n_294, n_431, n_318, n_380, n_419, n_653, n_611, n_444, n_642, n_469, n_615, n_82, n_194, n_316, n_785, n_389, n_549, n_684, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_705, n_619, n_408, n_61, n_678, n_664, n_376, n_697, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_776, n_667, n_515, n_57, n_353, n_351, n_367, n_620, n_643, n_452, n_397, n_493, n_111, n_525, n_703, n_698, n_483, n_544, n_683, n_155, n_780, n_649, n_552, n_547, n_43, n_721, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_725, n_139, n_38, n_105, n_280, n_744, n_590, n_629, n_672, n_4, n_378, n_551, n_762, n_17, n_581, n_688, n_382, n_554, n_254, n_690, n_33, n_23, n_583, n_671, n_718, n_302, n_265, n_526, n_719, n_293, n_372, n_443, n_244, n_677, n_47, n_173, n_198, n_714, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_753, n_100, n_455, n_674, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_689, n_738, n_606, n_559, n_275, n_640, n_252, n_624, n_26, n_295, n_133, n_330, n_508, n_739, n_506, n_2, n_737, n_610, n_692, n_755, n_6, n_509, n_568, n_39, n_147, n_373, n_757, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_758, n_668, n_733, n_375, n_301, n_779, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_659, n_51, n_63, n_492, n_563, n_171, n_153, n_756, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_741, n_548, n_543, n_260, n_298, n_650, n_320, n_694, n_518, n_505, n_286, n_122, n_282, n_752, n_331, n_10, n_24, n_406, n_519, n_470, n_782, n_325, n_449, n_132, n_90, n_724, n_546, n_101, n_760, n_658, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_731, n_31, n_456, n_13, n_371, n_481, n_535, n_709, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_769, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_654, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_751, n_484, n_775, n_219, n_442, n_157, n_131, n_192, n_636, n_786, n_600, n_660, n_223, n_392, n_158, n_655, n_704, n_138, n_264, n_109, n_669, n_472, n_742, n_750, n_454, n_387, n_771, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_763, n_169, n_59, n_522, n_550, n_255, n_696, n_215, n_350, n_196, n_662, n_459, n_646, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_723, n_386, n_578, n_287, n_344, n_555, n_783, n_473, n_422, n_475, n_777, n_72, n_661, n_104, n_41, n_682, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_670, n_15, n_336, n_584, n_681, n_591, n_145, n_48, n_521, n_614, n_663, n_50, n_337, n_430, n_313, n_631, n_673, n_88, n_479, n_528, n_510, n_216, n_680, n_168, n_395, n_164, n_432, n_553, n_727, n_311, n_773, n_208, n_142, n_743, n_214, n_328, n_140, n_299, n_303, n_369, n_675, n_296, n_613, n_241, n_637, n_357, n_598, n_685, n_608, n_184, n_446, n_445, n_65, n_78, n_749, n_144, n_114, n_96, n_772, n_691, n_717, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_734, n_638, n_700, n_197, n_107, n_573, n_69, n_236, n_388, n_761, n_1, n_249, n_740, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_693, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_652, n_778, n_29, n_79, n_151, n_25, n_306, n_722, n_458, n_288, n_770, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_711, n_781, n_474, n_112, n_765, n_542, n_85, n_463, n_488, n_595, n_736, n_502, n_239, n_466, n_420, n_630, n_489, n_632, n_699, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_748, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_745, n_627, n_767, n_172, n_206, n_217, n_440, n_726, n_478, n_545, n_441, n_450, n_648, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_641, n_628, n_365, n_774, n_91, n_729, n_730, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_679, n_707, n_710, n_695, n_180, n_560, n_656, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_665, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_720, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_117, n_326, n_768, n_233, n_404, n_686, n_205, n_366, n_572, n_113, n_712, n_754, n_246, n_596, n_179, n_125, n_410, n_558, n_708, n_269, n_529, n_128, n_735, n_702, n_285, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_728, n_202, n_266, n_272, n_491, n_427, n_732, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_716, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_159, n_334, n_599, n_766, n_541, n_391, n_701, n_434, n_645, n_539, n_175, n_538, n_666, n_262, n_238, n_639, n_99, n_687, n_715, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_764, n_200, n_162, n_64, n_759, n_222, n_28, n_89, n_438, n_115, n_713, n_324, n_634, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_424, n_7, n_706, n_746, n_256, n_305, n_533, n_747, n_52, n_278, n_784, n_110, n_3830);

input n_137;
input n_676;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_785;
input n_389;
input n_549;
input n_684;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_705;
input n_619;
input n_408;
input n_61;
input n_678;
input n_664;
input n_376;
input n_697;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_776;
input n_667;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_703;
input n_698;
input n_483;
input n_544;
input n_683;
input n_155;
input n_780;
input n_649;
input n_552;
input n_547;
input n_43;
input n_721;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_725;
input n_139;
input n_38;
input n_105;
input n_280;
input n_744;
input n_590;
input n_629;
input n_672;
input n_4;
input n_378;
input n_551;
input n_762;
input n_17;
input n_581;
input n_688;
input n_382;
input n_554;
input n_254;
input n_690;
input n_33;
input n_23;
input n_583;
input n_671;
input n_718;
input n_302;
input n_265;
input n_526;
input n_719;
input n_293;
input n_372;
input n_443;
input n_244;
input n_677;
input n_47;
input n_173;
input n_198;
input n_714;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_753;
input n_100;
input n_455;
input n_674;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_689;
input n_738;
input n_606;
input n_559;
input n_275;
input n_640;
input n_252;
input n_624;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_739;
input n_506;
input n_2;
input n_737;
input n_610;
input n_692;
input n_755;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_757;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_758;
input n_668;
input n_733;
input n_375;
input n_301;
input n_779;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_659;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_756;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_741;
input n_548;
input n_543;
input n_260;
input n_298;
input n_650;
input n_320;
input n_694;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_752;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_782;
input n_325;
input n_449;
input n_132;
input n_90;
input n_724;
input n_546;
input n_101;
input n_760;
input n_658;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_731;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_709;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_769;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_654;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_751;
input n_484;
input n_775;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_636;
input n_786;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_704;
input n_138;
input n_264;
input n_109;
input n_669;
input n_472;
input n_742;
input n_750;
input n_454;
input n_387;
input n_771;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_763;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_696;
input n_215;
input n_350;
input n_196;
input n_662;
input n_459;
input n_646;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_723;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_783;
input n_473;
input n_422;
input n_475;
input n_777;
input n_72;
input n_661;
input n_104;
input n_41;
input n_682;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_670;
input n_15;
input n_336;
input n_584;
input n_681;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_663;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_673;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_680;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_727;
input n_311;
input n_773;
input n_208;
input n_142;
input n_743;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_675;
input n_296;
input n_613;
input n_241;
input n_637;
input n_357;
input n_598;
input n_685;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_749;
input n_144;
input n_114;
input n_96;
input n_772;
input n_691;
input n_717;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_734;
input n_638;
input n_700;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_761;
input n_1;
input n_249;
input n_740;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_693;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_778;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_722;
input n_458;
input n_288;
input n_770;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_711;
input n_781;
input n_474;
input n_112;
input n_765;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_736;
input n_502;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_699;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_748;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_745;
input n_627;
input n_767;
input n_172;
input n_206;
input n_217;
input n_440;
input n_726;
input n_478;
input n_545;
input n_441;
input n_450;
input n_648;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_641;
input n_628;
input n_365;
input n_774;
input n_91;
input n_729;
input n_730;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_679;
input n_707;
input n_710;
input n_695;
input n_180;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_665;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_720;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_768;
input n_233;
input n_404;
input n_686;
input n_205;
input n_366;
input n_572;
input n_113;
input n_712;
input n_754;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_708;
input n_269;
input n_529;
input n_128;
input n_735;
input n_702;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_728;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_732;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_716;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_159;
input n_334;
input n_599;
input n_766;
input n_541;
input n_391;
input n_701;
input n_434;
input n_645;
input n_539;
input n_175;
input n_538;
input n_666;
input n_262;
input n_238;
input n_639;
input n_99;
input n_687;
input n_715;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_764;
input n_200;
input n_162;
input n_64;
input n_759;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_713;
input n_324;
input n_634;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_424;
input n_7;
input n_706;
input n_746;
input n_256;
input n_305;
input n_533;
input n_747;
input n_52;
input n_278;
input n_784;
input n_110;

output n_3830;

wire n_924;
wire n_1263;
wire n_3304;
wire n_1378;
wire n_977;
wire n_2253;
wire n_2417;
wire n_2756;
wire n_1423;
wire n_1126;
wire n_1729;
wire n_2739;
wire n_2380;
wire n_1166;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_3241;
wire n_2617;
wire n_2200;
wire n_3261;
wire n_3006;
wire n_1161;
wire n_3795;
wire n_3027;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_3179;
wire n_3127;
wire n_1780;
wire n_3256;
wire n_3732;
wire n_1488;
wire n_2899;
wire n_2955;
wire n_790;
wire n_3619;
wire n_1055;
wire n_3541;
wire n_3622;
wire n_2386;
wire n_3596;
wire n_1501;
wire n_2395;
wire n_880;
wire n_3086;
wire n_3297;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1360;
wire n_1198;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_3641;
wire n_956;
wire n_1738;
wire n_2021;
wire n_3728;
wire n_2134;
wire n_3064;
wire n_2391;
wire n_3088;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_3713;
wire n_2853;
wire n_3615;
wire n_2059;
wire n_1323;
wire n_3663;
wire n_1466;
wire n_1695;
wire n_2487;
wire n_3766;
wire n_1353;
wire n_800;
wire n_3595;
wire n_3246;
wire n_3202;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_3813;
wire n_1789;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_3341;
wire n_1947;
wire n_1264;
wire n_3587;
wire n_2114;
wire n_3445;
wire n_2001;
wire n_1494;
wire n_3407;
wire n_3571;
wire n_3599;
wire n_3785;
wire n_1462;
wire n_1799;
wire n_854;
wire n_2069;
wire n_2396;
wire n_3621;
wire n_1580;
wire n_1939;
wire n_2486;
wire n_3434;
wire n_1806;
wire n_933;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_1152;
wire n_3501;
wire n_3448;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_3039;
wire n_3019;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_3776;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_3163;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_3710;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1728;
wire n_1107;
wire n_2031;
wire n_2076;
wire n_3036;
wire n_2482;
wire n_2677;
wire n_1230;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_3010;
wire n_3180;
wire n_3379;
wire n_3532;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_902;
wire n_1104;
wire n_1705;
wire n_1294;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_3188;
wire n_3325;
wire n_3107;
wire n_3531;
wire n_3403;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2963;
wire n_3624;
wire n_2142;
wire n_3186;
wire n_3461;
wire n_3082;
wire n_1154;
wire n_2189;
wire n_3796;
wire n_3332;
wire n_1242;
wire n_3283;
wire n_1135;
wire n_3048;
wire n_3258;
wire n_3696;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_2959;
wire n_3340;
wire n_2047;
wire n_1280;
wire n_3277;
wire n_3782;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_3650;
wire n_3786;
wire n_2761;
wire n_1483;
wire n_2888;
wire n_3638;
wire n_1314;
wire n_1512;
wire n_3157;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2983;
wire n_3763;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_3214;
wire n_2306;
wire n_920;
wire n_2515;
wire n_3022;
wire n_3810;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_3631;
wire n_2715;
wire n_3806;
wire n_3087;
wire n_2085;
wire n_3489;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_2936;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_3060;
wire n_2651;
wire n_3490;
wire n_3656;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_3013;
wire n_3183;
wire n_1984;
wire n_3437;
wire n_2099;
wire n_2408;
wire n_3446;
wire n_3353;
wire n_1877;
wire n_3687;
wire n_1831;
wire n_1598;
wire n_3049;
wire n_1723;
wire n_955;
wire n_1850;
wire n_3028;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1097;
wire n_1749;
wire n_1036;
wire n_3156;
wire n_3101;
wire n_3669;
wire n_897;
wire n_798;
wire n_3376;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_3653;
wire n_1414;
wire n_1216;
wire n_2693;
wire n_3798;
wire n_3702;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_3389;
wire n_1852;
wire n_2159;
wire n_2976;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_3089;
wire n_1547;
wire n_1070;
wire n_2089;
wire n_3420;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_3222;
wire n_1561;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_1513;
wire n_2908;
wire n_2970;
wire n_3361;
wire n_1600;
wire n_3744;
wire n_845;
wire n_2235;
wire n_1862;
wire n_837;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_3291;
wire n_1473;
wire n_1587;
wire n_2682;
wire n_901;
wire n_3755;
wire n_2432;
wire n_3668;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_3440;
wire n_3405;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_3563;
wire n_2934;
wire n_1672;
wire n_2506;
wire n_2699;
wire n_1880;
wire n_888;
wire n_2769;
wire n_3542;
wire n_2337;
wire n_3550;
wire n_1167;
wire n_1626;
wire n_3436;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_2985;
wire n_1151;
wire n_2944;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_3418;
wire n_2932;
wire n_2753;
wire n_2980;
wire n_1582;
wire n_3637;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_3262;
wire n_3136;
wire n_1836;
wire n_2868;
wire n_3395;
wire n_1450;
wire n_3141;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_3164;
wire n_2738;
wire n_1750;
wire n_3570;
wire n_3690;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_3716;
wire n_2968;
wire n_1700;
wire n_2833;
wire n_3191;
wire n_1585;
wire n_2712;
wire n_2684;
wire n_3593;
wire n_3193;
wire n_1971;
wire n_1599;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3507;
wire n_3273;
wire n_3821;
wire n_2713;
wire n_3544;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_3367;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_3008;
wire n_3709;
wire n_907;
wire n_1447;
wire n_2251;
wire n_3096;
wire n_1377;
wire n_2370;
wire n_3496;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_3339;
wire n_2055;
wire n_3427;
wire n_3025;
wire n_3349;
wire n_1403;
wire n_3735;
wire n_2248;
wire n_2356;
wire n_892;
wire n_3320;
wire n_3007;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_3714;
wire n_1463;
wire n_1581;
wire n_1002;
wire n_2100;
wire n_3071;
wire n_3739;
wire n_3651;
wire n_3310;
wire n_3487;
wire n_2258;
wire n_1667;
wire n_1058;
wire n_3359;
wire n_838;
wire n_2784;
wire n_3718;
wire n_2919;
wire n_3092;
wire n_1053;
wire n_3470;
wire n_1224;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_3676;
wire n_2150;
wire n_3146;
wire n_2241;
wire n_2757;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_963;
wire n_1052;
wire n_954;
wire n_3781;
wire n_1385;
wire n_793;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_3580;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_2987;
wire n_1527;
wire n_2042;
wire n_3106;
wire n_1882;
wire n_884;
wire n_3328;
wire n_944;
wire n_1754;
wire n_3611;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2674;
wire n_2606;
wire n_3187;
wire n_1565;
wire n_3508;
wire n_2828;
wire n_3682;
wire n_3371;
wire n_1809;
wire n_1856;
wire n_3433;
wire n_3392;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_2305;
wire n_3430;
wire n_2636;
wire n_2450;
wire n_3208;
wire n_1319;
wire n_2379;
wire n_3331;
wire n_3447;
wire n_2616;
wire n_2911;
wire n_3305;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_3528;
wire n_3649;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_3257;
wire n_3625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2331;
wire n_2945;
wire n_2293;
wire n_2837;
wire n_847;
wire n_3804;
wire n_1393;
wire n_2319;
wire n_1775;
wire n_2979;
wire n_3296;
wire n_2028;
wire n_1368;
wire n_3481;
wire n_2762;
wire n_3655;
wire n_2808;
wire n_1276;
wire n_3009;
wire n_2548;
wire n_1412;
wire n_822;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_2108;
wire n_3640;
wire n_1538;
wire n_1162;
wire n_2930;
wire n_1838;
wire n_1847;
wire n_1199;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_3514;
wire n_3116;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_3602;
wire n_1038;
wire n_2967;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_3207;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_3224;
wire n_2698;
wire n_3752;
wire n_809;
wire n_870;
wire n_931;
wire n_1711;
wire n_1891;
wire n_1662;
wire n_1481;
wire n_2626;
wire n_3441;
wire n_3042;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_3047;
wire n_3526;
wire n_868;
wire n_2454;
wire n_2804;
wire n_914;
wire n_3659;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_3120;
wire n_965;
wire n_1876;
wire n_1743;
wire n_3790;
wire n_3491;
wire n_935;
wire n_817;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_1888;
wire n_2009;
wire n_3643;
wire n_2222;
wire n_1892;
wire n_3510;
wire n_3745;
wire n_806;
wire n_2990;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_3218;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_3119;
wire n_1189;
wire n_2690;
wire n_3370;
wire n_2215;
wire n_3479;
wire n_1259;
wire n_1690;
wire n_3819;
wire n_1649;
wire n_3150;
wire n_2064;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_3500;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_3660;
wire n_2297;
wire n_1815;
wire n_3279;
wire n_2621;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_3747;
wire n_1537;
wire n_913;
wire n_865;
wire n_2227;
wire n_3775;
wire n_2671;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_3346;
wire n_1798;
wire n_2022;
wire n_3814;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_3416;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_3133;
wire n_3513;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_2992;
wire n_1674;
wire n_3725;
wire n_1833;
wire n_3138;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_3128;
wire n_1734;
wire n_3038;
wire n_3770;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_3068;
wire n_1767;
wire n_3144;
wire n_2943;
wire n_2913;
wire n_2336;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_1233;
wire n_3469;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_3317;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_3355;
wire n_2007;
wire n_3220;
wire n_949;
wire n_2539;
wire n_3263;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_3765;
wire n_1468;
wire n_1559;
wire n_3823;
wire n_1765;
wire n_3455;
wire n_1866;
wire n_3158;
wire n_1624;
wire n_3000;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_3113;
wire n_1231;
wire n_1406;
wire n_1279;
wire n_3108;
wire n_3111;
wire n_2718;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_2577;
wire n_3760;
wire n_1760;
wire n_2875;
wire n_936;
wire n_1500;
wire n_2960;
wire n_1090;
wire n_2796;
wire n_3280;
wire n_2342;
wire n_2856;
wire n_3471;
wire n_1832;
wire n_1851;
wire n_999;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_2937;
wire n_3666;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_3828;
wire n_2290;
wire n_1656;
wire n_3564;
wire n_3288;
wire n_1158;
wire n_3095;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_3199;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_3667;
wire n_1145;
wire n_878;
wire n_3457;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_1639;
wire n_1306;
wire n_3703;
wire n_1068;
wire n_3030;
wire n_3558;
wire n_1871;
wire n_2580;
wire n_3630;
wire n_2545;
wire n_2787;
wire n_3685;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_1163;
wire n_906;
wire n_3271;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_3753;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_3648;
wire n_2035;
wire n_2061;
wire n_3773;
wire n_3555;
wire n_3579;
wire n_3075;
wire n_3173;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_3236;
wire n_2398;
wire n_1362;
wire n_2857;
wire n_1586;
wire n_959;
wire n_2459;
wire n_3031;
wire n_3396;
wire n_3701;
wire n_940;
wire n_1445;
wire n_3516;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1923;
wire n_1773;
wire n_3243;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_2982;
wire n_3385;
wire n_1017;
wire n_2481;
wire n_2947;
wire n_3545;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_3343;
wire n_3515;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_1079;
wire n_1045;
wire n_2093;
wire n_2339;
wire n_2038;
wire n_2320;
wire n_2473;
wire n_1208;
wire n_3287;
wire n_2137;
wire n_3378;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_3767;
wire n_3426;
wire n_3454;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_3820;
wire n_3741;
wire n_3410;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_2029;
wire n_995;
wire n_3221;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_3629;
wire n_3021;
wire n_1989;
wire n_3818;
wire n_2359;
wire n_2941;
wire n_3674;
wire n_1887;
wire n_3502;
wire n_2523;
wire n_1383;
wire n_3098;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_2312;
wire n_962;
wire n_3475;
wire n_1215;
wire n_3015;
wire n_1171;
wire n_1578;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_3719;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_3681;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_3672;
wire n_2399;
wire n_3058;
wire n_2812;
wire n_2048;
wire n_3197;
wire n_3109;
wire n_3607;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_3505;
wire n_3002;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_3730;
wire n_1177;
wire n_3276;
wire n_1355;
wire n_2565;
wire n_974;
wire n_1159;
wire n_957;
wire n_3787;
wire n_2124;
wire n_3001;
wire n_2081;
wire n_3149;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_3268;
wire n_3597;
wire n_2418;
wire n_3827;
wire n_829;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_3614;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_3301;
wire n_3466;
wire n_3458;
wire n_1237;
wire n_1420;
wire n_3185;
wire n_1132;
wire n_3330;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_3248;
wire n_2277;
wire n_2477;
wire n_3523;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_1006;
wire n_3411;
wire n_2110;
wire n_3811;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_1486;
wire n_3586;
wire n_1332;
wire n_3519;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2879;
wire n_2474;
wire n_2604;
wire n_2090;
wire n_3374;
wire n_3153;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_3453;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_3399;
wire n_2896;
wire n_1111;
wire n_3213;
wire n_1365;
wire n_1927;
wire n_3065;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_3645;
wire n_1041;
wire n_1265;
wire n_3223;
wire n_1909;
wire n_3077;
wire n_2681;
wire n_1562;
wire n_3103;
wire n_834;
wire n_3474;
wire n_3675;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_3387;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_2878;
wire n_1823;
wire n_3679;
wire n_3779;
wire n_874;
wire n_2464;
wire n_3422;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_3557;
wire n_2230;
wire n_3498;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_3707;
wire n_987;
wire n_3189;
wire n_1846;
wire n_3037;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_3429;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_3154;
wire n_860;
wire n_3229;
wire n_2849;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_3692;
wire n_948;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_1849;
wire n_3788;
wire n_2410;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_2922;
wire n_1430;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2467;
wire n_3366;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_3421;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1044;
wire n_2436;
wire n_1205;
wire n_1209;
wire n_3029;
wire n_3242;
wire n_1552;
wire n_2508;
wire n_3592;
wire n_3618;
wire n_3525;
wire n_2593;
wire n_3486;
wire n_1435;
wire n_879;
wire n_3394;
wire n_3793;
wire n_3683;
wire n_2416;
wire n_2405;
wire n_3642;
wire n_3286;
wire n_2088;
wire n_2953;
wire n_3808;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_1684;
wire n_921;
wire n_996;
wire n_2658;
wire n_3590;
wire n_1717;
wire n_2895;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_3097;
wire n_3483;
wire n_1821;
wire n_2929;
wire n_3424;
wire n_3478;
wire n_1381;
wire n_2555;
wire n_3751;
wire n_2662;
wire n_2740;
wire n_3824;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_3388;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_3583;
wire n_2890;
wire n_3560;
wire n_3059;
wire n_3524;
wire n_2554;
wire n_3465;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_3215;
wire n_1438;
wire n_3698;
wire n_1082;
wire n_1840;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_3589;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_3171;
wire n_1229;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_3658;
wire n_3449;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_3559;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2989;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_3026;
wire n_2216;
wire n_3020;
wire n_3677;
wire n_1757;
wire n_890;
wire n_1897;
wire n_1919;
wire n_1424;
wire n_1056;
wire n_960;
wire n_3462;
wire n_3588;
wire n_2933;
wire n_2308;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_3419;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_3546;
wire n_1206;
wire n_2647;
wire n_3784;
wire n_3160;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_2969;
wire n_3195;
wire n_1519;
wire n_950;
wire n_3190;
wire n_2428;
wire n_1553;
wire n_3678;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_3456;
wire n_1346;
wire n_3053;
wire n_1299;
wire n_3244;
wire n_2158;
wire n_1808;
wire n_3290;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_3130;
wire n_2465;
wire n_2824;
wire n_3033;
wire n_2650;
wire n_3298;
wire n_3548;
wire n_912;
wire n_968;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_3334;
wire n_967;
wire n_1442;
wire n_2923;
wire n_3665;
wire n_3494;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_3264;
wire n_2333;
wire n_885;
wire n_2916;
wire n_3166;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_3771;
wire n_1632;
wire n_3110;
wire n_2998;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_3800;
wire n_2402;
wire n_1157;
wire n_3073;
wire n_2403;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_3162;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_3554;
wire n_3377;
wire n_2870;
wire n_3777;
wire n_1305;
wire n_3749;
wire n_3178;
wire n_873;
wire n_1826;
wire n_1112;
wire n_3134;
wire n_2304;
wire n_2999;
wire n_1644;
wire n_1283;
wire n_2334;
wire n_2637;
wire n_3695;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_3537;
wire n_2289;
wire n_3080;
wire n_3051;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_3362;
wire n_2881;
wire n_1631;
wire n_1203;
wire n_3750;
wire n_3282;
wire n_2472;
wire n_821;
wire n_3816;
wire n_1763;
wire n_2341;
wire n_3105;
wire n_3231;
wire n_1966;
wire n_3632;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_2993;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_3569;
wire n_2309;
wire n_2415;
wire n_2948;
wire n_3274;
wire n_3041;
wire n_3299;
wire n_2646;
wire n_1560;
wire n_3715;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_3209;
wire n_972;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_3040;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_3568;
wire n_3664;
wire n_2589;
wire n_3203;
wire n_1363;
wire n_1668;
wire n_1301;
wire n_3737;
wire n_1185;
wire n_991;
wire n_2903;
wire n_3417;
wire n_3482;
wire n_828;
wire n_1967;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_3717;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_3255;
wire n_1439;
wire n_1312;
wire n_804;
wire n_2827;
wire n_1688;
wire n_3052;
wire n_945;
wire n_2997;
wire n_3743;
wire n_3327;
wire n_1504;
wire n_943;
wire n_3326;
wire n_3572;
wire n_992;
wire n_3067;
wire n_1932;
wire n_3375;
wire n_2755;
wire n_842;
wire n_3734;
wire n_984;
wire n_3237;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_3167;
wire n_3400;
wire n_1594;
wire n_1400;
wire n_1342;
wire n_1214;
wire n_3423;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_3382;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3574;
wire n_918;
wire n_3529;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1977;
wire n_1557;
wire n_2153;
wire n_1147;
wire n_2468;
wire n_1610;
wire n_1422;
wire n_1077;
wire n_3196;
wire n_3078;
wire n_2364;
wire n_2533;
wire n_3492;
wire n_3094;
wire n_896;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2860;
wire n_3316;
wire n_2291;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_3253;
wire n_1730;
wire n_3601;
wire n_3603;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_3633;
wire n_3363;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_2973;
wire n_1470;
wire n_2094;
wire n_1096;
wire n_2670;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2318;
wire n_2393;
wire n_3689;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_3801;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_2974;
wire n_988;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_814;
wire n_2707;
wire n_2751;
wire n_2793;
wire n_3372;
wire n_3451;
wire n_2971;
wire n_3442;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_3240;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_3147;
wire n_2758;
wire n_1458;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1176;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_2559;
wire n_3230;
wire n_1020;
wire n_1062;
wire n_3342;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_3386;
wire n_3708;
wire n_1204;
wire n_2840;
wire n_3729;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_3488;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_3780;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_2893;
wire n_3636;
wire n_1188;
wire n_2588;
wire n_2962;
wire n_1722;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_2600;
wire n_849;
wire n_2795;
wire n_1638;
wire n_1786;
wire n_2981;
wire n_2002;
wire n_2282;
wire n_3608;
wire n_2800;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_3233;
wire n_3829;
wire n_3380;
wire n_3177;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_3409;
wire n_3460;
wire n_2352;
wire n_3538;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_3085;
wire n_2444;
wire n_2068;
wire n_3552;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_3123;
wire n_3684;
wire n_3137;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_939;
wire n_3697;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_789;
wire n_3393;
wire n_1603;
wire n_1232;
wire n_2638;
wire n_866;
wire n_1401;
wire n_969;
wire n_3520;
wire n_2492;
wire n_1998;
wire n_1019;
wire n_1105;
wire n_3759;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_2270;
wire n_1506;
wire n_3206;
wire n_2653;
wire n_3578;
wire n_836;
wire n_990;
wire n_2867;
wire n_3812;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_1465;
wire n_3145;
wire n_3124;
wire n_1122;
wire n_3192;
wire n_2608;
wire n_3764;
wire n_2657;
wire n_2995;
wire n_1375;
wire n_2494;
wire n_3547;
wire n_2649;
wire n_1102;
wire n_3727;
wire n_2852;
wire n_3774;
wire n_2392;
wire n_3459;
wire n_3093;
wire n_1843;
wire n_1499;
wire n_3061;
wire n_3155;
wire n_1187;
wire n_3517;
wire n_2633;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_3324;
wire n_3356;
wire n_3758;
wire n_2835;
wire n_2558;
wire n_1371;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_3803;
wire n_3182;
wire n_1572;
wire n_1968;
wire n_3742;
wire n_3269;
wire n_2564;
wire n_2252;
wire n_1516;
wire n_876;
wire n_3736;
wire n_1190;
wire n_3506;
wire n_1736;
wire n_3605;
wire n_1685;
wire n_2409;
wire n_917;
wire n_3450;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_3402;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_3565;
wire n_3174;
wire n_982;
wire n_2575;
wire n_2988;
wire n_3390;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_3746;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_2766;
wire n_3817;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2745;
wire n_2117;
wire n_2722;
wire n_3408;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_3432;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1345;
wire n_1059;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_3401;
wire n_1899;
wire n_3226;
wire n_1410;
wire n_1005;
wire n_1003;
wire n_3090;
wire n_2067;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_3762;
wire n_3533;
wire n_2877;
wire n_3318;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_3485;
wire n_1584;
wire n_1726;
wire n_1835;
wire n_3035;
wire n_3654;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_3333;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_3034;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_2811;
wire n_1496;
wire n_3348;
wire n_1125;
wire n_3014;
wire n_2547;
wire n_3639;
wire n_1812;
wire n_2501;
wire n_3079;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_3791;
wire n_3308;
wire n_2665;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_1533;
wire n_2224;
wire n_3368;
wire n_2924;
wire n_3467;
wire n_808;
wire n_2484;
wire n_797;
wire n_3530;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_3731;
wire n_2765;
wire n_3329;
wire n_2994;
wire n_1067;
wire n_3805;
wire n_3825;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_3135;
wire n_3657;
wire n_2003;
wire n_1457;
wire n_2692;
wire n_3573;
wire n_3148;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_3534;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_3757;
wire n_3438;
wire n_872;
wire n_2012;
wire n_3792;
wire n_1291;
wire n_3381;
wire n_3503;
wire n_1753;
wire n_1297;
wire n_2283;
wire n_2866;
wire n_3278;
wire n_1782;
wire n_2245;
wire n_3561;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_869;
wire n_810;
wire n_2965;
wire n_3536;
wire n_3661;
wire n_3635;
wire n_827;
wire n_3217;
wire n_3404;
wire n_3425;
wire n_1703;
wire n_3312;
wire n_1352;
wire n_2926;
wire n_2197;
wire n_2199;
wire n_3540;
wire n_1650;
wire n_3670;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_3046;
wire n_2213;
wire n_1170;
wire n_2023;
wire n_3826;
wire n_3249;
wire n_3211;
wire n_3285;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_2103;
wire n_2160;
wire n_3337;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_850;
wire n_3074;
wire n_3204;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_3673;
wire n_2480;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_3397;
wire n_3740;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_3005;
wire n_2332;
wire n_1235;
wire n_980;
wire n_1115;
wire n_2433;
wire n_3293;
wire n_3129;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_2977;
wire n_3606;
wire n_2601;
wire n_3043;
wire n_998;
wire n_3802;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_3600;
wire n_823;
wire n_2686;
wire n_2528;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_2316;
wire n_1985;
wire n_3055;
wire n_1898;
wire n_2107;
wire n_3294;
wire n_3219;
wire n_3711;
wire n_3315;
wire n_2906;
wire n_1625;
wire n_2130;
wire n_3415;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_3239;
wire n_3139;
wire n_2773;
wire n_3172;
wire n_3292;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_1452;
wire n_2687;
wire n_3023;
wire n_3553;
wire n_1120;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_2850;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_2654;
wire n_997;
wire n_3431;
wire n_3104;
wire n_932;
wire n_3169;
wire n_3151;
wire n_3822;
wire n_3131;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_3070;
wire n_3284;
wire n_3647;
wire n_3176;
wire n_2884;
wire n_1268;
wire n_2996;
wire n_825;
wire n_2819;
wire n_3126;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_1718;
wire n_3700;
wire n_3609;
wire n_986;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_3581;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_3576;
wire n_1063;
wire n_3720;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_1489;
wire n_1922;
wire n_2966;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_3495;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_2950;
wire n_792;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_3140;
wire n_3170;
wire n_3724;
wire n_812;
wire n_2104;
wire n_2748;
wire n_3311;
wire n_2057;
wire n_3272;
wire n_3011;
wire n_1772;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_3345;
wire n_862;
wire n_3584;
wire n_1425;
wire n_1901;
wire n_3069;
wire n_3756;
wire n_1900;
wire n_1620;
wire n_3032;
wire n_3628;
wire n_2889;
wire n_3691;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_3018;
wire n_1675;
wire n_3072;
wire n_1924;
wire n_2573;
wire n_3084;
wire n_3081;
wire n_3313;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_2939;
wire n_1745;
wire n_2735;
wire n_2497;
wire n_2006;
wire n_3412;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_3807;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_3761;
wire n_886;
wire n_3439;
wire n_2014;
wire n_3056;
wire n_1221;
wire n_2345;
wire n_2986;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_2774;
wire n_2726;
wire n_3295;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_2382;
wire n_1707;
wire n_853;
wire n_3062;
wire n_3161;
wire n_2317;
wire n_3289;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_3477;
wire n_3017;
wire n_3626;
wire n_2476;
wire n_787;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_2984;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_3364;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_930;
wire n_1873;
wire n_1411;
wire n_3201;
wire n_3054;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_3671;
wire n_1087;
wire n_3472;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_3344;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_3302;
wire n_3235;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_3391;
wire n_1567;
wire n_2567;
wire n_3543;
wire n_1247;
wire n_2709;
wire n_3102;
wire n_922;
wire n_3122;
wire n_816;
wire n_1648;
wire n_1536;
wire n_3050;
wire n_3265;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_3627;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_2957;
wire n_1769;
wire n_3551;
wire n_839;
wire n_1210;
wire n_3518;
wire n_2964;
wire n_3769;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_3733;
wire n_2183;
wire n_2742;
wire n_2673;
wire n_3314;
wire n_2360;
wire n_3254;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_3722;
wire n_1842;
wire n_871;
wire n_2442;
wire n_3309;
wire n_3738;
wire n_928;
wire n_1367;
wire n_1943;
wire n_3634;
wire n_1460;
wire n_2018;
wire n_3464;
wire n_3260;
wire n_1555;
wire n_3117;
wire n_2834;
wire n_3245;
wire n_3357;
wire n_2531;
wire n_1589;
wire n_3428;
wire n_2961;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_3351;
wire n_1619;
wire n_3527;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_3754;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_2883;
wire n_3115;
wire n_3509;
wire n_3352;
wire n_2208;
wire n_3076;
wire n_1404;
wire n_3063;
wire n_3617;
wire n_2912;
wire n_1794;
wire n_3535;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_3251;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_3118;
wire n_3227;
wire n_3300;
wire n_2321;
wire n_3511;
wire n_1226;
wire n_1277;
wire n_3680;
wire n_2591;
wire n_3443;
wire n_2146;
wire n_844;
wire n_3384;
wire n_852;
wire n_3497;
wire n_1487;
wire n_1864;
wire n_3644;
wire n_1601;
wire n_1028;
wire n_3336;
wire n_2940;
wire n_3435;
wire n_3521;
wire n_3575;
wire n_1546;
wire n_3562;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_979;
wire n_1515;
wire n_2841;
wire n_3165;
wire n_1627;
wire n_2918;
wire n_3232;
wire n_3322;
wire n_3652;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_2832;
wire n_1975;
wire n_1321;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_3250;
wire n_1739;
wire n_3181;
wire n_2958;
wire n_2278;
wire n_2594;
wire n_3114;
wire n_3125;
wire n_2394;
wire n_3234;
wire n_1914;
wire n_3612;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_3493;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_3004;
wire n_3323;
wire n_2569;
wire n_3112;
wire n_2349;
wire n_1103;
wire n_3132;
wire n_3556;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_3591;
wire n_3024;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_3512;
wire n_1761;
wire n_3238;
wire n_3210;
wire n_3175;
wire n_3522;
wire n_2036;
wire n_1325;
wire n_3267;
wire n_1595;
wire n_2161;
wire n_795;
wire n_2404;
wire n_2083;
wire n_3281;
wire n_3307;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_3266;
wire n_2485;
wire n_3772;
wire n_1956;
wire n_1936;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_2655;
wire n_2027;
wire n_2642;
wire n_1130;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_3726;
wire n_2210;
wire n_805;
wire n_3247;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_3091;
wire n_2695;
wire n_1764;
wire n_3480;
wire n_2892;
wire n_3057;
wire n_3194;
wire n_3582;
wire n_3066;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_3577;
wire n_3539;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_3662;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_3347;
wire n_2004;
wire n_3216;
wire n_1621;
wire n_2708;
wire n_3809;
wire n_2113;
wire n_2586;
wire n_3694;
wire n_1448;
wire n_2225;
wire n_3567;
wire n_3613;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_3444;
wire n_1505;
wire n_1181;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_1340;
wire n_2274;
wire n_2972;
wire n_811;
wire n_3225;
wire n_1558;
wire n_807;
wire n_3321;
wire n_2166;
wire n_2938;
wire n_3212;
wire n_835;
wire n_3319;
wire n_1433;
wire n_3594;
wire n_1704;
wire n_2256;
wire n_3152;
wire n_3721;
wire n_3335;
wire n_1254;
wire n_3799;
wire n_1026;
wire n_3413;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_2044;
wire n_1089;
wire n_2013;
wire n_927;
wire n_1138;
wire n_1990;
wire n_2689;
wire n_2920;
wire n_3259;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_2991;
wire n_3688;
wire n_3383;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_3016;
wire n_1693;
wire n_3585;
wire n_2975;
wire n_3473;
wire n_2599;
wire n_2704;
wire n_904;
wire n_2839;
wire n_3338;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_3414;
wire n_3463;
wire n_3699;
wire n_1827;
wire n_1180;
wire n_3360;
wire n_2524;
wire n_1271;
wire n_3705;
wire n_2802;
wire n_1542;
wire n_1251;
wire n_3693;
wire n_3159;
wire n_2728;
wire n_2268;
wire n_3778;

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_96),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_754),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_636),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_376),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_632),
.Y(n_791)
);

BUFx10_ASAP7_75t_L g792 ( 
.A(n_204),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_681),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_698),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_253),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_634),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_289),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_59),
.Y(n_798)
);

INVx1_ASAP7_75t_SL g799 ( 
.A(n_449),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_132),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_519),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_439),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_202),
.Y(n_803)
);

INVx1_ASAP7_75t_SL g804 ( 
.A(n_123),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_204),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_624),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_745),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_537),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_383),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_560),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_427),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_576),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_481),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_779),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_386),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_519),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_91),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_414),
.Y(n_818)
);

INVxp33_ASAP7_75t_L g819 ( 
.A(n_457),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_290),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_773),
.Y(n_821)
);

INVx1_ASAP7_75t_SL g822 ( 
.A(n_542),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_589),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_605),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_539),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_758),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_782),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_314),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_255),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_596),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_772),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_412),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_144),
.Y(n_833)
);

CKINVDCx14_ASAP7_75t_R g834 ( 
.A(n_115),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_753),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_239),
.Y(n_836)
);

BUFx10_ASAP7_75t_L g837 ( 
.A(n_703),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_689),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_771),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_152),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_18),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_647),
.Y(n_842)
);

CKINVDCx20_ASAP7_75t_R g843 ( 
.A(n_701),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_209),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_395),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_293),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_323),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_513),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_505),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_377),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_16),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_266),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_436),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_526),
.Y(n_854)
);

CKINVDCx16_ASAP7_75t_R g855 ( 
.A(n_309),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_677),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_620),
.Y(n_857)
);

INVx1_ASAP7_75t_SL g858 ( 
.A(n_770),
.Y(n_858)
);

CKINVDCx11_ASAP7_75t_R g859 ( 
.A(n_118),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_517),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_500),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_285),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_348),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_685),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_10),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_358),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_184),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_736),
.Y(n_868)
);

CKINVDCx16_ASAP7_75t_R g869 ( 
.A(n_469),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_540),
.Y(n_870)
);

BUFx3_ASAP7_75t_L g871 ( 
.A(n_355),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_374),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_640),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_651),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_126),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_185),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_303),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_95),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_31),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_9),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_444),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_8),
.Y(n_882)
);

CKINVDCx16_ASAP7_75t_R g883 ( 
.A(n_149),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_275),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_746),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_344),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_710),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_315),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_622),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_431),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_487),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_643),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_227),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_130),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_96),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_149),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_750),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_178),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_609),
.Y(n_899)
);

BUFx10_ASAP7_75t_L g900 ( 
.A(n_99),
.Y(n_900)
);

INVxp33_ASAP7_75t_SL g901 ( 
.A(n_504),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_436),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_275),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_310),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_192),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_299),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_49),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_459),
.Y(n_908)
);

INVxp33_ASAP7_75t_SL g909 ( 
.A(n_26),
.Y(n_909)
);

CKINVDCx20_ASAP7_75t_R g910 ( 
.A(n_508),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_672),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_705),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_29),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_521),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_539),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_358),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_7),
.Y(n_917)
);

BUFx8_ASAP7_75t_SL g918 ( 
.A(n_715),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_476),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_518),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_662),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_402),
.Y(n_922)
);

BUFx3_ASAP7_75t_L g923 ( 
.A(n_341),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_36),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_392),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_509),
.Y(n_926)
);

BUFx10_ASAP7_75t_L g927 ( 
.A(n_508),
.Y(n_927)
);

BUFx5_ASAP7_75t_L g928 ( 
.A(n_255),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_497),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_39),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_291),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_3),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_402),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_367),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_297),
.Y(n_935)
);

INVxp67_ASAP7_75t_L g936 ( 
.A(n_530),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_90),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_475),
.Y(n_938)
);

CKINVDCx16_ASAP7_75t_R g939 ( 
.A(n_470),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_777),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_99),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_764),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_757),
.Y(n_943)
);

CKINVDCx14_ASAP7_75t_R g944 ( 
.A(n_451),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_769),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_603),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_540),
.Y(n_947)
);

CKINVDCx20_ASAP7_75t_R g948 ( 
.A(n_721),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_679),
.Y(n_949)
);

INVx1_ASAP7_75t_SL g950 ( 
.A(n_385),
.Y(n_950)
);

CKINVDCx20_ASAP7_75t_R g951 ( 
.A(n_365),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_140),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_2),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_106),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_107),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_439),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_472),
.Y(n_957)
);

CKINVDCx14_ASAP7_75t_R g958 ( 
.A(n_162),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_728),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_727),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_212),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_283),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_355),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_502),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_712),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_494),
.Y(n_966)
);

BUFx10_ASAP7_75t_L g967 ( 
.A(n_403),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_94),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_776),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_47),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_324),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_230),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_756),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_175),
.Y(n_974)
);

BUFx3_ASAP7_75t_L g975 ( 
.A(n_183),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_543),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_138),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_627),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_347),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_617),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_36),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_780),
.Y(n_982)
);

BUFx5_ASAP7_75t_L g983 ( 
.A(n_762),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_719),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_263),
.Y(n_985)
);

CKINVDCx20_ASAP7_75t_R g986 ( 
.A(n_166),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_646),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_17),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_197),
.Y(n_989)
);

CKINVDCx16_ASAP7_75t_R g990 ( 
.A(n_512),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_676),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_234),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_562),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_470),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_156),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_239),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_350),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_33),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_763),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_612),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_579),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_500),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_648),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_56),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_143),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_546),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_495),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_228),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_222),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_235),
.Y(n_1010)
);

BUFx8_ASAP7_75t_SL g1011 ( 
.A(n_137),
.Y(n_1011)
);

INVx1_ASAP7_75t_SL g1012 ( 
.A(n_289),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_337),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_25),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_70),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_62),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_248),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_718),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_11),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_475),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_248),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_709),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_170),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_13),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_172),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_644),
.Y(n_1026)
);

INVx2_ASAP7_75t_SL g1027 ( 
.A(n_422),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_244),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_254),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_456),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_559),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_120),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_574),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_140),
.Y(n_1034)
);

BUFx5_ASAP7_75t_L g1035 ( 
.A(n_550),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_319),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_435),
.Y(n_1037)
);

CKINVDCx16_ASAP7_75t_R g1038 ( 
.A(n_378),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_SL g1039 ( 
.A(n_187),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_70),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_532),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_541),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_557),
.Y(n_1043)
);

BUFx10_ASAP7_75t_L g1044 ( 
.A(n_449),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_488),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_378),
.Y(n_1046)
);

INVx2_ASAP7_75t_SL g1047 ( 
.A(n_546),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_329),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_734),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_238),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_503),
.Y(n_1051)
);

INVx1_ASAP7_75t_SL g1052 ( 
.A(n_699),
.Y(n_1052)
);

CKINVDCx20_ASAP7_75t_R g1053 ( 
.A(n_524),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_348),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_761),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_731),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_748),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_380),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_306),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_510),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_460),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_571),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_366),
.Y(n_1063)
);

INVx1_ASAP7_75t_SL g1064 ( 
.A(n_254),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_495),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_732),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_125),
.Y(n_1067)
);

CKINVDCx20_ASAP7_75t_R g1068 ( 
.A(n_308),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_428),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_213),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_536),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_184),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_103),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_607),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_11),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_545),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_53),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_92),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_578),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_590),
.Y(n_1080)
);

BUFx5_ASAP7_75t_L g1081 ( 
.A(n_446),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_552),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_464),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_236),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_327),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_584),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_434),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_175),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_440),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_244),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_455),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_453),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_437),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_95),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_231),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_463),
.Y(n_1096)
);

INVx1_ASAP7_75t_SL g1097 ( 
.A(n_257),
.Y(n_1097)
);

CKINVDCx20_ASAP7_75t_R g1098 ( 
.A(n_641),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_240),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_541),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_116),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_269),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_131),
.Y(n_1103)
);

CKINVDCx16_ASAP7_75t_R g1104 ( 
.A(n_191),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_498),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_4),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_469),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_148),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_544),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_558),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_467),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_165),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_464),
.Y(n_1113)
);

CKINVDCx20_ASAP7_75t_R g1114 ( 
.A(n_784),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_714),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_525),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_205),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_344),
.Y(n_1118)
);

BUFx2_ASAP7_75t_L g1119 ( 
.A(n_85),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_534),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_713),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_509),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_555),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_507),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_215),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_536),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_225),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_89),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_173),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_538),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_435),
.Y(n_1131)
);

INVx2_ASAP7_75t_SL g1132 ( 
.A(n_177),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_260),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_430),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_395),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_249),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_362),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_100),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_549),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_529),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_616),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_535),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_373),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_18),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_273),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_194),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_522),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_768),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_633),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_391),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_370),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_410),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_502),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_447),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_226),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_760),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_128),
.Y(n_1157)
);

CKINVDCx20_ASAP7_75t_R g1158 ( 
.A(n_499),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_133),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_708),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_61),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_515),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_160),
.Y(n_1163)
);

CKINVDCx14_ASAP7_75t_R g1164 ( 
.A(n_141),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_682),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_528),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_53),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_265),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_586),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_68),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_479),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_687),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_691),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_285),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_90),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_45),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_333),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_87),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_205),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_485),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_245),
.Y(n_1181)
);

CKINVDCx20_ASAP7_75t_R g1182 ( 
.A(n_3),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_477),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_626),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_251),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_27),
.Y(n_1186)
);

INVxp67_ASAP7_75t_L g1187 ( 
.A(n_343),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_207),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_9),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_30),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_514),
.Y(n_1191)
);

CKINVDCx20_ASAP7_75t_R g1192 ( 
.A(n_210),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_241),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_716),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_44),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_767),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_774),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_755),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_31),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_128),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_511),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_197),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_720),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_506),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_10),
.Y(n_1206)
);

INVx1_ASAP7_75t_SL g1207 ( 
.A(n_236),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_60),
.Y(n_1208)
);

BUFx2_ASAP7_75t_L g1209 ( 
.A(n_142),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_330),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_42),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_174),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_501),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_591),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_249),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_220),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_447),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_247),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_485),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_751),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_446),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_361),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_110),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_63),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_775),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_441),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_364),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_637),
.Y(n_1228)
);

INVx1_ASAP7_75t_SL g1229 ( 
.A(n_23),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_749),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_383),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_270),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_115),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_303),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_198),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_59),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_357),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_352),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_530),
.Y(n_1239)
);

BUFx10_ASAP7_75t_L g1240 ( 
.A(n_12),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_330),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_126),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_212),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_759),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_533),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_207),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_157),
.Y(n_1247)
);

BUFx10_ASAP7_75t_L g1248 ( 
.A(n_361),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_572),
.Y(n_1249)
);

CKINVDCx16_ASAP7_75t_R g1250 ( 
.A(n_538),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_392),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_510),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_523),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_35),
.Y(n_1254)
);

BUFx10_ASAP7_75t_L g1255 ( 
.A(n_497),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_664),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_700),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_296),
.Y(n_1258)
);

INVx1_ASAP7_75t_SL g1259 ( 
.A(n_258),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_328),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_737),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_531),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_336),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_404),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_729),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_387),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_253),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_693),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_63),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_663),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_785),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_103),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_725),
.Y(n_1273)
);

INVx1_ASAP7_75t_SL g1274 ( 
.A(n_730),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_49),
.Y(n_1275)
);

INVx1_ASAP7_75t_SL g1276 ( 
.A(n_752),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_511),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_766),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_91),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_527),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_688),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_629),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_286),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_744),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_516),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_747),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_176),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_405),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_608),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_178),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_434),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_166),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_397),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_489),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_93),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_765),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_575),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_214),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_577),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_327),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_8),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_597),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_403),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_738),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_411),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_92),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_87),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_241),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_551),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_442),
.Y(n_1310)
);

INVx1_ASAP7_75t_SL g1311 ( 
.A(n_267),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_413),
.Y(n_1312)
);

INVx2_ASAP7_75t_SL g1313 ( 
.A(n_110),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_496),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_783),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_363),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_213),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_273),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_520),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_601),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_1),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_454),
.Y(n_1322)
);

CKINVDCx14_ASAP7_75t_R g1323 ( 
.A(n_450),
.Y(n_1323)
);

INVxp33_ASAP7_75t_SL g1324 ( 
.A(n_997),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_928),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_928),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_862),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_928),
.Y(n_1328)
);

INVxp67_ASAP7_75t_SL g1329 ( 
.A(n_862),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_928),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_859),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_859),
.Y(n_1332)
);

CKINVDCx20_ASAP7_75t_R g1333 ( 
.A(n_948),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_819),
.B(n_0),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_1284),
.Y(n_1335)
);

CKINVDCx16_ASAP7_75t_R g1336 ( 
.A(n_855),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_928),
.Y(n_1337)
);

CKINVDCx16_ASAP7_75t_R g1338 ( 
.A(n_869),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_928),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_928),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1081),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1081),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_1011),
.Y(n_1343)
);

INVxp33_ASAP7_75t_L g1344 ( 
.A(n_1040),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1081),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1081),
.Y(n_1346)
);

CKINVDCx20_ASAP7_75t_R g1347 ( 
.A(n_843),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_1011),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1081),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1081),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1081),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_828),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_828),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_862),
.Y(n_1354)
);

INVxp67_ASAP7_75t_SL g1355 ( 
.A(n_862),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_871),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_871),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_923),
.Y(n_1358)
);

INVxp33_ASAP7_75t_L g1359 ( 
.A(n_1157),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_788),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_923),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_935),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_935),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_789),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_994),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_975),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_975),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_976),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_976),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_998),
.Y(n_1370)
);

INVxp33_ASAP7_75t_L g1371 ( 
.A(n_1288),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_998),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_843),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1060),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_994),
.Y(n_1375)
);

INVxp67_ASAP7_75t_SL g1376 ( 
.A(n_994),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1060),
.Y(n_1377)
);

INVxp33_ASAP7_75t_SL g1378 ( 
.A(n_1021),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_994),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1016),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1016),
.Y(n_1381)
);

CKINVDCx20_ASAP7_75t_R g1382 ( 
.A(n_1066),
.Y(n_1382)
);

INVxp67_ASAP7_75t_SL g1383 ( 
.A(n_1016),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_814),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1016),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1106),
.Y(n_1386)
);

CKINVDCx20_ASAP7_75t_R g1387 ( 
.A(n_1066),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1106),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1106),
.Y(n_1389)
);

CKINVDCx16_ASAP7_75t_R g1390 ( 
.A(n_883),
.Y(n_1390)
);

INVx1_ASAP7_75t_SL g1391 ( 
.A(n_1023),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1106),
.Y(n_1392)
);

CKINVDCx16_ASAP7_75t_R g1393 ( 
.A(n_939),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_821),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1133),
.Y(n_1395)
);

CKINVDCx20_ASAP7_75t_R g1396 ( 
.A(n_1080),
.Y(n_1396)
);

INVxp67_ASAP7_75t_L g1397 ( 
.A(n_1045),
.Y(n_1397)
);

INVxp67_ASAP7_75t_SL g1398 ( 
.A(n_1133),
.Y(n_1398)
);

INVxp67_ASAP7_75t_SL g1399 ( 
.A(n_1133),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1133),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_792),
.Y(n_1401)
);

INVxp33_ASAP7_75t_SL g1402 ( 
.A(n_1069),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1171),
.Y(n_1403)
);

INVx4_ASAP7_75t_R g1404 ( 
.A(n_1039),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1171),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1171),
.Y(n_1406)
);

INVxp67_ASAP7_75t_SL g1407 ( 
.A(n_1171),
.Y(n_1407)
);

INVxp33_ASAP7_75t_SL g1408 ( 
.A(n_1119),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_790),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_797),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_802),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_808),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_844),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_846),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_983),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_847),
.Y(n_1416)
);

INVxp67_ASAP7_75t_SL g1417 ( 
.A(n_800),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_851),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_853),
.Y(n_1419)
);

INVxp67_ASAP7_75t_SL g1420 ( 
.A(n_800),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_861),
.Y(n_1421)
);

INVxp67_ASAP7_75t_SL g1422 ( 
.A(n_836),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_824),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_863),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_867),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_870),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_880),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_881),
.Y(n_1428)
);

INVxp33_ASAP7_75t_SL g1429 ( 
.A(n_1209),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_890),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_898),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_903),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_983),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_904),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_983),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_907),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_919),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_925),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_836),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_931),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_983),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_826),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_932),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_953),
.Y(n_1444)
);

INVx1_ASAP7_75t_SL g1445 ( 
.A(n_910),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_954),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_794),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_964),
.Y(n_1448)
);

INVxp67_ASAP7_75t_SL g1449 ( 
.A(n_879),
.Y(n_1449)
);

CKINVDCx20_ASAP7_75t_R g1450 ( 
.A(n_1080),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_974),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_816),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_879),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_981),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_983),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_983),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_988),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_983),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_989),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_966),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_992),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1006),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1331),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1354),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1329),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1360),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1447),
.B(n_834),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1365),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1329),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_L g1470 ( 
.A(n_1375),
.Y(n_1470)
);

INVx5_ASAP7_75t_L g1471 ( 
.A(n_1327),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1364),
.B(n_823),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1405),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1384),
.B(n_834),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1332),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1355),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1378),
.A2(n_944),
.B1(n_1164),
.B2(n_958),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1327),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1394),
.B(n_944),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1379),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1355),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1376),
.B(n_1184),
.Y(n_1482)
);

BUFx6f_ASAP7_75t_L g1483 ( 
.A(n_1380),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1423),
.B(n_1281),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1442),
.B(n_1086),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1376),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1383),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1344),
.B(n_958),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1381),
.Y(n_1489)
);

BUFx6f_ASAP7_75t_L g1490 ( 
.A(n_1385),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1352),
.Y(n_1491)
);

AOI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1402),
.A2(n_1323),
.B1(n_1164),
.B2(n_909),
.Y(n_1492)
);

BUFx12f_ASAP7_75t_L g1493 ( 
.A(n_1343),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1386),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1324),
.B(n_1323),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1383),
.B(n_794),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1398),
.Y(n_1497)
);

INVxp67_ASAP7_75t_L g1498 ( 
.A(n_1401),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1353),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1388),
.Y(n_1500)
);

OA21x2_ASAP7_75t_L g1501 ( 
.A1(n_1325),
.A2(n_965),
.B(n_887),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1389),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1392),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1326),
.A2(n_965),
.B(n_887),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1398),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1391),
.B(n_990),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1408),
.A2(n_901),
.B1(n_1104),
.B2(n_1038),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1359),
.B(n_1250),
.Y(n_1508)
);

AND2x6_ASAP7_75t_L g1509 ( 
.A(n_1328),
.B(n_793),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1395),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1415),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1399),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1400),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1399),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1407),
.Y(n_1515)
);

BUFx12f_ASAP7_75t_L g1516 ( 
.A(n_1348),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1403),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1407),
.Y(n_1518)
);

INVx4_ASAP7_75t_L g1519 ( 
.A(n_1433),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1406),
.Y(n_1520)
);

AOI22x1_ASAP7_75t_SL g1521 ( 
.A1(n_1347),
.A2(n_795),
.B1(n_840),
.B2(n_833),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1330),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1397),
.B(n_946),
.Y(n_1523)
);

BUFx6f_ASAP7_75t_L g1524 ( 
.A(n_1337),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1417),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1339),
.A2(n_1001),
.B(n_969),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1397),
.B(n_946),
.Y(n_1527)
);

BUFx3_ASAP7_75t_L g1528 ( 
.A(n_1356),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1357),
.B(n_1172),
.Y(n_1529)
);

BUFx6f_ASAP7_75t_L g1530 ( 
.A(n_1340),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1333),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1358),
.B(n_1172),
.Y(n_1532)
);

OA21x2_ASAP7_75t_L g1533 ( 
.A1(n_1341),
.A2(n_1001),
.B(n_969),
.Y(n_1533)
);

BUFx6f_ASAP7_75t_L g1534 ( 
.A(n_1342),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1361),
.B(n_1362),
.Y(n_1535)
);

INVx5_ASAP7_75t_L g1536 ( 
.A(n_1336),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1363),
.B(n_1249),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1345),
.Y(n_1538)
);

OA21x2_ASAP7_75t_L g1539 ( 
.A1(n_1346),
.A2(n_1249),
.B(n_796),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1349),
.Y(n_1540)
);

AND2x2_ASAP7_75t_SL g1541 ( 
.A(n_1338),
.B(n_906),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1359),
.B(n_1371),
.Y(n_1542)
);

BUFx6f_ASAP7_75t_L g1543 ( 
.A(n_1350),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1366),
.B(n_1367),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1351),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1417),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1409),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1368),
.B(n_791),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1429),
.B(n_819),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1369),
.B(n_806),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1410),
.Y(n_1551)
);

BUFx6f_ASAP7_75t_L g1552 ( 
.A(n_1411),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1370),
.Y(n_1553)
);

BUFx6f_ASAP7_75t_L g1554 ( 
.A(n_1412),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1413),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1372),
.B(n_807),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1414),
.Y(n_1557)
);

BUFx3_ASAP7_75t_L g1558 ( 
.A(n_1374),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1335),
.Y(n_1559)
);

BUFx3_ASAP7_75t_L g1560 ( 
.A(n_1377),
.Y(n_1560)
);

AOI22xp5_ASAP7_75t_SL g1561 ( 
.A1(n_1373),
.A2(n_795),
.B1(n_840),
.B2(n_833),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1416),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1390),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1420),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1418),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_L g1566 ( 
.A(n_1419),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1420),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1422),
.B(n_810),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1452),
.B(n_812),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1422),
.Y(n_1570)
);

OAI21x1_ASAP7_75t_L g1571 ( 
.A1(n_1435),
.A2(n_838),
.B(n_830),
.Y(n_1571)
);

OAI21x1_ASAP7_75t_L g1572 ( 
.A1(n_1441),
.A2(n_874),
.B(n_856),
.Y(n_1572)
);

AOI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1393),
.A2(n_1114),
.B1(n_1244),
.B2(n_1098),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1449),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1421),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1382),
.Y(n_1576)
);

BUFx6f_ASAP7_75t_L g1577 ( 
.A(n_1424),
.Y(n_1577)
);

INVx3_ASAP7_75t_L g1578 ( 
.A(n_1425),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1449),
.Y(n_1579)
);

BUFx6f_ASAP7_75t_L g1580 ( 
.A(n_1426),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1427),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1428),
.Y(n_1582)
);

OA21x2_ASAP7_75t_L g1583 ( 
.A1(n_1455),
.A2(n_892),
.B(n_889),
.Y(n_1583)
);

OA21x2_ASAP7_75t_L g1584 ( 
.A1(n_1456),
.A2(n_943),
.B(n_921),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1371),
.B(n_837),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1387),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1439),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1452),
.B(n_837),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1470),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1470),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1542),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1545),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1496),
.B(n_1430),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1488),
.B(n_1460),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1465),
.B(n_1334),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1545),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1524),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_1470),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1524),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1524),
.Y(n_1600)
);

INVxp67_ASAP7_75t_L g1601 ( 
.A(n_1506),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1563),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1530),
.Y(n_1603)
);

BUFx3_ASAP7_75t_L g1604 ( 
.A(n_1465),
.Y(n_1604)
);

NAND2xp33_ASAP7_75t_L g1605 ( 
.A(n_1484),
.B(n_1474),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1530),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1483),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1530),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1534),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1483),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1483),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1490),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1522),
.B(n_1458),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1496),
.B(n_1431),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1534),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1534),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1538),
.Y(n_1617)
);

BUFx8_ASAP7_75t_L g1618 ( 
.A(n_1586),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1541),
.B(n_793),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1538),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1538),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1490),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1543),
.Y(n_1623)
);

BUFx2_ASAP7_75t_L g1624 ( 
.A(n_1508),
.Y(n_1624)
);

BUFx6f_ASAP7_75t_L g1625 ( 
.A(n_1543),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1525),
.B(n_1432),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1467),
.Y(n_1627)
);

INVx3_ASAP7_75t_L g1628 ( 
.A(n_1490),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1510),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1543),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1469),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1469),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1497),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1497),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1510),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1540),
.B(n_1035),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1512),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1511),
.B(n_1035),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1510),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1513),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1512),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1585),
.B(n_1460),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1513),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1476),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1513),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1546),
.B(n_1434),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1481),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1486),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1564),
.B(n_1436),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1588),
.B(n_1445),
.Y(n_1650)
);

NAND2xp33_ASAP7_75t_SL g1651 ( 
.A(n_1477),
.B(n_1098),
.Y(n_1651)
);

BUFx6f_ASAP7_75t_L g1652 ( 
.A(n_1517),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1517),
.Y(n_1653)
);

BUFx2_ASAP7_75t_L g1654 ( 
.A(n_1498),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1487),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1505),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1517),
.Y(n_1657)
);

BUFx6f_ASAP7_75t_L g1658 ( 
.A(n_1571),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1514),
.Y(n_1659)
);

INVx3_ASAP7_75t_L g1660 ( 
.A(n_1511),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1549),
.B(n_1439),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1515),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1464),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1518),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1519),
.B(n_1035),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1491),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1468),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1495),
.B(n_1114),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1473),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1480),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1482),
.Y(n_1671)
);

INVx3_ASAP7_75t_L g1672 ( 
.A(n_1519),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1466),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1489),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1501),
.B(n_1035),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1499),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1528),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1553),
.Y(n_1678)
);

INVx3_ASAP7_75t_L g1679 ( 
.A(n_1552),
.Y(n_1679)
);

BUFx6f_ASAP7_75t_L g1680 ( 
.A(n_1572),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1558),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1560),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1482),
.Y(n_1683)
);

BUFx3_ASAP7_75t_L g1684 ( 
.A(n_1544),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1494),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1500),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1555),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1555),
.Y(n_1688)
);

BUFx6f_ASAP7_75t_L g1689 ( 
.A(n_1552),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1552),
.Y(n_1690)
);

BUFx6f_ASAP7_75t_L g1691 ( 
.A(n_1554),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1554),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1554),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1557),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1557),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1567),
.B(n_1334),
.Y(n_1696)
);

BUFx6f_ASAP7_75t_L g1697 ( 
.A(n_1557),
.Y(n_1697)
);

INVx3_ASAP7_75t_L g1698 ( 
.A(n_1566),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1566),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1566),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1577),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1577),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1577),
.Y(n_1703)
);

AND3x1_ASAP7_75t_L g1704 ( 
.A(n_1507),
.B(n_1047),
.C(n_1027),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1502),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1580),
.Y(n_1706)
);

INVxp67_ASAP7_75t_L g1707 ( 
.A(n_1587),
.Y(n_1707)
);

INVx3_ASAP7_75t_L g1708 ( 
.A(n_1580),
.Y(n_1708)
);

AND3x1_ASAP7_75t_L g1709 ( 
.A(n_1492),
.B(n_1132),
.C(n_1117),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1479),
.B(n_1453),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_SL g1711 ( 
.A(n_1570),
.B(n_793),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1574),
.B(n_1453),
.Y(n_1712)
);

INVx3_ASAP7_75t_L g1713 ( 
.A(n_1580),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1551),
.Y(n_1714)
);

INVxp67_ASAP7_75t_L g1715 ( 
.A(n_1472),
.Y(n_1715)
);

BUFx8_ASAP7_75t_L g1716 ( 
.A(n_1463),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_SL g1717 ( 
.A(n_1536),
.B(n_1244),
.Y(n_1717)
);

BUFx2_ASAP7_75t_L g1718 ( 
.A(n_1573),
.Y(n_1718)
);

INVx1_ASAP7_75t_SL g1719 ( 
.A(n_1576),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1503),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1562),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1478),
.Y(n_1722)
);

XNOR2xp5_ASAP7_75t_L g1723 ( 
.A(n_1531),
.B(n_1396),
.Y(n_1723)
);

INVx4_ASAP7_75t_L g1724 ( 
.A(n_1539),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1520),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1565),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1687),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1642),
.B(n_1536),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_SL g1729 ( 
.A1(n_1718),
.A2(n_1450),
.B1(n_1561),
.B2(n_1521),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1684),
.Y(n_1730)
);

INVx4_ASAP7_75t_L g1731 ( 
.A(n_1689),
.Y(n_1731)
);

AND2x6_ASAP7_75t_L g1732 ( 
.A(n_1675),
.B(n_1523),
.Y(n_1732)
);

NOR2x1p5_ASAP7_75t_L g1733 ( 
.A(n_1673),
.B(n_1493),
.Y(n_1733)
);

OAI22xp5_ASAP7_75t_L g1734 ( 
.A1(n_1715),
.A2(n_1683),
.B1(n_1671),
.B2(n_1601),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1688),
.Y(n_1735)
);

BUFx6f_ASAP7_75t_L g1736 ( 
.A(n_1689),
.Y(n_1736)
);

AND2x6_ASAP7_75t_L g1737 ( 
.A(n_1675),
.B(n_1595),
.Y(n_1737)
);

AND2x6_ASAP7_75t_L g1738 ( 
.A(n_1595),
.B(n_1523),
.Y(n_1738)
);

AND2x6_ASAP7_75t_L g1739 ( 
.A(n_1650),
.B(n_1527),
.Y(n_1739)
);

INVx2_ASAP7_75t_SL g1740 ( 
.A(n_1712),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1591),
.B(n_1475),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1631),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1632),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1633),
.Y(n_1744)
);

INVx4_ASAP7_75t_L g1745 ( 
.A(n_1689),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_SL g1746 ( 
.A(n_1671),
.B(n_1536),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1634),
.Y(n_1747)
);

BUFx10_ASAP7_75t_L g1748 ( 
.A(n_1696),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_SL g1749 ( 
.A(n_1683),
.B(n_1485),
.Y(n_1749)
);

INVx4_ASAP7_75t_SL g1750 ( 
.A(n_1710),
.Y(n_1750)
);

INVx1_ASAP7_75t_SL g1751 ( 
.A(n_1654),
.Y(n_1751)
);

AOI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1605),
.A2(n_1579),
.B1(n_1548),
.B2(n_1568),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_L g1753 ( 
.A1(n_1696),
.A2(n_1539),
.B1(n_1584),
.B2(n_1583),
.Y(n_1753)
);

OAI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1715),
.A2(n_1052),
.B1(n_1256),
.B2(n_858),
.Y(n_1754)
);

INVx5_ASAP7_75t_L g1755 ( 
.A(n_1625),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1663),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1667),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_SL g1758 ( 
.A(n_1601),
.B(n_1527),
.Y(n_1758)
);

BUFx8_ASAP7_75t_SL g1759 ( 
.A(n_1602),
.Y(n_1759)
);

INVxp33_ASAP7_75t_L g1760 ( 
.A(n_1723),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_SL g1761 ( 
.A(n_1593),
.B(n_1529),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1591),
.B(n_1559),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1669),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1707),
.B(n_1516),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1637),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1619),
.A2(n_1548),
.B1(n_1276),
.B2(n_1274),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1641),
.Y(n_1767)
);

INVx3_ASAP7_75t_L g1768 ( 
.A(n_1691),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1660),
.B(n_1583),
.Y(n_1769)
);

INVxp67_ASAP7_75t_SL g1770 ( 
.A(n_1660),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1672),
.B(n_1584),
.Y(n_1771)
);

BUFx6f_ASAP7_75t_L g1772 ( 
.A(n_1691),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1661),
.B(n_1529),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_SL g1774 ( 
.A(n_1719),
.B(n_918),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1670),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1674),
.Y(n_1776)
);

NAND3xp33_ASAP7_75t_L g1777 ( 
.A(n_1707),
.B(n_1556),
.C(n_1550),
.Y(n_1777)
);

AND2x4_ASAP7_75t_L g1778 ( 
.A(n_1593),
.B(n_1544),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_1719),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1644),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1647),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1685),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1594),
.B(n_1532),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1686),
.Y(n_1784)
);

AND2x6_ASAP7_75t_L g1785 ( 
.A(n_1658),
.B(n_793),
.Y(n_1785)
);

AOI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1619),
.A2(n_1532),
.B1(n_831),
.B2(n_835),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1648),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1655),
.Y(n_1788)
);

INVx4_ASAP7_75t_L g1789 ( 
.A(n_1691),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1672),
.B(n_1501),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1705),
.Y(n_1791)
);

BUFx3_ASAP7_75t_L g1792 ( 
.A(n_1618),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1656),
.Y(n_1793)
);

BUFx3_ASAP7_75t_L g1794 ( 
.A(n_1618),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_SL g1795 ( 
.A(n_1614),
.B(n_1624),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1668),
.B(n_1535),
.Y(n_1796)
);

INVx5_ASAP7_75t_L g1797 ( 
.A(n_1625),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1592),
.B(n_1533),
.Y(n_1798)
);

INVx2_ASAP7_75t_SL g1799 ( 
.A(n_1614),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1717),
.B(n_1604),
.Y(n_1800)
);

BUFx3_ASAP7_75t_L g1801 ( 
.A(n_1666),
.Y(n_1801)
);

NAND3xp33_ASAP7_75t_L g1802 ( 
.A(n_1651),
.B(n_1569),
.C(n_798),
.Y(n_1802)
);

AOI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1724),
.A2(n_1533),
.B1(n_1537),
.B2(n_1569),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1627),
.B(n_1537),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1720),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1659),
.Y(n_1806)
);

AND2x6_ASAP7_75t_L g1807 ( 
.A(n_1658),
.B(n_987),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_L g1808 ( 
.A(n_1662),
.B(n_799),
.Y(n_1808)
);

AOI22xp33_ASAP7_75t_L g1809 ( 
.A1(n_1724),
.A2(n_973),
.B1(n_978),
.B2(n_945),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1596),
.B(n_1664),
.Y(n_1810)
);

INVx2_ASAP7_75t_SL g1811 ( 
.A(n_1626),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_L g1812 ( 
.A(n_1627),
.B(n_804),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1597),
.B(n_1509),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1722),
.Y(n_1814)
);

AOI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1626),
.A2(n_982),
.B1(n_991),
.B2(n_980),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1599),
.B(n_1509),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1676),
.B(n_815),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1714),
.Y(n_1818)
);

BUFx2_ASAP7_75t_L g1819 ( 
.A(n_1709),
.Y(n_1819)
);

INVx4_ASAP7_75t_L g1820 ( 
.A(n_1625),
.Y(n_1820)
);

INVx4_ASAP7_75t_L g1821 ( 
.A(n_1697),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1721),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_SL g1823 ( 
.A1(n_1716),
.A2(n_1521),
.B1(n_894),
.B2(n_896),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1646),
.B(n_1547),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_SL g1825 ( 
.A(n_1697),
.B(n_827),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1600),
.B(n_1509),
.Y(n_1826)
);

CKINVDCx20_ASAP7_75t_R g1827 ( 
.A(n_1716),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1725),
.Y(n_1828)
);

AND2x2_ASAP7_75t_SL g1829 ( 
.A(n_1704),
.B(n_1404),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_L g1830 ( 
.A(n_1677),
.B(n_822),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1726),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1646),
.Y(n_1832)
);

INVx3_ASAP7_75t_L g1833 ( 
.A(n_1697),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1598),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1603),
.B(n_1509),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1598),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_SL g1837 ( 
.A(n_1678),
.B(n_918),
.Y(n_1837)
);

CKINVDCx20_ASAP7_75t_R g1838 ( 
.A(n_1681),
.Y(n_1838)
);

OR2x6_ASAP7_75t_L g1839 ( 
.A(n_1682),
.B(n_1313),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1649),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1649),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1613),
.Y(n_1842)
);

INVx2_ASAP7_75t_SL g1843 ( 
.A(n_1589),
.Y(n_1843)
);

INVx2_ASAP7_75t_SL g1844 ( 
.A(n_1590),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_1679),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1679),
.B(n_1547),
.Y(n_1846)
);

BUFx6f_ASAP7_75t_L g1847 ( 
.A(n_1652),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1613),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1638),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1638),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1698),
.B(n_1578),
.Y(n_1851)
);

INVx3_ASAP7_75t_L g1852 ( 
.A(n_1698),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1606),
.B(n_1578),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_SL g1854 ( 
.A(n_1708),
.B(n_839),
.Y(n_1854)
);

AND3x2_ASAP7_75t_L g1855 ( 
.A(n_1690),
.B(n_1187),
.C(n_936),
.Y(n_1855)
);

INVx2_ASAP7_75t_SL g1856 ( 
.A(n_1692),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1665),
.Y(n_1857)
);

BUFx3_ASAP7_75t_L g1858 ( 
.A(n_1693),
.Y(n_1858)
);

INVx5_ASAP7_75t_L g1859 ( 
.A(n_1652),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1628),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1708),
.B(n_1575),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1608),
.B(n_999),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1665),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1628),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_L g1865 ( 
.A(n_1694),
.B(n_947),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1695),
.B(n_950),
.Y(n_1866)
);

OAI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1711),
.A2(n_1031),
.B1(n_1079),
.B2(n_1000),
.Y(n_1867)
);

INVx3_ASAP7_75t_L g1868 ( 
.A(n_1713),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1636),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1636),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1609),
.B(n_1082),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1699),
.B(n_1012),
.Y(n_1872)
);

AOI22xp33_ASAP7_75t_L g1873 ( 
.A1(n_1658),
.A2(n_1160),
.B1(n_1196),
.B2(n_1148),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1700),
.B(n_1064),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_L g1875 ( 
.A(n_1701),
.B(n_1097),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1615),
.B(n_1214),
.Y(n_1876)
);

BUFx6f_ASAP7_75t_L g1877 ( 
.A(n_1652),
.Y(n_1877)
);

INVx4_ASAP7_75t_L g1878 ( 
.A(n_1713),
.Y(n_1878)
);

BUFx3_ASAP7_75t_L g1879 ( 
.A(n_1702),
.Y(n_1879)
);

AOI22xp33_ASAP7_75t_L g1880 ( 
.A1(n_1680),
.A2(n_1257),
.B1(n_1265),
.B2(n_1225),
.Y(n_1880)
);

BUFx2_ASAP7_75t_L g1881 ( 
.A(n_1709),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1704),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1703),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1706),
.Y(n_1884)
);

INVxp67_ASAP7_75t_SL g1885 ( 
.A(n_1635),
.Y(n_1885)
);

AND3x2_ASAP7_75t_L g1886 ( 
.A(n_1607),
.B(n_924),
.C(n_906),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1610),
.Y(n_1887)
);

BUFx2_ASAP7_75t_L g1888 ( 
.A(n_1611),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1727),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1735),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1748),
.B(n_1612),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1842),
.B(n_1616),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1742),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1848),
.B(n_1737),
.Y(n_1894)
);

NOR2xp33_ASAP7_75t_SL g1895 ( 
.A(n_1779),
.B(n_1751),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1737),
.B(n_1617),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_SL g1897 ( 
.A(n_1748),
.B(n_1622),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1756),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_SL g1899 ( 
.A(n_1740),
.B(n_1629),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1737),
.B(n_1620),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1757),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1743),
.Y(n_1902)
);

INVxp33_ASAP7_75t_L g1903 ( 
.A(n_1759),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_L g1904 ( 
.A(n_1741),
.B(n_1621),
.Y(n_1904)
);

INVx1_ASAP7_75t_SL g1905 ( 
.A(n_1762),
.Y(n_1905)
);

NOR2xp33_ASAP7_75t_L g1906 ( 
.A(n_1800),
.B(n_1623),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1763),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1744),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1775),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1770),
.B(n_1630),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1849),
.B(n_1711),
.Y(n_1911)
);

NAND2xp33_ASAP7_75t_L g1912 ( 
.A(n_1738),
.B(n_1680),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1747),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1850),
.B(n_1635),
.Y(n_1914)
);

AOI22xp5_ASAP7_75t_L g1915 ( 
.A1(n_1738),
.A2(n_1640),
.B1(n_1643),
.B2(n_1639),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1857),
.B(n_1645),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1738),
.A2(n_1657),
.B1(n_1653),
.B2(n_1680),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1863),
.B(n_1270),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1765),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_SL g1920 ( 
.A(n_1796),
.B(n_842),
.Y(n_1920)
);

NAND2x1_ASAP7_75t_L g1921 ( 
.A(n_1820),
.B(n_1581),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_SL g1922 ( 
.A(n_1811),
.B(n_857),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1776),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1782),
.Y(n_1924)
);

AOI22xp33_ASAP7_75t_L g1925 ( 
.A1(n_1869),
.A2(n_1289),
.B1(n_1296),
.B2(n_1273),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_SL g1926 ( 
.A(n_1773),
.B(n_1799),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1812),
.B(n_1582),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1870),
.B(n_1302),
.Y(n_1928)
);

AOI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1790),
.A2(n_1526),
.B(n_1504),
.Y(n_1929)
);

INVxp67_ASAP7_75t_L g1930 ( 
.A(n_1817),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1767),
.B(n_1320),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1780),
.Y(n_1932)
);

NAND2xp33_ASAP7_75t_SL g1933 ( 
.A(n_1733),
.B(n_1819),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1749),
.B(n_934),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1781),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1783),
.B(n_792),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1784),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1734),
.B(n_1312),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1787),
.B(n_864),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_L g1940 ( 
.A(n_1795),
.B(n_894),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1791),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1805),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1814),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1788),
.B(n_868),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1793),
.B(n_1806),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1803),
.B(n_873),
.Y(n_1946)
);

INVx2_ASAP7_75t_SL g1947 ( 
.A(n_1804),
.Y(n_1947)
);

AOI22xp33_ASAP7_75t_L g1948 ( 
.A1(n_1732),
.A2(n_1035),
.B1(n_987),
.B2(n_837),
.Y(n_1948)
);

NAND2xp33_ASAP7_75t_L g1949 ( 
.A(n_1732),
.B(n_1035),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1810),
.B(n_885),
.Y(n_1950)
);

OR2x2_ASAP7_75t_L g1951 ( 
.A(n_1758),
.B(n_1207),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1808),
.B(n_897),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_L g1953 ( 
.A(n_1754),
.B(n_1764),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1824),
.B(n_899),
.Y(n_1954)
);

NOR2xp33_ASAP7_75t_L g1955 ( 
.A(n_1730),
.B(n_895),
.Y(n_1955)
);

NOR2xp33_ASAP7_75t_L g1956 ( 
.A(n_1802),
.B(n_895),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1846),
.B(n_911),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1851),
.B(n_912),
.Y(n_1958)
);

AOI22xp5_ASAP7_75t_L g1959 ( 
.A1(n_1732),
.A2(n_940),
.B1(n_949),
.B2(n_942),
.Y(n_1959)
);

INVx4_ASAP7_75t_L g1960 ( 
.A(n_1736),
.Y(n_1960)
);

BUFx6f_ASAP7_75t_L g1961 ( 
.A(n_1736),
.Y(n_1961)
);

OR2x6_ASAP7_75t_L g1962 ( 
.A(n_1792),
.B(n_924),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1752),
.B(n_959),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1888),
.Y(n_1964)
);

INVxp67_ASAP7_75t_L g1965 ( 
.A(n_1830),
.Y(n_1965)
);

INVx4_ASAP7_75t_L g1966 ( 
.A(n_1772),
.Y(n_1966)
);

BUFx6f_ASAP7_75t_L g1967 ( 
.A(n_1772),
.Y(n_1967)
);

INVx2_ASAP7_75t_SL g1968 ( 
.A(n_1801),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1777),
.B(n_960),
.Y(n_1969)
);

INVx2_ASAP7_75t_SL g1970 ( 
.A(n_1778),
.Y(n_1970)
);

NOR2xp67_ASAP7_75t_L g1971 ( 
.A(n_1766),
.B(n_1437),
.Y(n_1971)
);

AOI22xp33_ASAP7_75t_L g1972 ( 
.A1(n_1809),
.A2(n_1035),
.B1(n_987),
.B2(n_951),
.Y(n_1972)
);

BUFx6f_ASAP7_75t_L g1973 ( 
.A(n_1847),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1888),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1828),
.Y(n_1975)
);

NOR2xp67_ASAP7_75t_L g1976 ( 
.A(n_1786),
.B(n_1438),
.Y(n_1976)
);

AND2x4_ASAP7_75t_L g1977 ( 
.A(n_1778),
.B(n_1440),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1861),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1818),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1822),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1831),
.Y(n_1981)
);

INVxp67_ASAP7_75t_L g1982 ( 
.A(n_1865),
.Y(n_1982)
);

NAND2x1p5_ASAP7_75t_L g1983 ( 
.A(n_1755),
.B(n_1471),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1834),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1832),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1882),
.B(n_896),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_SL g1987 ( 
.A(n_1750),
.B(n_984),
.Y(n_1987)
);

BUFx3_ASAP7_75t_L g1988 ( 
.A(n_1838),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_SL g1989 ( 
.A(n_1750),
.B(n_993),
.Y(n_1989)
);

INVx4_ASAP7_75t_L g1990 ( 
.A(n_1847),
.Y(n_1990)
);

NOR2xp33_ASAP7_75t_L g1991 ( 
.A(n_1840),
.B(n_1841),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_SL g1992 ( 
.A(n_1755),
.B(n_1003),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1883),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_1794),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1866),
.B(n_1018),
.Y(n_1995)
);

NAND3xp33_ASAP7_75t_L g1996 ( 
.A(n_1872),
.B(n_801),
.C(n_787),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1874),
.B(n_792),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1875),
.B(n_1022),
.Y(n_1998)
);

AND2x4_ASAP7_75t_L g1999 ( 
.A(n_1858),
.B(n_1443),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1769),
.B(n_1026),
.Y(n_2000)
);

INVx2_ASAP7_75t_SL g2001 ( 
.A(n_1839),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1836),
.Y(n_2002)
);

OR2x6_ASAP7_75t_L g2003 ( 
.A(n_1819),
.B(n_938),
.Y(n_2003)
);

AOI22xp33_ASAP7_75t_L g2004 ( 
.A1(n_1739),
.A2(n_987),
.B1(n_951),
.B2(n_986),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_SL g2005 ( 
.A(n_1774),
.B(n_985),
.Y(n_2005)
);

INVx3_ASAP7_75t_L g2006 ( 
.A(n_1877),
.Y(n_2006)
);

NOR2xp33_ASAP7_75t_L g2007 ( 
.A(n_1881),
.B(n_985),
.Y(n_2007)
);

INVx2_ASAP7_75t_SL g2008 ( 
.A(n_1839),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1860),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1864),
.Y(n_2010)
);

BUFx2_ASAP7_75t_L g2011 ( 
.A(n_1739),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1884),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1771),
.B(n_1033),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1739),
.B(n_1043),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1887),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1852),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_1827),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1853),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1868),
.Y(n_2019)
);

NOR2xp33_ASAP7_75t_L g2020 ( 
.A(n_1881),
.B(n_986),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1885),
.B(n_1049),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1768),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1833),
.Y(n_2023)
);

BUFx6f_ASAP7_75t_L g2024 ( 
.A(n_1877),
.Y(n_2024)
);

NOR2xp33_ASAP7_75t_L g2025 ( 
.A(n_1728),
.B(n_1004),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1843),
.Y(n_2026)
);

AND2x6_ASAP7_75t_L g2027 ( 
.A(n_1798),
.B(n_938),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1844),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1753),
.B(n_1055),
.Y(n_2029)
);

AOI22xp5_ASAP7_75t_L g2030 ( 
.A1(n_1761),
.A2(n_1057),
.B1(n_1062),
.B2(n_1056),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1879),
.Y(n_2031)
);

INVx2_ASAP7_75t_SL g2032 ( 
.A(n_1886),
.Y(n_2032)
);

AND2x6_ASAP7_75t_L g2033 ( 
.A(n_1813),
.B(n_1008),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1856),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1815),
.B(n_1074),
.Y(n_2035)
);

AOI21xp5_ASAP7_75t_L g2036 ( 
.A1(n_1816),
.A2(n_1115),
.B(n_1110),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_SL g2037 ( 
.A(n_1755),
.B(n_1121),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_SL g2038 ( 
.A(n_1797),
.B(n_1123),
.Y(n_2038)
);

NOR2xp33_ASAP7_75t_SL g2039 ( 
.A(n_1837),
.B(n_1004),
.Y(n_2039)
);

A2O1A1Ixp33_ASAP7_75t_L g2040 ( 
.A1(n_1862),
.A2(n_1259),
.B(n_1311),
.C(n_1229),
.Y(n_2040)
);

OR2x2_ASAP7_75t_L g2041 ( 
.A(n_1760),
.B(n_1444),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1820),
.Y(n_2042)
);

AND2x4_ASAP7_75t_L g2043 ( 
.A(n_1845),
.B(n_1446),
.Y(n_2043)
);

NOR2xp33_ASAP7_75t_R g2044 ( 
.A(n_1829),
.B(n_1139),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1871),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1876),
.Y(n_2046)
);

INVx3_ASAP7_75t_L g2047 ( 
.A(n_1731),
.Y(n_2047)
);

INVxp67_ASAP7_75t_L g2048 ( 
.A(n_1746),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1729),
.B(n_900),
.Y(n_2049)
);

BUFx6f_ASAP7_75t_L g2050 ( 
.A(n_1797),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_SL g2051 ( 
.A(n_1797),
.B(n_1141),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1878),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1873),
.B(n_1149),
.Y(n_2053)
);

NOR2xp33_ASAP7_75t_L g2054 ( 
.A(n_1825),
.B(n_1014),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_L g2055 ( 
.A(n_1854),
.B(n_1014),
.Y(n_2055)
);

AOI22xp33_ASAP7_75t_L g2056 ( 
.A1(n_1880),
.A2(n_1068),
.B1(n_1093),
.B2(n_1053),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1785),
.B(n_1156),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1826),
.Y(n_2058)
);

BUFx6f_ASAP7_75t_L g2059 ( 
.A(n_1859),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_SL g2060 ( 
.A(n_1859),
.B(n_1165),
.Y(n_2060)
);

BUFx6f_ASAP7_75t_L g2061 ( 
.A(n_1859),
.Y(n_2061)
);

AOI21xp5_ASAP7_75t_L g2062 ( 
.A1(n_1835),
.A2(n_1173),
.B(n_1169),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1930),
.B(n_1785),
.Y(n_2063)
);

NOR2x2_ASAP7_75t_L g2064 ( 
.A(n_2003),
.B(n_1823),
.Y(n_2064)
);

NAND2x1p5_ASAP7_75t_L g2065 ( 
.A(n_2047),
.B(n_1960),
.Y(n_2065)
);

AOI22xp33_ASAP7_75t_L g2066 ( 
.A1(n_1953),
.A2(n_1867),
.B1(n_1785),
.B2(n_1807),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_SL g2067 ( 
.A(n_1965),
.B(n_1895),
.Y(n_2067)
);

AOI22xp33_ASAP7_75t_L g2068 ( 
.A1(n_1956),
.A2(n_1807),
.B1(n_1789),
.B2(n_1745),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_1997),
.B(n_1855),
.Y(n_2069)
);

BUFx3_ASAP7_75t_L g2070 ( 
.A(n_1988),
.Y(n_2070)
);

NOR2x1p5_ASAP7_75t_L g2071 ( 
.A(n_2041),
.B(n_1821),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1889),
.Y(n_2072)
);

HB1xp67_ASAP7_75t_L g2073 ( 
.A(n_1964),
.Y(n_2073)
);

INVxp67_ASAP7_75t_SL g2074 ( 
.A(n_1974),
.Y(n_2074)
);

A2O1A1Ixp33_ASAP7_75t_L g2075 ( 
.A1(n_1934),
.A2(n_1010),
.B(n_1015),
.C(n_1007),
.Y(n_2075)
);

AOI21xp5_ASAP7_75t_L g2076 ( 
.A1(n_1912),
.A2(n_1807),
.B(n_1197),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_1947),
.Y(n_2077)
);

NAND3xp33_ASAP7_75t_L g2078 ( 
.A(n_1938),
.B(n_805),
.C(n_803),
.Y(n_2078)
);

OR2x2_ASAP7_75t_L g2079 ( 
.A(n_1905),
.B(n_1448),
.Y(n_2079)
);

BUFx3_ASAP7_75t_L g2080 ( 
.A(n_1961),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1980),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1890),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1893),
.Y(n_2083)
);

BUFx2_ASAP7_75t_L g2084 ( 
.A(n_2003),
.Y(n_2084)
);

BUFx2_ASAP7_75t_L g2085 ( 
.A(n_1961),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1902),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1908),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1982),
.B(n_1194),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1927),
.B(n_1198),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_2045),
.B(n_1204),
.Y(n_2090)
);

BUFx4f_ASAP7_75t_L g2091 ( 
.A(n_1967),
.Y(n_2091)
);

A2O1A1Ixp33_ASAP7_75t_L g2092 ( 
.A1(n_2055),
.A2(n_1017),
.B(n_1030),
.C(n_1029),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2046),
.B(n_2018),
.Y(n_2093)
);

AOI22xp33_ASAP7_75t_SL g2094 ( 
.A1(n_2039),
.A2(n_1068),
.B1(n_1158),
.B2(n_1053),
.Y(n_2094)
);

NOR2xp33_ASAP7_75t_L g2095 ( 
.A(n_1940),
.B(n_1955),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_1952),
.B(n_1906),
.Y(n_2096)
);

NAND2xp33_ASAP7_75t_SL g2097 ( 
.A(n_2044),
.B(n_1093),
.Y(n_2097)
);

INVx4_ASAP7_75t_L g2098 ( 
.A(n_2050),
.Y(n_2098)
);

INVx2_ASAP7_75t_SL g2099 ( 
.A(n_2043),
.Y(n_2099)
);

BUFx4f_ASAP7_75t_L g2100 ( 
.A(n_2050),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_1968),
.B(n_1220),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1913),
.B(n_1228),
.Y(n_2102)
);

NOR2xp33_ASAP7_75t_R g2103 ( 
.A(n_1933),
.B(n_1107),
.Y(n_2103)
);

INVx2_ASAP7_75t_SL g2104 ( 
.A(n_2043),
.Y(n_2104)
);

AND2x4_ASAP7_75t_L g2105 ( 
.A(n_1970),
.B(n_1451),
.Y(n_2105)
);

NOR2xp33_ASAP7_75t_L g2106 ( 
.A(n_2007),
.B(n_1107),
.Y(n_2106)
);

NOR2xp33_ASAP7_75t_R g2107 ( 
.A(n_1994),
.B(n_1155),
.Y(n_2107)
);

INVx2_ASAP7_75t_SL g2108 ( 
.A(n_1977),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1919),
.B(n_1230),
.Y(n_2109)
);

OR2x2_ASAP7_75t_L g2110 ( 
.A(n_1951),
.B(n_1454),
.Y(n_2110)
);

NOR2xp33_ASAP7_75t_L g2111 ( 
.A(n_2020),
.B(n_1155),
.Y(n_2111)
);

INVx3_ASAP7_75t_L g2112 ( 
.A(n_2050),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1945),
.B(n_1261),
.Y(n_2113)
);

NOR2x1p5_ASAP7_75t_L g2114 ( 
.A(n_2017),
.B(n_809),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_SL g2115 ( 
.A(n_1978),
.B(n_1995),
.Y(n_2115)
);

INVx4_ASAP7_75t_L g2116 ( 
.A(n_2059),
.Y(n_2116)
);

AOI22xp33_ASAP7_75t_L g2117 ( 
.A1(n_2054),
.A2(n_1182),
.B1(n_1192),
.B2(n_1158),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1932),
.Y(n_2118)
);

INVx3_ASAP7_75t_L g2119 ( 
.A(n_2059),
.Y(n_2119)
);

HB1xp67_ASAP7_75t_L g2120 ( 
.A(n_1967),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1935),
.B(n_1268),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1898),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1892),
.B(n_1998),
.Y(n_2123)
);

AOI22xp5_ASAP7_75t_L g2124 ( 
.A1(n_1926),
.A2(n_1315),
.B1(n_1278),
.B2(n_1282),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1979),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1950),
.B(n_1271),
.Y(n_2126)
);

INVx3_ASAP7_75t_SL g2127 ( 
.A(n_1962),
.Y(n_2127)
);

O2A1O1Ixp33_ASAP7_75t_SL g2128 ( 
.A1(n_1894),
.A2(n_1042),
.B(n_1059),
.C(n_1058),
.Y(n_2128)
);

BUFx3_ASAP7_75t_L g2129 ( 
.A(n_1973),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_1904),
.B(n_1286),
.Y(n_2130)
);

CKINVDCx5p33_ASAP7_75t_R g2131 ( 
.A(n_1973),
.Y(n_2131)
);

NOR2xp33_ASAP7_75t_R g2132 ( 
.A(n_2011),
.B(n_2006),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1981),
.Y(n_2133)
);

NAND2x1_ASAP7_75t_L g2134 ( 
.A(n_2059),
.B(n_1457),
.Y(n_2134)
);

BUFx3_ASAP7_75t_L g2135 ( 
.A(n_2024),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1985),
.Y(n_2136)
);

NAND2xp33_ASAP7_75t_R g2137 ( 
.A(n_1986),
.B(n_1297),
.Y(n_2137)
);

BUFx3_ASAP7_75t_L g2138 ( 
.A(n_2024),
.Y(n_2138)
);

CKINVDCx20_ASAP7_75t_R g2139 ( 
.A(n_1987),
.Y(n_2139)
);

AOI22xp5_ASAP7_75t_L g2140 ( 
.A1(n_1920),
.A2(n_1304),
.B1(n_1309),
.B2(n_1299),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1918),
.B(n_811),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_SL g2142 ( 
.A(n_2034),
.B(n_1182),
.Y(n_2142)
);

AND2x4_ASAP7_75t_L g2143 ( 
.A(n_1977),
.B(n_1459),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1901),
.Y(n_2144)
);

BUFx6f_ASAP7_75t_L g2145 ( 
.A(n_2061),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1907),
.Y(n_2146)
);

AOI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_1991),
.A2(n_1242),
.B1(n_1252),
.B2(n_1192),
.Y(n_2147)
);

NOR3xp33_ASAP7_75t_SL g2148 ( 
.A(n_2025),
.B(n_817),
.C(n_813),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1993),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_1909),
.Y(n_2150)
);

INVxp67_ASAP7_75t_L g2151 ( 
.A(n_1936),
.Y(n_2151)
);

AND2x4_ASAP7_75t_L g2152 ( 
.A(n_2031),
.B(n_1461),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_1923),
.Y(n_2153)
);

INVx2_ASAP7_75t_SL g2154 ( 
.A(n_1999),
.Y(n_2154)
);

AND2x4_ASAP7_75t_L g2155 ( 
.A(n_2016),
.B(n_1462),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1911),
.B(n_818),
.Y(n_2156)
);

NAND2x1p5_ASAP7_75t_L g2157 ( 
.A(n_1966),
.B(n_1990),
.Y(n_2157)
);

INVx2_ASAP7_75t_SL g2158 ( 
.A(n_1999),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_1924),
.Y(n_2159)
);

AND2x4_ASAP7_75t_L g2160 ( 
.A(n_2019),
.B(n_1063),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_SL g2161 ( 
.A(n_1954),
.B(n_1242),
.Y(n_2161)
);

NOR2xp33_ASAP7_75t_L g2162 ( 
.A(n_2048),
.B(n_1252),
.Y(n_2162)
);

AND2x4_ASAP7_75t_L g2163 ( 
.A(n_2012),
.B(n_1070),
.Y(n_2163)
);

OR2x2_ASAP7_75t_L g2164 ( 
.A(n_2056),
.B(n_820),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1937),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1941),
.Y(n_2166)
);

BUFx3_ASAP7_75t_L g2167 ( 
.A(n_2001),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2015),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_1942),
.Y(n_2169)
);

AND2x4_ASAP7_75t_L g2170 ( 
.A(n_1899),
.B(n_1072),
.Y(n_2170)
);

NOR2xp33_ASAP7_75t_L g2171 ( 
.A(n_2049),
.B(n_1275),
.Y(n_2171)
);

AOI21xp5_ASAP7_75t_L g2172 ( 
.A1(n_2029),
.A2(n_1471),
.B(n_1089),
.Y(n_2172)
);

OAI22xp5_ASAP7_75t_L g2173 ( 
.A1(n_1946),
.A2(n_1928),
.B1(n_1917),
.B2(n_1914),
.Y(n_2173)
);

AOI21x1_ASAP7_75t_L g2174 ( 
.A1(n_1896),
.A2(n_1091),
.B(n_1087),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1943),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_2004),
.B(n_2040),
.Y(n_2176)
);

INVxp67_ASAP7_75t_L g2177 ( 
.A(n_2008),
.Y(n_2177)
);

AOI22xp5_ASAP7_75t_L g2178 ( 
.A1(n_1976),
.A2(n_1317),
.B1(n_1275),
.B2(n_829),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_SL g2179 ( 
.A(n_2061),
.B(n_1317),
.Y(n_2179)
);

INVx5_ASAP7_75t_L g2180 ( 
.A(n_2061),
.Y(n_2180)
);

INVx2_ASAP7_75t_SL g2181 ( 
.A(n_1962),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_1975),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1916),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_1984),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_1971),
.B(n_900),
.Y(n_2185)
);

OR2x2_ASAP7_75t_L g2186 ( 
.A(n_1939),
.B(n_825),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_2002),
.Y(n_2187)
);

BUFx2_ASAP7_75t_L g2188 ( 
.A(n_2032),
.Y(n_2188)
);

OR2x2_ASAP7_75t_L g2189 ( 
.A(n_1944),
.B(n_832),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_1957),
.B(n_841),
.Y(n_2190)
);

BUFx3_ASAP7_75t_L g2191 ( 
.A(n_2026),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1958),
.B(n_845),
.Y(n_2192)
);

AND2x4_ASAP7_75t_L g2193 ( 
.A(n_2028),
.B(n_1092),
.Y(n_2193)
);

NOR2xp33_ASAP7_75t_R g2194 ( 
.A(n_2005),
.B(n_848),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2009),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_1931),
.B(n_849),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_2010),
.Y(n_2197)
);

BUFx3_ASAP7_75t_L g2198 ( 
.A(n_2022),
.Y(n_2198)
);

BUFx3_ASAP7_75t_L g2199 ( 
.A(n_2023),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_SL g2200 ( 
.A(n_1996),
.B(n_1471),
.Y(n_2200)
);

AND2x4_ASAP7_75t_L g2201 ( 
.A(n_1891),
.B(n_1094),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_2000),
.B(n_2013),
.Y(n_2202)
);

AND2x6_ASAP7_75t_SL g2203 ( 
.A(n_1969),
.B(n_1102),
.Y(n_2203)
);

AOI22xp5_ASAP7_75t_L g2204 ( 
.A1(n_1963),
.A2(n_852),
.B1(n_854),
.B2(n_850),
.Y(n_2204)
);

BUFx2_ASAP7_75t_L g2205 ( 
.A(n_2033),
.Y(n_2205)
);

NAND2xp33_ASAP7_75t_L g2206 ( 
.A(n_2027),
.B(n_1298),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1910),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_2042),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1900),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2058),
.Y(n_2210)
);

NOR2xp33_ASAP7_75t_L g2211 ( 
.A(n_1897),
.B(n_860),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1921),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2052),
.Y(n_2213)
);

BUFx2_ASAP7_75t_L g2214 ( 
.A(n_2033),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1915),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_2027),
.B(n_865),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_SL g2217 ( 
.A(n_2021),
.B(n_866),
.Y(n_2217)
);

INVx2_ASAP7_75t_SL g2218 ( 
.A(n_1989),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2027),
.B(n_872),
.Y(n_2219)
);

NOR2xp33_ASAP7_75t_R g2220 ( 
.A(n_2131),
.B(n_2097),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2072),
.Y(n_2221)
);

AND3x2_ASAP7_75t_SL g2222 ( 
.A(n_2081),
.B(n_1118),
.C(n_1008),
.Y(n_2222)
);

AND2x4_ASAP7_75t_L g2223 ( 
.A(n_2099),
.B(n_1922),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2096),
.B(n_2093),
.Y(n_2224)
);

AND2x4_ASAP7_75t_L g2225 ( 
.A(n_2104),
.B(n_2014),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2095),
.B(n_1925),
.Y(n_2226)
);

AND2x4_ASAP7_75t_L g2227 ( 
.A(n_2154),
.B(n_1992),
.Y(n_2227)
);

NOR2xp33_ASAP7_75t_L g2228 ( 
.A(n_2106),
.B(n_2030),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2082),
.Y(n_2229)
);

BUFx3_ASAP7_75t_L g2230 ( 
.A(n_2091),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2207),
.B(n_2035),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_2083),
.Y(n_2232)
);

INVx2_ASAP7_75t_SL g2233 ( 
.A(n_2080),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_2086),
.Y(n_2234)
);

HB1xp67_ASAP7_75t_L g2235 ( 
.A(n_2073),
.Y(n_2235)
);

BUFx3_ASAP7_75t_L g2236 ( 
.A(n_2129),
.Y(n_2236)
);

AOI22xp33_ASAP7_75t_L g2237 ( 
.A1(n_2111),
.A2(n_1972),
.B1(n_2053),
.B2(n_2033),
.Y(n_2237)
);

INVxp67_ASAP7_75t_SL g2238 ( 
.A(n_2074),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2087),
.Y(n_2239)
);

BUFx6f_ASAP7_75t_L g2240 ( 
.A(n_2100),
.Y(n_2240)
);

INVx3_ASAP7_75t_L g2241 ( 
.A(n_2180),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_2118),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2125),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_2171),
.B(n_1903),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_2133),
.Y(n_2245)
);

AND2x4_ASAP7_75t_L g2246 ( 
.A(n_2158),
.B(n_2037),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_2149),
.Y(n_2247)
);

A2O1A1Ixp33_ASAP7_75t_SL g2248 ( 
.A1(n_2211),
.A2(n_1948),
.B(n_1949),
.C(n_1959),
.Y(n_2248)
);

INVx4_ASAP7_75t_L g2249 ( 
.A(n_2180),
.Y(n_2249)
);

A2O1A1Ixp33_ASAP7_75t_L g2250 ( 
.A1(n_2176),
.A2(n_2062),
.B(n_2036),
.C(n_2057),
.Y(n_2250)
);

BUFx8_ASAP7_75t_SL g2251 ( 
.A(n_2070),
.Y(n_2251)
);

OR2x6_ASAP7_75t_L g2252 ( 
.A(n_2157),
.B(n_1983),
.Y(n_2252)
);

AND3x2_ASAP7_75t_SL g2253 ( 
.A(n_2213),
.B(n_1125),
.C(n_1118),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2136),
.Y(n_2254)
);

BUFx2_ASAP7_75t_L g2255 ( 
.A(n_2135),
.Y(n_2255)
);

OR2x2_ASAP7_75t_L g2256 ( 
.A(n_2110),
.B(n_2038),
.Y(n_2256)
);

AND3x1_ASAP7_75t_SL g2257 ( 
.A(n_2114),
.B(n_1322),
.C(n_1319),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2168),
.Y(n_2258)
);

CKINVDCx16_ASAP7_75t_R g2259 ( 
.A(n_2107),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_SL g2260 ( 
.A(n_2094),
.B(n_2051),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2122),
.Y(n_2261)
);

INVxp67_ASAP7_75t_SL g2262 ( 
.A(n_2077),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2123),
.B(n_2060),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_2162),
.B(n_900),
.Y(n_2264)
);

BUFx3_ASAP7_75t_L g2265 ( 
.A(n_2138),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2210),
.Y(n_2266)
);

AOI22xp5_ASAP7_75t_L g2267 ( 
.A1(n_2137),
.A2(n_2161),
.B1(n_2139),
.B2(n_2067),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2183),
.B(n_2089),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_2144),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2175),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2146),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2150),
.Y(n_2272)
);

OAI21xp5_ASAP7_75t_L g2273 ( 
.A1(n_2202),
.A2(n_1929),
.B(n_1109),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2156),
.B(n_1103),
.Y(n_2274)
);

AOI22xp5_ASAP7_75t_L g2275 ( 
.A1(n_2069),
.A2(n_876),
.B1(n_877),
.B2(n_875),
.Y(n_2275)
);

OR2x6_ASAP7_75t_L g2276 ( 
.A(n_2065),
.B(n_1125),
.Y(n_2276)
);

INVx4_ASAP7_75t_L g2277 ( 
.A(n_2180),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2130),
.B(n_2141),
.Y(n_2278)
);

INVx2_ASAP7_75t_SL g2279 ( 
.A(n_2100),
.Y(n_2279)
);

NOR2x2_ASAP7_75t_L g2280 ( 
.A(n_2153),
.B(n_1135),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2159),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2165),
.Y(n_2282)
);

AO22x1_ASAP7_75t_L g2283 ( 
.A1(n_2127),
.A2(n_882),
.B1(n_884),
.B2(n_878),
.Y(n_2283)
);

BUFx2_ASAP7_75t_L g2284 ( 
.A(n_2085),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2166),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2169),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2182),
.Y(n_2287)
);

BUFx2_ASAP7_75t_L g2288 ( 
.A(n_2084),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2143),
.B(n_927),
.Y(n_2289)
);

AND2x4_ASAP7_75t_SL g2290 ( 
.A(n_2098),
.B(n_927),
.Y(n_2290)
);

INVx3_ASAP7_75t_L g2291 ( 
.A(n_2098),
.Y(n_2291)
);

AND3x1_ASAP7_75t_SL g2292 ( 
.A(n_2071),
.B(n_1307),
.C(n_1306),
.Y(n_2292)
);

NOR2xp33_ASAP7_75t_L g2293 ( 
.A(n_2088),
.B(n_886),
.Y(n_2293)
);

CKINVDCx5p33_ASAP7_75t_R g2294 ( 
.A(n_2103),
.Y(n_2294)
);

AND2x4_ASAP7_75t_L g2295 ( 
.A(n_2108),
.B(n_1112),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2209),
.B(n_1113),
.Y(n_2296)
);

BUFx2_ASAP7_75t_L g2297 ( 
.A(n_2120),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2195),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2184),
.Y(n_2299)
);

HB1xp67_ASAP7_75t_L g2300 ( 
.A(n_2188),
.Y(n_2300)
);

NOR2xp33_ASAP7_75t_L g2301 ( 
.A(n_2147),
.B(n_888),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_SL g2302 ( 
.A(n_2194),
.B(n_927),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2090),
.B(n_1120),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2113),
.B(n_1126),
.Y(n_2304)
);

INVxp67_ASAP7_75t_SL g2305 ( 
.A(n_2191),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_2187),
.Y(n_2306)
);

AOI22x1_ASAP7_75t_L g2307 ( 
.A1(n_2172),
.A2(n_1143),
.B1(n_1147),
.B2(n_1135),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_SL g2308 ( 
.A(n_2178),
.B(n_967),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_SL g2309 ( 
.A(n_2151),
.B(n_967),
.Y(n_2309)
);

NOR2xp33_ASAP7_75t_L g2310 ( 
.A(n_2179),
.B(n_891),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2197),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2190),
.B(n_1129),
.Y(n_2312)
);

NOR2xp33_ASAP7_75t_L g2313 ( 
.A(n_2117),
.B(n_893),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_SL g2314 ( 
.A(n_2079),
.B(n_967),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2192),
.B(n_1131),
.Y(n_2315)
);

HB1xp67_ASAP7_75t_L g2316 ( 
.A(n_2143),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2155),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2163),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2163),
.Y(n_2319)
);

INVx4_ASAP7_75t_L g2320 ( 
.A(n_2145),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2155),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2160),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2208),
.Y(n_2323)
);

NAND3xp33_ASAP7_75t_L g2324 ( 
.A(n_2078),
.B(n_905),
.C(n_902),
.Y(n_2324)
);

BUFx6f_ASAP7_75t_L g2325 ( 
.A(n_2145),
.Y(n_2325)
);

NOR2xp33_ASAP7_75t_L g2326 ( 
.A(n_2142),
.B(n_908),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2105),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2160),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_2105),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2196),
.B(n_2115),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2126),
.B(n_1138),
.Y(n_2331)
);

NOR2xp33_ASAP7_75t_L g2332 ( 
.A(n_2186),
.B(n_913),
.Y(n_2332)
);

HB1xp67_ASAP7_75t_L g2333 ( 
.A(n_2145),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2189),
.B(n_1144),
.Y(n_2334)
);

AND2x4_ASAP7_75t_L g2335 ( 
.A(n_2198),
.B(n_2199),
.Y(n_2335)
);

A2O1A1Ixp33_ASAP7_75t_L g2336 ( 
.A1(n_2215),
.A2(n_1152),
.B(n_1168),
.C(n_1150),
.Y(n_2336)
);

INVx3_ASAP7_75t_L g2337 ( 
.A(n_2116),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2170),
.B(n_1175),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2170),
.B(n_1178),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2102),
.B(n_1183),
.Y(n_2340)
);

AND2x4_ASAP7_75t_SL g2341 ( 
.A(n_2116),
.B(n_1044),
.Y(n_2341)
);

BUFx2_ASAP7_75t_SL g2342 ( 
.A(n_2167),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2109),
.B(n_1186),
.Y(n_2343)
);

AND2x2_ASAP7_75t_L g2344 ( 
.A(n_2185),
.B(n_1044),
.Y(n_2344)
);

NOR2xp33_ASAP7_75t_L g2345 ( 
.A(n_2164),
.B(n_914),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2121),
.B(n_1188),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_SL g2347 ( 
.A(n_2132),
.B(n_1044),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2218),
.B(n_1191),
.Y(n_2348)
);

AND3x1_ASAP7_75t_SL g2349 ( 
.A(n_2064),
.B(n_1206),
.C(n_1195),
.Y(n_2349)
);

NOR2xp33_ASAP7_75t_R g2350 ( 
.A(n_2112),
.B(n_547),
.Y(n_2350)
);

NOR2x1p5_ASAP7_75t_L g2351 ( 
.A(n_2134),
.B(n_915),
.Y(n_2351)
);

NOR2xp33_ASAP7_75t_L g2352 ( 
.A(n_2063),
.B(n_2217),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2152),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2152),
.Y(n_2354)
);

HB1xp67_ASAP7_75t_L g2355 ( 
.A(n_2177),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_SL g2356 ( 
.A(n_2148),
.B(n_2181),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2201),
.B(n_1210),
.Y(n_2357)
);

NOR2xp33_ASAP7_75t_L g2358 ( 
.A(n_2204),
.B(n_916),
.Y(n_2358)
);

HB1xp67_ASAP7_75t_L g2359 ( 
.A(n_2112),
.Y(n_2359)
);

BUFx3_ASAP7_75t_L g2360 ( 
.A(n_2119),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_2193),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2193),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2174),
.Y(n_2363)
);

AOI22xp33_ASAP7_75t_L g2364 ( 
.A1(n_2201),
.A2(n_1248),
.B1(n_1255),
.B2(n_1240),
.Y(n_2364)
);

BUFx5_ASAP7_75t_L g2365 ( 
.A(n_2212),
.Y(n_2365)
);

AOI22xp33_ASAP7_75t_L g2366 ( 
.A1(n_2206),
.A2(n_1248),
.B1(n_1255),
.B2(n_1240),
.Y(n_2366)
);

AOI22xp33_ASAP7_75t_L g2367 ( 
.A1(n_2219),
.A2(n_1248),
.B1(n_1255),
.B2(n_1240),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2075),
.B(n_917),
.Y(n_2368)
);

AOI22xp33_ASAP7_75t_L g2369 ( 
.A1(n_2216),
.A2(n_1217),
.B1(n_1218),
.B2(n_1211),
.Y(n_2369)
);

NAND3xp33_ASAP7_75t_SL g2370 ( 
.A(n_2092),
.B(n_922),
.C(n_920),
.Y(n_2370)
);

O2A1O1Ixp5_ASAP7_75t_L g2371 ( 
.A1(n_2173),
.A2(n_1147),
.B(n_1180),
.C(n_1143),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2205),
.B(n_1221),
.Y(n_2372)
);

OAI21x1_ASAP7_75t_L g2373 ( 
.A1(n_2371),
.A2(n_2273),
.B(n_2363),
.Y(n_2373)
);

INVx5_ASAP7_75t_L g2374 ( 
.A(n_2240),
.Y(n_2374)
);

BUFx2_ASAP7_75t_L g2375 ( 
.A(n_2238),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2266),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2232),
.Y(n_2377)
);

CKINVDCx5p33_ASAP7_75t_R g2378 ( 
.A(n_2251),
.Y(n_2378)
);

OR2x2_ASAP7_75t_L g2379 ( 
.A(n_2224),
.B(n_2214),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2234),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2242),
.Y(n_2381)
);

OR2x2_ASAP7_75t_L g2382 ( 
.A(n_2268),
.B(n_2200),
.Y(n_2382)
);

A2O1A1Ixp33_ASAP7_75t_L g2383 ( 
.A1(n_2228),
.A2(n_2066),
.B(n_2140),
.C(n_2076),
.Y(n_2383)
);

AOI21x1_ASAP7_75t_L g2384 ( 
.A1(n_2278),
.A2(n_2263),
.B(n_2296),
.Y(n_2384)
);

AO21x2_ASAP7_75t_L g2385 ( 
.A1(n_2250),
.A2(n_2128),
.B(n_2101),
.Y(n_2385)
);

AO31x2_ASAP7_75t_L g2386 ( 
.A1(n_2352),
.A2(n_1200),
.A3(n_1219),
.B(n_1180),
.Y(n_2386)
);

OAI21x1_ASAP7_75t_L g2387 ( 
.A1(n_2307),
.A2(n_2068),
.B(n_2119),
.Y(n_2387)
);

NOR2xp33_ASAP7_75t_L g2388 ( 
.A(n_2267),
.B(n_2203),
.Y(n_2388)
);

BUFx12f_ASAP7_75t_L g2389 ( 
.A(n_2240),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_SL g2390 ( 
.A(n_2226),
.B(n_2124),
.Y(n_2390)
);

AND2x4_ASAP7_75t_L g2391 ( 
.A(n_2236),
.B(n_1222),
.Y(n_2391)
);

OA22x2_ASAP7_75t_L g2392 ( 
.A1(n_2308),
.A2(n_929),
.B1(n_930),
.B2(n_926),
.Y(n_2392)
);

OAI21x1_ASAP7_75t_L g2393 ( 
.A1(n_2270),
.A2(n_1219),
.B(n_1200),
.Y(n_2393)
);

AOI21xp5_ASAP7_75t_L g2394 ( 
.A1(n_2248),
.A2(n_2231),
.B(n_2330),
.Y(n_2394)
);

A2O1A1Ixp33_ASAP7_75t_L g2395 ( 
.A1(n_2358),
.A2(n_1290),
.B(n_1295),
.C(n_1287),
.Y(n_2395)
);

AO21x1_ASAP7_75t_L g2396 ( 
.A1(n_2293),
.A2(n_1231),
.B(n_1224),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_2245),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2345),
.B(n_933),
.Y(n_2398)
);

AND2x2_ASAP7_75t_L g2399 ( 
.A(n_2344),
.B(n_1234),
.Y(n_2399)
);

OAI22x1_ASAP7_75t_L g2400 ( 
.A1(n_2260),
.A2(n_2301),
.B1(n_2313),
.B2(n_2302),
.Y(n_2400)
);

INVx3_ASAP7_75t_L g2401 ( 
.A(n_2230),
.Y(n_2401)
);

AO21x1_ASAP7_75t_L g2402 ( 
.A1(n_2274),
.A2(n_1246),
.B(n_1238),
.Y(n_2402)
);

OAI21x1_ASAP7_75t_L g2403 ( 
.A1(n_2298),
.A2(n_1290),
.B(n_1287),
.Y(n_2403)
);

AOI22xp5_ASAP7_75t_L g2404 ( 
.A1(n_2244),
.A2(n_941),
.B1(n_952),
.B2(n_937),
.Y(n_2404)
);

AOI22xp33_ASAP7_75t_L g2405 ( 
.A1(n_2370),
.A2(n_1260),
.B1(n_1263),
.B2(n_1253),
.Y(n_2405)
);

OAI21xp5_ASAP7_75t_L g2406 ( 
.A1(n_2332),
.A2(n_2303),
.B(n_2331),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2264),
.B(n_955),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2247),
.Y(n_2408)
);

OAI21x1_ASAP7_75t_L g2409 ( 
.A1(n_2221),
.A2(n_1314),
.B(n_1295),
.Y(n_2409)
);

HB1xp67_ASAP7_75t_L g2410 ( 
.A(n_2235),
.Y(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_2327),
.B(n_2329),
.Y(n_2411)
);

NAND2x1p5_ASAP7_75t_L g2412 ( 
.A(n_2249),
.B(n_1280),
.Y(n_2412)
);

A2O1A1Ixp33_ASAP7_75t_L g2413 ( 
.A1(n_2237),
.A2(n_2324),
.B(n_2304),
.C(n_2315),
.Y(n_2413)
);

OAI21x1_ASAP7_75t_SL g2414 ( 
.A1(n_2229),
.A2(n_1314),
.B(n_1292),
.Y(n_2414)
);

AOI211x1_ASAP7_75t_L g2415 ( 
.A1(n_2356),
.A2(n_957),
.B(n_961),
.C(n_956),
.Y(n_2415)
);

AO31x2_ASAP7_75t_L g2416 ( 
.A1(n_2336),
.A2(n_553),
.A3(n_554),
.B(n_548),
.Y(n_2416)
);

O2A1O1Ixp33_ASAP7_75t_L g2417 ( 
.A1(n_2314),
.A2(n_963),
.B(n_968),
.C(n_962),
.Y(n_2417)
);

NAND2xp33_ASAP7_75t_L g2418 ( 
.A(n_2240),
.B(n_970),
.Y(n_2418)
);

NAND2x1p5_ASAP7_75t_L g2419 ( 
.A(n_2249),
.B(n_556),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2316),
.B(n_971),
.Y(n_2420)
);

AO21x1_ASAP7_75t_L g2421 ( 
.A1(n_2312),
.A2(n_0),
.B(n_2),
.Y(n_2421)
);

OAI21xp5_ASAP7_75t_L g2422 ( 
.A1(n_2340),
.A2(n_2346),
.B(n_2343),
.Y(n_2422)
);

AOI21x1_ASAP7_75t_L g2423 ( 
.A1(n_2334),
.A2(n_563),
.B(n_561),
.Y(n_2423)
);

INVx1_ASAP7_75t_SL g2424 ( 
.A(n_2284),
.Y(n_2424)
);

OAI21x1_ASAP7_75t_L g2425 ( 
.A1(n_2239),
.A2(n_565),
.B(n_564),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2326),
.B(n_972),
.Y(n_2426)
);

OA21x2_ASAP7_75t_L g2427 ( 
.A1(n_2243),
.A2(n_979),
.B(n_977),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2254),
.Y(n_2428)
);

BUFx3_ASAP7_75t_L g2429 ( 
.A(n_2265),
.Y(n_2429)
);

OAI21x1_ASAP7_75t_SL g2430 ( 
.A1(n_2258),
.A2(n_4),
.B(n_5),
.Y(n_2430)
);

NAND2x1p5_ASAP7_75t_L g2431 ( 
.A(n_2277),
.B(n_566),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2310),
.B(n_995),
.Y(n_2432)
);

OAI21x1_ASAP7_75t_L g2433 ( 
.A1(n_2323),
.A2(n_568),
.B(n_567),
.Y(n_2433)
);

OAI21x1_ASAP7_75t_L g2434 ( 
.A1(n_2271),
.A2(n_570),
.B(n_569),
.Y(n_2434)
);

BUFx3_ASAP7_75t_L g2435 ( 
.A(n_2255),
.Y(n_2435)
);

AO22x2_ASAP7_75t_L g2436 ( 
.A1(n_2322),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_2436)
);

NOR2x1_ASAP7_75t_L g2437 ( 
.A(n_2277),
.B(n_996),
.Y(n_2437)
);

AND2x4_ASAP7_75t_L g2438 ( 
.A(n_2335),
.B(n_573),
.Y(n_2438)
);

OAI21x1_ASAP7_75t_L g2439 ( 
.A1(n_2272),
.A2(n_581),
.B(n_580),
.Y(n_2439)
);

NAND3xp33_ASAP7_75t_L g2440 ( 
.A(n_2366),
.B(n_1005),
.C(n_1002),
.Y(n_2440)
);

OAI21x1_ASAP7_75t_L g2441 ( 
.A1(n_2281),
.A2(n_583),
.B(n_582),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2305),
.B(n_2256),
.Y(n_2442)
);

OAI21xp5_ASAP7_75t_L g2443 ( 
.A1(n_2368),
.A2(n_2348),
.B(n_2372),
.Y(n_2443)
);

NOR2xp33_ASAP7_75t_L g2444 ( 
.A(n_2259),
.B(n_2355),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2335),
.B(n_1009),
.Y(n_2445)
);

OAI22xp5_ASAP7_75t_L g2446 ( 
.A1(n_2262),
.A2(n_1019),
.B1(n_1020),
.B2(n_1013),
.Y(n_2446)
);

OAI21x1_ASAP7_75t_L g2447 ( 
.A1(n_2282),
.A2(n_587),
.B(n_585),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2317),
.B(n_1024),
.Y(n_2448)
);

OA22x2_ASAP7_75t_L g2449 ( 
.A1(n_2275),
.A2(n_1028),
.B1(n_1032),
.B2(n_1025),
.Y(n_2449)
);

INVx2_ASAP7_75t_SL g2450 ( 
.A(n_2233),
.Y(n_2450)
);

BUFx2_ASAP7_75t_L g2451 ( 
.A(n_2288),
.Y(n_2451)
);

AOI21xp5_ASAP7_75t_L g2452 ( 
.A1(n_2225),
.A2(n_592),
.B(n_588),
.Y(n_2452)
);

OAI21x1_ASAP7_75t_L g2453 ( 
.A1(n_2286),
.A2(n_594),
.B(n_593),
.Y(n_2453)
);

AOI21xp5_ASAP7_75t_L g2454 ( 
.A1(n_2225),
.A2(n_598),
.B(n_595),
.Y(n_2454)
);

AND2x2_ASAP7_75t_L g2455 ( 
.A(n_2361),
.B(n_1034),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_SL g2456 ( 
.A(n_2328),
.B(n_1300),
.Y(n_2456)
);

OAI21x1_ASAP7_75t_L g2457 ( 
.A1(n_2287),
.A2(n_600),
.B(n_599),
.Y(n_2457)
);

OAI21xp5_ASAP7_75t_L g2458 ( 
.A1(n_2369),
.A2(n_1308),
.B(n_1305),
.Y(n_2458)
);

OAI21xp5_ASAP7_75t_L g2459 ( 
.A1(n_2367),
.A2(n_1316),
.B(n_1310),
.Y(n_2459)
);

OAI21x1_ASAP7_75t_L g2460 ( 
.A1(n_2299),
.A2(n_604),
.B(n_602),
.Y(n_2460)
);

BUFx2_ASAP7_75t_L g2461 ( 
.A(n_2297),
.Y(n_2461)
);

OR2x6_ASAP7_75t_L g2462 ( 
.A(n_2342),
.B(n_606),
.Y(n_2462)
);

OAI22xp5_ASAP7_75t_L g2463 ( 
.A1(n_2354),
.A2(n_1037),
.B1(n_1041),
.B2(n_1036),
.Y(n_2463)
);

OAI21x1_ASAP7_75t_L g2464 ( 
.A1(n_2311),
.A2(n_611),
.B(n_610),
.Y(n_2464)
);

AND2x4_ASAP7_75t_L g2465 ( 
.A(n_2279),
.B(n_613),
.Y(n_2465)
);

AOI21x1_ASAP7_75t_L g2466 ( 
.A1(n_2338),
.A2(n_615),
.B(n_614),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2353),
.B(n_2357),
.Y(n_2467)
);

OAI22xp5_ASAP7_75t_L g2468 ( 
.A1(n_2300),
.A2(n_1048),
.B1(n_1050),
.B2(n_1046),
.Y(n_2468)
);

BUFx4_ASAP7_75t_SL g2469 ( 
.A(n_2360),
.Y(n_2469)
);

AOI21xp5_ASAP7_75t_L g2470 ( 
.A1(n_2321),
.A2(n_619),
.B(n_618),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2261),
.Y(n_2471)
);

BUFx2_ASAP7_75t_L g2472 ( 
.A(n_2333),
.Y(n_2472)
);

OAI21x1_ASAP7_75t_L g2473 ( 
.A1(n_2269),
.A2(n_2306),
.B(n_2285),
.Y(n_2473)
);

BUFx2_ASAP7_75t_L g2474 ( 
.A(n_2359),
.Y(n_2474)
);

AOI21xp5_ASAP7_75t_L g2475 ( 
.A1(n_2223),
.A2(n_623),
.B(n_621),
.Y(n_2475)
);

OAI21x1_ASAP7_75t_L g2476 ( 
.A1(n_2291),
.A2(n_628),
.B(n_625),
.Y(n_2476)
);

AOI21xp5_ASAP7_75t_L g2477 ( 
.A1(n_2223),
.A2(n_631),
.B(n_630),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2339),
.B(n_2318),
.Y(n_2478)
);

AOI21xp5_ASAP7_75t_L g2479 ( 
.A1(n_2227),
.A2(n_638),
.B(n_635),
.Y(n_2479)
);

AOI221xp5_ASAP7_75t_SL g2480 ( 
.A1(n_2364),
.A2(n_1061),
.B1(n_1065),
.B2(n_1054),
.C(n_1051),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2319),
.B(n_1067),
.Y(n_2481)
);

BUFx2_ASAP7_75t_L g2482 ( 
.A(n_2365),
.Y(n_2482)
);

OAI21x1_ASAP7_75t_L g2483 ( 
.A1(n_2291),
.A2(n_642),
.B(n_639),
.Y(n_2483)
);

OAI21x1_ASAP7_75t_L g2484 ( 
.A1(n_2337),
.A2(n_649),
.B(n_645),
.Y(n_2484)
);

AO221x2_ASAP7_75t_L g2485 ( 
.A1(n_2283),
.A2(n_13),
.B1(n_6),
.B2(n_12),
.C(n_14),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_2362),
.B(n_1071),
.Y(n_2486)
);

NAND2x1_ASAP7_75t_L g2487 ( 
.A(n_2337),
.B(n_650),
.Y(n_2487)
);

OAI21x1_ASAP7_75t_L g2488 ( 
.A1(n_2365),
.A2(n_653),
.B(n_652),
.Y(n_2488)
);

AOI221x1_ASAP7_75t_L g2489 ( 
.A1(n_2253),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.C(n_17),
.Y(n_2489)
);

OR2x6_ASAP7_75t_L g2490 ( 
.A(n_2252),
.B(n_654),
.Y(n_2490)
);

INVx3_ASAP7_75t_L g2491 ( 
.A(n_2320),
.Y(n_2491)
);

OAI21x1_ASAP7_75t_L g2492 ( 
.A1(n_2365),
.A2(n_656),
.B(n_655),
.Y(n_2492)
);

AOI21xp5_ASAP7_75t_L g2493 ( 
.A1(n_2227),
.A2(n_658),
.B(n_657),
.Y(n_2493)
);

CKINVDCx11_ASAP7_75t_R g2494 ( 
.A(n_2325),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2289),
.B(n_1073),
.Y(n_2495)
);

OAI21x1_ASAP7_75t_L g2496 ( 
.A1(n_2365),
.A2(n_660),
.B(n_659),
.Y(n_2496)
);

OAI21x1_ASAP7_75t_L g2497 ( 
.A1(n_2241),
.A2(n_665),
.B(n_661),
.Y(n_2497)
);

AND2x4_ASAP7_75t_L g2498 ( 
.A(n_2246),
.B(n_2252),
.Y(n_2498)
);

BUFx6f_ASAP7_75t_L g2499 ( 
.A(n_2325),
.Y(n_2499)
);

OAI21x1_ASAP7_75t_L g2500 ( 
.A1(n_2351),
.A2(n_2309),
.B(n_2347),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2295),
.B(n_2294),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2295),
.B(n_1075),
.Y(n_2502)
);

AOI21xp5_ASAP7_75t_L g2503 ( 
.A1(n_2246),
.A2(n_667),
.B(n_666),
.Y(n_2503)
);

AOI21xp5_ASAP7_75t_L g2504 ( 
.A1(n_2276),
.A2(n_669),
.B(n_668),
.Y(n_2504)
);

AOI21xp5_ASAP7_75t_L g2505 ( 
.A1(n_2276),
.A2(n_671),
.B(n_670),
.Y(n_2505)
);

AOI21xp5_ASAP7_75t_L g2506 ( 
.A1(n_2320),
.A2(n_674),
.B(n_673),
.Y(n_2506)
);

AOI21xp5_ASAP7_75t_L g2507 ( 
.A1(n_2325),
.A2(n_678),
.B(n_675),
.Y(n_2507)
);

OA22x2_ASAP7_75t_L g2508 ( 
.A1(n_2290),
.A2(n_1077),
.B1(n_1078),
.B2(n_1076),
.Y(n_2508)
);

AO31x2_ASAP7_75t_L g2509 ( 
.A1(n_2222),
.A2(n_683),
.A3(n_684),
.B(n_680),
.Y(n_2509)
);

OAI22xp5_ASAP7_75t_L g2510 ( 
.A1(n_2341),
.A2(n_1084),
.B1(n_1085),
.B2(n_1083),
.Y(n_2510)
);

AO31x2_ASAP7_75t_L g2511 ( 
.A1(n_2292),
.A2(n_690),
.A3(n_692),
.B(n_686),
.Y(n_2511)
);

OAI22x1_ASAP7_75t_L g2512 ( 
.A1(n_2349),
.A2(n_1090),
.B1(n_1095),
.B2(n_1088),
.Y(n_2512)
);

OAI21x1_ASAP7_75t_L g2513 ( 
.A1(n_2257),
.A2(n_695),
.B(n_694),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2220),
.B(n_1096),
.Y(n_2514)
);

AND2x4_ASAP7_75t_L g2515 ( 
.A(n_2280),
.B(n_696),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2350),
.B(n_1099),
.Y(n_2516)
);

OAI21xp5_ASAP7_75t_L g2517 ( 
.A1(n_2228),
.A2(n_1269),
.B(n_1267),
.Y(n_2517)
);

NOR2xp67_ASAP7_75t_L g2518 ( 
.A(n_2442),
.B(n_697),
.Y(n_2518)
);

INVx2_ASAP7_75t_L g2519 ( 
.A(n_2397),
.Y(n_2519)
);

INVx6_ASAP7_75t_L g2520 ( 
.A(n_2374),
.Y(n_2520)
);

AND2x2_ASAP7_75t_L g2521 ( 
.A(n_2411),
.B(n_2379),
.Y(n_2521)
);

OAI21x1_ASAP7_75t_L g2522 ( 
.A1(n_2409),
.A2(n_704),
.B(n_702),
.Y(n_2522)
);

OAI22xp33_ASAP7_75t_L g2523 ( 
.A1(n_2400),
.A2(n_1285),
.B1(n_1291),
.B2(n_1283),
.Y(n_2523)
);

INVxp67_ASAP7_75t_L g2524 ( 
.A(n_2410),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2443),
.B(n_706),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2382),
.B(n_707),
.Y(n_2526)
);

INVxp67_ASAP7_75t_L g2527 ( 
.A(n_2461),
.Y(n_2527)
);

BUFx3_ASAP7_75t_L g2528 ( 
.A(n_2429),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2406),
.B(n_2384),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2471),
.Y(n_2530)
);

NOR2xp33_ASAP7_75t_SL g2531 ( 
.A(n_2378),
.B(n_1100),
.Y(n_2531)
);

AND2x6_ASAP7_75t_L g2532 ( 
.A(n_2498),
.B(n_711),
.Y(n_2532)
);

O2A1O1Ixp33_ASAP7_75t_L g2533 ( 
.A1(n_2413),
.A2(n_1321),
.B(n_1318),
.C(n_1105),
.Y(n_2533)
);

HB1xp67_ASAP7_75t_L g2534 ( 
.A(n_2474),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2422),
.B(n_1245),
.Y(n_2535)
);

OAI22xp5_ASAP7_75t_L g2536 ( 
.A1(n_2388),
.A2(n_1108),
.B1(n_1111),
.B2(n_1101),
.Y(n_2536)
);

INVx1_ASAP7_75t_SL g2537 ( 
.A(n_2424),
.Y(n_2537)
);

AO21x2_ASAP7_75t_L g2538 ( 
.A1(n_2394),
.A2(n_1122),
.B(n_1116),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2478),
.B(n_1264),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2376),
.Y(n_2540)
);

BUFx6f_ASAP7_75t_L g2541 ( 
.A(n_2494),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2467),
.B(n_1266),
.Y(n_2542)
);

AOI22xp33_ASAP7_75t_L g2543 ( 
.A1(n_2485),
.A2(n_1127),
.B1(n_1128),
.B2(n_1124),
.Y(n_2543)
);

NOR2xp33_ASAP7_75t_L g2544 ( 
.A(n_2444),
.B(n_1130),
.Y(n_2544)
);

BUFx3_ASAP7_75t_L g2545 ( 
.A(n_2435),
.Y(n_2545)
);

AND2x4_ASAP7_75t_L g2546 ( 
.A(n_2374),
.B(n_2451),
.Y(n_2546)
);

AND2x4_ASAP7_75t_L g2547 ( 
.A(n_2374),
.B(n_2472),
.Y(n_2547)
);

NOR2xp33_ASAP7_75t_L g2548 ( 
.A(n_2398),
.B(n_1134),
.Y(n_2548)
);

OAI21xp33_ASAP7_75t_L g2549 ( 
.A1(n_2517),
.A2(n_1303),
.B(n_1301),
.Y(n_2549)
);

INVx3_ASAP7_75t_L g2550 ( 
.A(n_2389),
.Y(n_2550)
);

AND2x2_ASAP7_75t_L g2551 ( 
.A(n_2427),
.B(n_717),
.Y(n_2551)
);

BUFx2_ASAP7_75t_L g2552 ( 
.A(n_2375),
.Y(n_2552)
);

BUFx6f_ASAP7_75t_L g2553 ( 
.A(n_2499),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2428),
.Y(n_2554)
);

O2A1O1Ixp33_ASAP7_75t_SL g2555 ( 
.A1(n_2383),
.A2(n_20),
.B(n_21),
.C(n_19),
.Y(n_2555)
);

INVx4_ASAP7_75t_L g2556 ( 
.A(n_2499),
.Y(n_2556)
);

BUFx2_ASAP7_75t_L g2557 ( 
.A(n_2375),
.Y(n_2557)
);

AOI21xp5_ASAP7_75t_L g2558 ( 
.A1(n_2390),
.A2(n_1137),
.B(n_1136),
.Y(n_2558)
);

AOI22xp33_ASAP7_75t_L g2559 ( 
.A1(n_2485),
.A2(n_1142),
.B1(n_1145),
.B2(n_1140),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_2377),
.B(n_1247),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2380),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2473),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2381),
.Y(n_2563)
);

OA21x2_ASAP7_75t_L g2564 ( 
.A1(n_2373),
.A2(n_2403),
.B(n_2393),
.Y(n_2564)
);

NAND2x1p5_ASAP7_75t_L g2565 ( 
.A(n_2491),
.B(n_2474),
.Y(n_2565)
);

NOR2x1_ASAP7_75t_L g2566 ( 
.A(n_2427),
.B(n_15),
.Y(n_2566)
);

OAI22xp5_ASAP7_75t_L g2567 ( 
.A1(n_2426),
.A2(n_1151),
.B1(n_1153),
.B2(n_1146),
.Y(n_2567)
);

INVx1_ASAP7_75t_SL g2568 ( 
.A(n_2469),
.Y(n_2568)
);

OR2x2_ASAP7_75t_L g2569 ( 
.A(n_2408),
.B(n_19),
.Y(n_2569)
);

OR2x6_ASAP7_75t_L g2570 ( 
.A(n_2462),
.B(n_722),
.Y(n_2570)
);

INVx3_ASAP7_75t_L g2571 ( 
.A(n_2401),
.Y(n_2571)
);

BUFx3_ASAP7_75t_L g2572 ( 
.A(n_2450),
.Y(n_2572)
);

HB1xp67_ASAP7_75t_L g2573 ( 
.A(n_2482),
.Y(n_2573)
);

BUFx2_ASAP7_75t_L g2574 ( 
.A(n_2482),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2399),
.B(n_723),
.Y(n_2575)
);

INVx3_ASAP7_75t_L g2576 ( 
.A(n_2438),
.Y(n_2576)
);

BUFx4f_ASAP7_75t_SL g2577 ( 
.A(n_2515),
.Y(n_2577)
);

AOI21xp5_ASAP7_75t_L g2578 ( 
.A1(n_2385),
.A2(n_1159),
.B(n_1154),
.Y(n_2578)
);

OAI22xp5_ASAP7_75t_L g2579 ( 
.A1(n_2405),
.A2(n_1162),
.B1(n_1163),
.B2(n_1161),
.Y(n_2579)
);

OR2x2_ASAP7_75t_L g2580 ( 
.A(n_2386),
.B(n_20),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2386),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2436),
.Y(n_2582)
);

INVx3_ASAP7_75t_SL g2583 ( 
.A(n_2391),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2396),
.B(n_2402),
.Y(n_2584)
);

NAND2x1p5_ASAP7_75t_L g2585 ( 
.A(n_2487),
.B(n_724),
.Y(n_2585)
);

NAND2x1_ASAP7_75t_L g2586 ( 
.A(n_2414),
.B(n_726),
.Y(n_2586)
);

AND2x2_ASAP7_75t_L g2587 ( 
.A(n_2455),
.B(n_733),
.Y(n_2587)
);

OAI21x1_ASAP7_75t_L g2588 ( 
.A1(n_2433),
.A2(n_739),
.B(n_735),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2436),
.Y(n_2589)
);

INVx3_ASAP7_75t_L g2590 ( 
.A(n_2465),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2415),
.B(n_1258),
.Y(n_2591)
);

OAI22xp5_ASAP7_75t_L g2592 ( 
.A1(n_2432),
.A2(n_1167),
.B1(n_1170),
.B2(n_1166),
.Y(n_2592)
);

AOI21xp5_ASAP7_75t_L g2593 ( 
.A1(n_2452),
.A2(n_1176),
.B(n_1174),
.Y(n_2593)
);

AO32x1_ASAP7_75t_L g2594 ( 
.A1(n_2446),
.A2(n_23),
.A3(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_2594)
);

AOI21xp5_ASAP7_75t_L g2595 ( 
.A1(n_2454),
.A2(n_1179),
.B(n_1177),
.Y(n_2595)
);

AND2x4_ASAP7_75t_L g2596 ( 
.A(n_2490),
.B(n_740),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2395),
.B(n_1237),
.Y(n_2597)
);

INVx3_ASAP7_75t_L g2598 ( 
.A(n_2490),
.Y(n_2598)
);

OR2x6_ASAP7_75t_L g2599 ( 
.A(n_2462),
.B(n_2419),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2421),
.Y(n_2600)
);

AND2x6_ASAP7_75t_L g2601 ( 
.A(n_2437),
.B(n_741),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2423),
.Y(n_2602)
);

AND2x2_ASAP7_75t_L g2603 ( 
.A(n_2392),
.B(n_2449),
.Y(n_2603)
);

INVx2_ASAP7_75t_SL g2604 ( 
.A(n_2501),
.Y(n_2604)
);

AND2x4_ASAP7_75t_L g2605 ( 
.A(n_2500),
.B(n_742),
.Y(n_2605)
);

OAI22xp5_ASAP7_75t_L g2606 ( 
.A1(n_2440),
.A2(n_1185),
.B1(n_1189),
.B2(n_1181),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2489),
.B(n_1262),
.Y(n_2607)
);

OR2x2_ASAP7_75t_L g2608 ( 
.A(n_2420),
.B(n_22),
.Y(n_2608)
);

AOI21xp5_ASAP7_75t_L g2609 ( 
.A1(n_2479),
.A2(n_2503),
.B(n_2493),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2416),
.Y(n_2610)
);

NOR2x1_ASAP7_75t_SL g2611 ( 
.A(n_2466),
.B(n_743),
.Y(n_2611)
);

BUFx3_ASAP7_75t_L g2612 ( 
.A(n_2445),
.Y(n_2612)
);

OA22x2_ASAP7_75t_L g2613 ( 
.A1(n_2430),
.A2(n_1193),
.B1(n_1199),
.B2(n_1190),
.Y(n_2613)
);

OAI22xp5_ASAP7_75t_L g2614 ( 
.A1(n_2516),
.A2(n_1202),
.B1(n_1203),
.B2(n_1201),
.Y(n_2614)
);

AOI21xp5_ASAP7_75t_L g2615 ( 
.A1(n_2475),
.A2(n_1208),
.B(n_1205),
.Y(n_2615)
);

OR2x6_ASAP7_75t_SL g2616 ( 
.A(n_2407),
.B(n_1212),
.Y(n_2616)
);

AOI21xp5_ASAP7_75t_L g2617 ( 
.A1(n_2477),
.A2(n_1215),
.B(n_1213),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2416),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2511),
.Y(n_2619)
);

O2A1O1Ixp33_ASAP7_75t_L g2620 ( 
.A1(n_2459),
.A2(n_2417),
.B(n_2458),
.C(n_2456),
.Y(n_2620)
);

AOI21xp5_ASAP7_75t_L g2621 ( 
.A1(n_2470),
.A2(n_1223),
.B(n_1216),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_2480),
.B(n_1254),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2502),
.B(n_1272),
.Y(n_2623)
);

OR2x2_ASAP7_75t_L g2624 ( 
.A(n_2552),
.B(n_2481),
.Y(n_2624)
);

AND2x4_ASAP7_75t_L g2625 ( 
.A(n_2552),
.B(n_2511),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2563),
.Y(n_2626)
);

HB1xp67_ASAP7_75t_L g2627 ( 
.A(n_2557),
.Y(n_2627)
);

A2O1A1Ixp33_ASAP7_75t_L g2628 ( 
.A1(n_2620),
.A2(n_2505),
.B(n_2504),
.C(n_2513),
.Y(n_2628)
);

CKINVDCx5p33_ASAP7_75t_R g2629 ( 
.A(n_2568),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2540),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_L g2631 ( 
.A(n_2521),
.B(n_2448),
.Y(n_2631)
);

NOR2xp67_ASAP7_75t_L g2632 ( 
.A(n_2571),
.B(n_2507),
.Y(n_2632)
);

A2O1A1Ixp33_ASAP7_75t_L g2633 ( 
.A1(n_2533),
.A2(n_2506),
.B(n_2404),
.C(n_2425),
.Y(n_2633)
);

INVxp67_ASAP7_75t_L g2634 ( 
.A(n_2534),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2561),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2529),
.B(n_2486),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2554),
.Y(n_2637)
);

BUFx2_ASAP7_75t_L g2638 ( 
.A(n_2565),
.Y(n_2638)
);

INVx1_ASAP7_75t_SL g2639 ( 
.A(n_2537),
.Y(n_2639)
);

NAND2x1p5_ASAP7_75t_L g2640 ( 
.A(n_2598),
.B(n_2488),
.Y(n_2640)
);

OR2x2_ASAP7_75t_L g2641 ( 
.A(n_2557),
.B(n_2495),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2573),
.Y(n_2642)
);

BUFx6f_ASAP7_75t_L g2643 ( 
.A(n_2528),
.Y(n_2643)
);

HB1xp67_ASAP7_75t_L g2644 ( 
.A(n_2574),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_SL g2645 ( 
.A(n_2518),
.B(n_2523),
.Y(n_2645)
);

AOI211xp5_ASAP7_75t_L g2646 ( 
.A1(n_2536),
.A2(n_2510),
.B(n_2463),
.C(n_2468),
.Y(n_2646)
);

AOI21xp5_ASAP7_75t_L g2647 ( 
.A1(n_2609),
.A2(n_2555),
.B(n_2535),
.Y(n_2647)
);

NOR2xp67_ASAP7_75t_L g2648 ( 
.A(n_2524),
.B(n_2514),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2582),
.B(n_2509),
.Y(n_2649)
);

AOI21x1_ASAP7_75t_SL g2650 ( 
.A1(n_2607),
.A2(n_2508),
.B(n_2512),
.Y(n_2650)
);

OR2x2_ASAP7_75t_L g2651 ( 
.A(n_2574),
.B(n_2509),
.Y(n_2651)
);

HB1xp67_ASAP7_75t_L g2652 ( 
.A(n_2589),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2519),
.Y(n_2653)
);

CKINVDCx11_ASAP7_75t_R g2654 ( 
.A(n_2541),
.Y(n_2654)
);

O2A1O1Ixp33_ASAP7_75t_SL g2655 ( 
.A1(n_2584),
.A2(n_2412),
.B(n_33),
.C(n_42),
.Y(n_2655)
);

AND2x4_ASAP7_75t_L g2656 ( 
.A(n_2547),
.B(n_2546),
.Y(n_2656)
);

A2O1A1Ixp33_ASAP7_75t_SL g2657 ( 
.A1(n_2600),
.A2(n_2418),
.B(n_2431),
.C(n_2497),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2527),
.B(n_1226),
.Y(n_2658)
);

OR2x2_ASAP7_75t_L g2659 ( 
.A(n_2569),
.B(n_2434),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2530),
.Y(n_2660)
);

AND2x2_ASAP7_75t_L g2661 ( 
.A(n_2604),
.B(n_2439),
.Y(n_2661)
);

OR2x2_ASAP7_75t_L g2662 ( 
.A(n_2580),
.B(n_2441),
.Y(n_2662)
);

AND2x2_ASAP7_75t_L g2663 ( 
.A(n_2526),
.B(n_2447),
.Y(n_2663)
);

O2A1O1Ixp5_ASAP7_75t_L g2664 ( 
.A1(n_2578),
.A2(n_2496),
.B(n_2492),
.C(n_2483),
.Y(n_2664)
);

AOI21xp5_ASAP7_75t_L g2665 ( 
.A1(n_2599),
.A2(n_2484),
.B(n_2476),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2612),
.B(n_1227),
.Y(n_2666)
);

NOR2x2_ASAP7_75t_L g2667 ( 
.A(n_2570),
.B(n_1232),
.Y(n_2667)
);

AND2x2_ASAP7_75t_L g2668 ( 
.A(n_2603),
.B(n_2453),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_SL g2669 ( 
.A(n_2605),
.B(n_2525),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2542),
.B(n_1233),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2581),
.Y(n_2671)
);

BUFx3_ASAP7_75t_L g2672 ( 
.A(n_2545),
.Y(n_2672)
);

NOR2xp33_ASAP7_75t_L g2673 ( 
.A(n_2544),
.B(n_1235),
.Y(n_2673)
);

NAND2x1p5_ASAP7_75t_L g2674 ( 
.A(n_2541),
.B(n_2457),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2619),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2562),
.Y(n_2676)
);

AND2x2_ASAP7_75t_L g2677 ( 
.A(n_2575),
.B(n_2460),
.Y(n_2677)
);

AND2x4_ASAP7_75t_L g2678 ( 
.A(n_2599),
.B(n_2464),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2539),
.B(n_1236),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2610),
.Y(n_2680)
);

OA21x2_ASAP7_75t_L g2681 ( 
.A1(n_2618),
.A2(n_2387),
.B(n_1241),
.Y(n_2681)
);

AND2x2_ASAP7_75t_L g2682 ( 
.A(n_2551),
.B(n_24),
.Y(n_2682)
);

OR2x2_ASAP7_75t_L g2683 ( 
.A(n_2608),
.B(n_25),
.Y(n_2683)
);

AND2x4_ASAP7_75t_L g2684 ( 
.A(n_2550),
.B(n_781),
.Y(n_2684)
);

AND2x4_ASAP7_75t_L g2685 ( 
.A(n_2572),
.B(n_786),
.Y(n_2685)
);

AOI21xp5_ASAP7_75t_L g2686 ( 
.A1(n_2538),
.A2(n_1243),
.B(n_1239),
.Y(n_2686)
);

INVx2_ASAP7_75t_L g2687 ( 
.A(n_2602),
.Y(n_2687)
);

AND2x2_ASAP7_75t_L g2688 ( 
.A(n_2590),
.B(n_2566),
.Y(n_2688)
);

O2A1O1Ixp5_ASAP7_75t_L g2689 ( 
.A1(n_2586),
.A2(n_1277),
.B(n_1279),
.C(n_1251),
.Y(n_2689)
);

HB1xp67_ASAP7_75t_L g2690 ( 
.A(n_2520),
.Y(n_2690)
);

A2O1A1Ixp33_ASAP7_75t_L g2691 ( 
.A1(n_2549),
.A2(n_1294),
.B(n_1293),
.C(n_28),
.Y(n_2691)
);

A2O1A1Ixp33_ASAP7_75t_L g2692 ( 
.A1(n_2615),
.A2(n_28),
.B(n_26),
.C(n_27),
.Y(n_2692)
);

AND2x2_ASAP7_75t_L g2693 ( 
.A(n_2576),
.B(n_29),
.Y(n_2693)
);

OAI22xp5_ASAP7_75t_SL g2694 ( 
.A1(n_2543),
.A2(n_34),
.B1(n_30),
.B2(n_32),
.Y(n_2694)
);

AND2x4_ASAP7_75t_L g2695 ( 
.A(n_2556),
.B(n_778),
.Y(n_2695)
);

OR2x2_ASAP7_75t_L g2696 ( 
.A(n_2560),
.B(n_32),
.Y(n_2696)
);

INVx1_ASAP7_75t_SL g2697 ( 
.A(n_2583),
.Y(n_2697)
);

A2O1A1Ixp33_ASAP7_75t_L g2698 ( 
.A1(n_2617),
.A2(n_37),
.B(n_34),
.C(n_35),
.Y(n_2698)
);

O2A1O1Ixp33_ASAP7_75t_L g2699 ( 
.A1(n_2622),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_2699)
);

AND2x2_ASAP7_75t_L g2700 ( 
.A(n_2587),
.B(n_38),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2594),
.Y(n_2701)
);

HB1xp67_ASAP7_75t_L g2702 ( 
.A(n_2652),
.Y(n_2702)
);

INVx2_ASAP7_75t_SL g2703 ( 
.A(n_2643),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2630),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2627),
.B(n_2548),
.Y(n_2705)
);

INVx3_ASAP7_75t_L g2706 ( 
.A(n_2656),
.Y(n_2706)
);

OR2x2_ASAP7_75t_L g2707 ( 
.A(n_2644),
.B(n_2642),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2637),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2635),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2675),
.Y(n_2710)
);

AO21x2_ASAP7_75t_L g2711 ( 
.A1(n_2647),
.A2(n_2611),
.B(n_2591),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2680),
.Y(n_2712)
);

AO21x1_ASAP7_75t_SL g2713 ( 
.A1(n_2649),
.A2(n_2597),
.B(n_2594),
.Y(n_2713)
);

BUFx2_ASAP7_75t_SL g2714 ( 
.A(n_2648),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2626),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2687),
.Y(n_2716)
);

AND2x2_ASAP7_75t_L g2717 ( 
.A(n_2634),
.B(n_2616),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2653),
.Y(n_2718)
);

AO21x1_ASAP7_75t_L g2719 ( 
.A1(n_2699),
.A2(n_2645),
.B(n_2636),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_2656),
.B(n_2570),
.Y(n_2720)
);

AOI21x1_ASAP7_75t_L g2721 ( 
.A1(n_2686),
.A2(n_2558),
.B(n_2621),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2625),
.B(n_2623),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2660),
.Y(n_2723)
);

INVx1_ASAP7_75t_SL g2724 ( 
.A(n_2641),
.Y(n_2724)
);

AND2x2_ASAP7_75t_L g2725 ( 
.A(n_2638),
.B(n_2531),
.Y(n_2725)
);

AO21x2_ASAP7_75t_L g2726 ( 
.A1(n_2665),
.A2(n_2595),
.B(n_2593),
.Y(n_2726)
);

AND2x4_ASAP7_75t_L g2727 ( 
.A(n_2625),
.B(n_2553),
.Y(n_2727)
);

OAI21x1_ASAP7_75t_L g2728 ( 
.A1(n_2664),
.A2(n_2522),
.B(n_2564),
.Y(n_2728)
);

INVx3_ASAP7_75t_L g2729 ( 
.A(n_2643),
.Y(n_2729)
);

BUFx12f_ASAP7_75t_L g2730 ( 
.A(n_2654),
.Y(n_2730)
);

AND2x2_ASAP7_75t_L g2731 ( 
.A(n_2639),
.B(n_2553),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2676),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2671),
.Y(n_2733)
);

BUFx2_ASAP7_75t_L g2734 ( 
.A(n_2690),
.Y(n_2734)
);

BUFx2_ASAP7_75t_SL g2735 ( 
.A(n_2643),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2651),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2624),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_2681),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2659),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2661),
.Y(n_2740)
);

HB1xp67_ASAP7_75t_L g2741 ( 
.A(n_2681),
.Y(n_2741)
);

INVx1_ASAP7_75t_SL g2742 ( 
.A(n_2688),
.Y(n_2742)
);

INVx2_ASAP7_75t_SL g2743 ( 
.A(n_2672),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2662),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2678),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2678),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2668),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2701),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2640),
.Y(n_2749)
);

AOI22xp33_ASAP7_75t_L g2750 ( 
.A1(n_2694),
.A2(n_2559),
.B1(n_2613),
.B2(n_2601),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2631),
.Y(n_2751)
);

AND2x4_ASAP7_75t_L g2752 ( 
.A(n_2663),
.B(n_2532),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2682),
.Y(n_2753)
);

OR2x2_ASAP7_75t_L g2754 ( 
.A(n_2683),
.B(n_2564),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2674),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2696),
.Y(n_2756)
);

CKINVDCx5p33_ASAP7_75t_R g2757 ( 
.A(n_2629),
.Y(n_2757)
);

OAI222xp33_ASAP7_75t_L g2758 ( 
.A1(n_2669),
.A2(n_2577),
.B1(n_2596),
.B2(n_2579),
.C1(n_2606),
.C2(n_2592),
.Y(n_2758)
);

OR2x6_ASAP7_75t_L g2759 ( 
.A(n_2677),
.B(n_2520),
.Y(n_2759)
);

INVx2_ASAP7_75t_L g2760 ( 
.A(n_2693),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2655),
.Y(n_2761)
);

AND2x2_ASAP7_75t_L g2762 ( 
.A(n_2697),
.B(n_2532),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2632),
.Y(n_2763)
);

CKINVDCx11_ASAP7_75t_R g2764 ( 
.A(n_2684),
.Y(n_2764)
);

INVx3_ASAP7_75t_L g2765 ( 
.A(n_2685),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2685),
.Y(n_2766)
);

AND2x2_ASAP7_75t_L g2767 ( 
.A(n_2700),
.B(n_2532),
.Y(n_2767)
);

INVx3_ASAP7_75t_L g2768 ( 
.A(n_2684),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2658),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2666),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2692),
.Y(n_2771)
);

AO31x2_ASAP7_75t_L g2772 ( 
.A1(n_2628),
.A2(n_2633),
.A3(n_2698),
.B(n_2691),
.Y(n_2772)
);

INVx2_ASAP7_75t_L g2773 ( 
.A(n_2695),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2670),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2744),
.Y(n_2775)
);

AND2x2_ASAP7_75t_L g2776 ( 
.A(n_2742),
.B(n_2588),
.Y(n_2776)
);

AND2x2_ASAP7_75t_L g2777 ( 
.A(n_2742),
.B(n_2695),
.Y(n_2777)
);

INVx3_ASAP7_75t_L g2778 ( 
.A(n_2746),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2702),
.Y(n_2779)
);

CKINVDCx5p33_ASAP7_75t_R g2780 ( 
.A(n_2757),
.Y(n_2780)
);

CKINVDCx5p33_ASAP7_75t_R g2781 ( 
.A(n_2757),
.Y(n_2781)
);

AND2x4_ASAP7_75t_L g2782 ( 
.A(n_2749),
.B(n_2601),
.Y(n_2782)
);

BUFx2_ASAP7_75t_L g2783 ( 
.A(n_2727),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2739),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2702),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2724),
.B(n_2679),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2710),
.Y(n_2787)
);

INVx2_ASAP7_75t_L g2788 ( 
.A(n_2712),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2724),
.B(n_2673),
.Y(n_2789)
);

NAND2x1p5_ASAP7_75t_L g2790 ( 
.A(n_2749),
.B(n_2657),
.Y(n_2790)
);

AND2x2_ASAP7_75t_L g2791 ( 
.A(n_2737),
.B(n_2689),
.Y(n_2791)
);

AOI22xp33_ASAP7_75t_L g2792 ( 
.A1(n_2771),
.A2(n_2719),
.B1(n_2750),
.B2(n_2761),
.Y(n_2792)
);

INVx2_ASAP7_75t_SL g2793 ( 
.A(n_2707),
.Y(n_2793)
);

OR2x2_ASAP7_75t_L g2794 ( 
.A(n_2736),
.B(n_2614),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2704),
.Y(n_2795)
);

AND2x2_ASAP7_75t_L g2796 ( 
.A(n_2747),
.B(n_2601),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_2754),
.Y(n_2797)
);

AND2x2_ASAP7_75t_L g2798 ( 
.A(n_2745),
.B(n_40),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2708),
.Y(n_2799)
);

INVx3_ASAP7_75t_L g2800 ( 
.A(n_2727),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2715),
.Y(n_2801)
);

AND2x2_ASAP7_75t_L g2802 ( 
.A(n_2706),
.B(n_2585),
.Y(n_2802)
);

OR2x2_ASAP7_75t_L g2803 ( 
.A(n_2740),
.B(n_2567),
.Y(n_2803)
);

OR2x2_ASAP7_75t_L g2804 ( 
.A(n_2748),
.B(n_40),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2715),
.Y(n_2805)
);

AND2x2_ASAP7_75t_L g2806 ( 
.A(n_2734),
.B(n_41),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2709),
.Y(n_2807)
);

INVx3_ASAP7_75t_L g2808 ( 
.A(n_2706),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2718),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2733),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_2716),
.Y(n_2811)
);

AND2x2_ASAP7_75t_L g2812 ( 
.A(n_2751),
.B(n_41),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_2722),
.B(n_2723),
.Y(n_2813)
);

OAI22xp5_ASAP7_75t_L g2814 ( 
.A1(n_2750),
.A2(n_2646),
.B1(n_2667),
.B2(n_2650),
.Y(n_2814)
);

OR2x2_ASAP7_75t_L g2815 ( 
.A(n_2756),
.B(n_43),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2732),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_L g2817 ( 
.A(n_2722),
.B(n_43),
.Y(n_2817)
);

INVx2_ASAP7_75t_L g2818 ( 
.A(n_2763),
.Y(n_2818)
);

AND2x2_ASAP7_75t_L g2819 ( 
.A(n_2753),
.B(n_44),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2787),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2787),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2791),
.B(n_2705),
.Y(n_2822)
);

BUFx2_ASAP7_75t_L g2823 ( 
.A(n_2800),
.Y(n_2823)
);

AND2x4_ASAP7_75t_L g2824 ( 
.A(n_2800),
.B(n_2755),
.Y(n_2824)
);

BUFx6f_ASAP7_75t_L g2825 ( 
.A(n_2790),
.Y(n_2825)
);

BUFx2_ASAP7_75t_L g2826 ( 
.A(n_2800),
.Y(n_2826)
);

INVx2_ASAP7_75t_L g2827 ( 
.A(n_2788),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2788),
.Y(n_2828)
);

OR2x2_ASAP7_75t_L g2829 ( 
.A(n_2793),
.B(n_2705),
.Y(n_2829)
);

BUFx2_ASAP7_75t_L g2830 ( 
.A(n_2783),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2810),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2791),
.B(n_2770),
.Y(n_2832)
);

OAI22xp5_ASAP7_75t_L g2833 ( 
.A1(n_2792),
.A2(n_2714),
.B1(n_2766),
.B2(n_2752),
.Y(n_2833)
);

AND2x2_ASAP7_75t_L g2834 ( 
.A(n_2808),
.B(n_2759),
.Y(n_2834)
);

AND2x2_ASAP7_75t_L g2835 ( 
.A(n_2777),
.B(n_2759),
.Y(n_2835)
);

AND2x2_ASAP7_75t_L g2836 ( 
.A(n_2777),
.B(n_2759),
.Y(n_2836)
);

AND2x2_ASAP7_75t_L g2837 ( 
.A(n_2808),
.B(n_2729),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2810),
.Y(n_2838)
);

INVx3_ASAP7_75t_L g2839 ( 
.A(n_2808),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2779),
.Y(n_2840)
);

INVx3_ASAP7_75t_L g2841 ( 
.A(n_2778),
.Y(n_2841)
);

AND2x2_ASAP7_75t_L g2842 ( 
.A(n_2797),
.B(n_2729),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2785),
.Y(n_2843)
);

BUFx3_ASAP7_75t_L g2844 ( 
.A(n_2780),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2795),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2818),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2813),
.B(n_2774),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2799),
.Y(n_2848)
);

AND2x2_ASAP7_75t_L g2849 ( 
.A(n_2797),
.B(n_2717),
.Y(n_2849)
);

BUFx12f_ASAP7_75t_L g2850 ( 
.A(n_2780),
.Y(n_2850)
);

CKINVDCx5p33_ASAP7_75t_R g2851 ( 
.A(n_2781),
.Y(n_2851)
);

OAI22xp5_ASAP7_75t_L g2852 ( 
.A1(n_2792),
.A2(n_2814),
.B1(n_2782),
.B2(n_2803),
.Y(n_2852)
);

AND2x2_ASAP7_75t_L g2853 ( 
.A(n_2778),
.B(n_2703),
.Y(n_2853)
);

AND2x2_ASAP7_75t_L g2854 ( 
.A(n_2778),
.B(n_2760),
.Y(n_2854)
);

INVx3_ASAP7_75t_L g2855 ( 
.A(n_2818),
.Y(n_2855)
);

AOI21xp33_ASAP7_75t_L g2856 ( 
.A1(n_2786),
.A2(n_2726),
.B(n_2711),
.Y(n_2856)
);

AND2x2_ASAP7_75t_L g2857 ( 
.A(n_2849),
.B(n_2793),
.Y(n_2857)
);

OR2x2_ASAP7_75t_L g2858 ( 
.A(n_2832),
.B(n_2822),
.Y(n_2858)
);

OR2x2_ASAP7_75t_L g2859 ( 
.A(n_2829),
.B(n_2794),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2845),
.Y(n_2860)
);

AND2x4_ASAP7_75t_L g2861 ( 
.A(n_2849),
.B(n_2782),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_L g2862 ( 
.A(n_2848),
.B(n_2809),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2840),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2843),
.Y(n_2864)
);

AND2x2_ASAP7_75t_L g2865 ( 
.A(n_2835),
.B(n_2796),
.Y(n_2865)
);

NOR2xp67_ASAP7_75t_L g2866 ( 
.A(n_2825),
.B(n_2730),
.Y(n_2866)
);

AND2x2_ASAP7_75t_L g2867 ( 
.A(n_2836),
.B(n_2796),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2820),
.Y(n_2868)
);

AND2x2_ASAP7_75t_L g2869 ( 
.A(n_2830),
.B(n_2776),
.Y(n_2869)
);

NAND2xp5_ASAP7_75t_L g2870 ( 
.A(n_2847),
.B(n_2807),
.Y(n_2870)
);

OR2x2_ASAP7_75t_L g2871 ( 
.A(n_2846),
.B(n_2789),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2821),
.Y(n_2872)
);

AND2x2_ASAP7_75t_L g2873 ( 
.A(n_2834),
.B(n_2842),
.Y(n_2873)
);

AND2x2_ASAP7_75t_L g2874 ( 
.A(n_2834),
.B(n_2776),
.Y(n_2874)
);

AND2x2_ASAP7_75t_L g2875 ( 
.A(n_2842),
.B(n_2782),
.Y(n_2875)
);

INVx2_ASAP7_75t_L g2876 ( 
.A(n_2855),
.Y(n_2876)
);

INVx4_ASAP7_75t_L g2877 ( 
.A(n_2850),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2828),
.B(n_2816),
.Y(n_2878)
);

INVx1_ASAP7_75t_SL g2879 ( 
.A(n_2844),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2831),
.Y(n_2880)
);

OR2x2_ASAP7_75t_L g2881 ( 
.A(n_2846),
.B(n_2775),
.Y(n_2881)
);

HB1xp67_ASAP7_75t_L g2882 ( 
.A(n_2827),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2838),
.B(n_2812),
.Y(n_2883)
);

AND2x2_ASAP7_75t_L g2884 ( 
.A(n_2837),
.B(n_2775),
.Y(n_2884)
);

HB1xp67_ASAP7_75t_L g2885 ( 
.A(n_2827),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2852),
.B(n_2812),
.Y(n_2886)
);

AND2x2_ASAP7_75t_L g2887 ( 
.A(n_2837),
.B(n_2798),
.Y(n_2887)
);

INVx2_ASAP7_75t_L g2888 ( 
.A(n_2855),
.Y(n_2888)
);

INVx2_ASAP7_75t_SL g2889 ( 
.A(n_2844),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2855),
.Y(n_2890)
);

INVx3_ASAP7_75t_L g2891 ( 
.A(n_2839),
.Y(n_2891)
);

HB1xp67_ASAP7_75t_L g2892 ( 
.A(n_2823),
.Y(n_2892)
);

AND2x2_ASAP7_75t_L g2893 ( 
.A(n_2853),
.B(n_2798),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2825),
.B(n_2811),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2883),
.Y(n_2895)
);

OAI31xp33_ASAP7_75t_SL g2896 ( 
.A1(n_2879),
.A2(n_2833),
.A3(n_2856),
.B(n_2806),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2883),
.Y(n_2897)
);

HB1xp67_ASAP7_75t_L g2898 ( 
.A(n_2892),
.Y(n_2898)
);

HB1xp67_ASAP7_75t_L g2899 ( 
.A(n_2892),
.Y(n_2899)
);

OR2x2_ASAP7_75t_SL g2900 ( 
.A(n_2886),
.B(n_2825),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2860),
.Y(n_2901)
);

OR2x2_ASAP7_75t_L g2902 ( 
.A(n_2859),
.B(n_2817),
.Y(n_2902)
);

INVx2_ASAP7_75t_L g2903 ( 
.A(n_2889),
.Y(n_2903)
);

NAND3xp33_ASAP7_75t_L g2904 ( 
.A(n_2886),
.B(n_2825),
.C(n_2804),
.Y(n_2904)
);

INVx3_ASAP7_75t_SL g2905 ( 
.A(n_2877),
.Y(n_2905)
);

OR2x2_ASAP7_75t_L g2906 ( 
.A(n_2871),
.B(n_2815),
.Y(n_2906)
);

AND2x2_ASAP7_75t_L g2907 ( 
.A(n_2875),
.B(n_2824),
.Y(n_2907)
);

NAND3xp33_ASAP7_75t_L g2908 ( 
.A(n_2877),
.B(n_2806),
.C(n_2769),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2862),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2862),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2863),
.Y(n_2911)
);

INVxp67_ASAP7_75t_SL g2912 ( 
.A(n_2866),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_2887),
.B(n_2819),
.Y(n_2913)
);

AOI22xp33_ASAP7_75t_L g2914 ( 
.A1(n_2861),
.A2(n_2726),
.B1(n_2711),
.B2(n_2752),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2893),
.B(n_2819),
.Y(n_2915)
);

OR2x2_ASAP7_75t_L g2916 ( 
.A(n_2858),
.B(n_2826),
.Y(n_2916)
);

OAI31xp33_ASAP7_75t_L g2917 ( 
.A1(n_2861),
.A2(n_2758),
.A3(n_2790),
.B(n_2762),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_2857),
.B(n_2854),
.Y(n_2918)
);

NOR2xp33_ASAP7_75t_L g2919 ( 
.A(n_2865),
.B(n_2850),
.Y(n_2919)
);

INVx2_ASAP7_75t_L g2920 ( 
.A(n_2873),
.Y(n_2920)
);

AOI221xp5_ASAP7_75t_L g2921 ( 
.A1(n_2864),
.A2(n_2758),
.B1(n_2741),
.B2(n_2824),
.C(n_2805),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2882),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2882),
.Y(n_2923)
);

INVx3_ASAP7_75t_L g2924 ( 
.A(n_2891),
.Y(n_2924)
);

OAI33xp33_ASAP7_75t_L g2925 ( 
.A1(n_2868),
.A2(n_2872),
.A3(n_2880),
.B1(n_2890),
.B2(n_2894),
.B3(n_2878),
.Y(n_2925)
);

AO21x2_ASAP7_75t_L g2926 ( 
.A1(n_2894),
.A2(n_2824),
.B(n_2853),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2885),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2870),
.B(n_2854),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2885),
.Y(n_2929)
);

AND2x2_ASAP7_75t_L g2930 ( 
.A(n_2912),
.B(n_2867),
.Y(n_2930)
);

OR2x2_ASAP7_75t_L g2931 ( 
.A(n_2904),
.B(n_2870),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2924),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_2903),
.B(n_2884),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2898),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2899),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2908),
.B(n_2869),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2908),
.B(n_2874),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2924),
.Y(n_2938)
);

HB1xp67_ASAP7_75t_L g2939 ( 
.A(n_2916),
.Y(n_2939)
);

NOR2x1_ASAP7_75t_L g2940 ( 
.A(n_2904),
.B(n_2919),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_L g2941 ( 
.A(n_2913),
.B(n_2878),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2929),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2922),
.Y(n_2943)
);

INVx2_ASAP7_75t_L g2944 ( 
.A(n_2926),
.Y(n_2944)
);

OR2x2_ASAP7_75t_L g2945 ( 
.A(n_2920),
.B(n_2881),
.Y(n_2945)
);

AND2x2_ASAP7_75t_L g2946 ( 
.A(n_2907),
.B(n_2851),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2923),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2927),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2901),
.Y(n_2949)
);

AND2x2_ASAP7_75t_L g2950 ( 
.A(n_2905),
.B(n_2851),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_SL g2951 ( 
.A(n_2917),
.B(n_2781),
.Y(n_2951)
);

AND2x2_ASAP7_75t_L g2952 ( 
.A(n_2906),
.B(n_2891),
.Y(n_2952)
);

OR2x6_ASAP7_75t_L g2953 ( 
.A(n_2902),
.B(n_2735),
.Y(n_2953)
);

OR2x2_ASAP7_75t_L g2954 ( 
.A(n_2900),
.B(n_2876),
.Y(n_2954)
);

AND2x2_ASAP7_75t_L g2955 ( 
.A(n_2915),
.B(n_2839),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_SL g2956 ( 
.A(n_2896),
.B(n_2839),
.Y(n_2956)
);

NAND4xp25_ASAP7_75t_L g2957 ( 
.A(n_2921),
.B(n_2725),
.C(n_2731),
.D(n_2876),
.Y(n_2957)
);

AND2x2_ASAP7_75t_L g2958 ( 
.A(n_2918),
.B(n_2888),
.Y(n_2958)
);

OR2x2_ASAP7_75t_L g2959 ( 
.A(n_2928),
.B(n_2888),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2911),
.Y(n_2960)
);

NAND2x1p5_ASAP7_75t_L g2961 ( 
.A(n_2909),
.B(n_2768),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_SL g2962 ( 
.A(n_2914),
.B(n_2743),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_2895),
.B(n_2841),
.Y(n_2963)
);

AND2x4_ASAP7_75t_SL g2964 ( 
.A(n_2910),
.B(n_2767),
.Y(n_2964)
);

AND2x2_ASAP7_75t_L g2965 ( 
.A(n_2897),
.B(n_2841),
.Y(n_2965)
);

AND2x2_ASAP7_75t_L g2966 ( 
.A(n_2926),
.B(n_2841),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2925),
.B(n_2811),
.Y(n_2967)
);

AND2x4_ASAP7_75t_L g2968 ( 
.A(n_2912),
.B(n_2720),
.Y(n_2968)
);

NOR2xp67_ASAP7_75t_L g2969 ( 
.A(n_2908),
.B(n_2801),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2898),
.Y(n_2970)
);

AND2x2_ASAP7_75t_L g2971 ( 
.A(n_2912),
.B(n_2802),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2924),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2898),
.Y(n_2973)
);

AND2x4_ASAP7_75t_SL g2974 ( 
.A(n_2903),
.B(n_2768),
.Y(n_2974)
);

INVxp33_ASAP7_75t_L g2975 ( 
.A(n_2919),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2950),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2934),
.Y(n_2977)
);

INVx2_ASAP7_75t_L g2978 ( 
.A(n_2930),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2934),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2939),
.B(n_2935),
.Y(n_2980)
);

INVx1_ASAP7_75t_SL g2981 ( 
.A(n_2946),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2935),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2970),
.Y(n_2983)
);

INVx2_ASAP7_75t_L g2984 ( 
.A(n_2968),
.Y(n_2984)
);

INVx2_ASAP7_75t_L g2985 ( 
.A(n_2968),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2970),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_SL g2987 ( 
.A(n_2969),
.B(n_2940),
.Y(n_2987)
);

INVx2_ASAP7_75t_L g2988 ( 
.A(n_2971),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2973),
.Y(n_2989)
);

AND2x4_ASAP7_75t_SL g2990 ( 
.A(n_2953),
.B(n_2765),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2973),
.Y(n_2991)
);

INVx3_ASAP7_75t_SL g2992 ( 
.A(n_2953),
.Y(n_2992)
);

OR2x2_ASAP7_75t_L g2993 ( 
.A(n_2936),
.B(n_2784),
.Y(n_2993)
);

NAND2xp67_ASAP7_75t_SL g2994 ( 
.A(n_2966),
.B(n_45),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2942),
.Y(n_2995)
);

NOR2xp33_ASAP7_75t_SL g2996 ( 
.A(n_2975),
.B(n_2741),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2932),
.B(n_2784),
.Y(n_2997)
);

INVx2_ASAP7_75t_L g2998 ( 
.A(n_2938),
.Y(n_2998)
);

INVx1_ASAP7_75t_SL g2999 ( 
.A(n_2954),
.Y(n_2999)
);

AND2x2_ASAP7_75t_L g3000 ( 
.A(n_2952),
.B(n_2765),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2942),
.Y(n_3001)
);

BUFx3_ASAP7_75t_L g3002 ( 
.A(n_2972),
.Y(n_3002)
);

INVx2_ASAP7_75t_SL g3003 ( 
.A(n_2974),
.Y(n_3003)
);

AOI22xp5_ASAP7_75t_L g3004 ( 
.A1(n_2951),
.A2(n_2764),
.B1(n_2766),
.B2(n_2773),
.Y(n_3004)
);

HB1xp67_ASAP7_75t_L g3005 ( 
.A(n_2944),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_L g3006 ( 
.A(n_2947),
.B(n_2772),
.Y(n_3006)
);

AND2x2_ASAP7_75t_L g3007 ( 
.A(n_2958),
.B(n_2773),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2943),
.Y(n_3008)
);

AND2x4_ASAP7_75t_SL g3009 ( 
.A(n_2955),
.B(n_2764),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2943),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2948),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2949),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_L g3013 ( 
.A(n_2937),
.B(n_2933),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2931),
.B(n_2772),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_L g3015 ( 
.A(n_2960),
.B(n_2772),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2945),
.Y(n_3016)
);

INVx1_ASAP7_75t_SL g3017 ( 
.A(n_2964),
.Y(n_3017)
);

OR2x2_ASAP7_75t_L g3018 ( 
.A(n_2941),
.B(n_2738),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_2967),
.B(n_2956),
.Y(n_3019)
);

AOI211xp5_ASAP7_75t_L g3020 ( 
.A1(n_2957),
.A2(n_2738),
.B(n_2728),
.C(n_48),
.Y(n_3020)
);

INVx3_ASAP7_75t_L g3021 ( 
.A(n_2961),
.Y(n_3021)
);

OR2x2_ASAP7_75t_L g3022 ( 
.A(n_2959),
.B(n_46),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2963),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_L g3024 ( 
.A(n_2965),
.B(n_46),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_L g3025 ( 
.A(n_2962),
.B(n_47),
.Y(n_3025)
);

INVxp67_ASAP7_75t_SL g3026 ( 
.A(n_2939),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2934),
.Y(n_3027)
);

OR2x2_ASAP7_75t_L g3028 ( 
.A(n_2936),
.B(n_48),
.Y(n_3028)
);

BUFx6f_ASAP7_75t_L g3029 ( 
.A(n_2950),
.Y(n_3029)
);

INVx1_ASAP7_75t_SL g3030 ( 
.A(n_2950),
.Y(n_3030)
);

OAI22xp5_ASAP7_75t_L g3031 ( 
.A1(n_2940),
.A2(n_2721),
.B1(n_2713),
.B2(n_52),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2930),
.B(n_50),
.Y(n_3032)
);

OAI21xp33_ASAP7_75t_L g3033 ( 
.A1(n_2940),
.A2(n_50),
.B(n_51),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2934),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2934),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2950),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2934),
.Y(n_3037)
);

NOR2xp33_ASAP7_75t_L g3038 ( 
.A(n_2975),
.B(n_51),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_SL g3039 ( 
.A(n_2950),
.B(n_52),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2930),
.B(n_54),
.Y(n_3040)
);

OR2x2_ASAP7_75t_L g3041 ( 
.A(n_2936),
.B(n_54),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2934),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_3026),
.B(n_55),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_SL g3044 ( 
.A(n_3029),
.B(n_55),
.Y(n_3044)
);

NOR3xp33_ASAP7_75t_L g3045 ( 
.A(n_3030),
.B(n_56),
.C(n_57),
.Y(n_3045)
);

HB1xp67_ASAP7_75t_L g3046 ( 
.A(n_2999),
.Y(n_3046)
);

NAND2xp33_ASAP7_75t_R g3047 ( 
.A(n_2980),
.B(n_57),
.Y(n_3047)
);

AND2x4_ASAP7_75t_L g3048 ( 
.A(n_2984),
.B(n_58),
.Y(n_3048)
);

AND2x4_ASAP7_75t_L g3049 ( 
.A(n_2985),
.B(n_58),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_3005),
.Y(n_3050)
);

OR2x2_ASAP7_75t_L g3051 ( 
.A(n_2978),
.B(n_60),
.Y(n_3051)
);

NOR3xp33_ASAP7_75t_L g3052 ( 
.A(n_2976),
.B(n_61),
.C(n_62),
.Y(n_3052)
);

AND2x2_ASAP7_75t_L g3053 ( 
.A(n_3029),
.B(n_64),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2977),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_3029),
.Y(n_3055)
);

AND2x2_ASAP7_75t_L g3056 ( 
.A(n_3009),
.B(n_64),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_L g3057 ( 
.A(n_2988),
.B(n_65),
.Y(n_3057)
);

OR2x2_ASAP7_75t_L g3058 ( 
.A(n_3028),
.B(n_65),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_L g3059 ( 
.A(n_3033),
.B(n_66),
.Y(n_3059)
);

INVxp67_ASAP7_75t_SL g3060 ( 
.A(n_2987),
.Y(n_3060)
);

NAND2x1p5_ASAP7_75t_L g3061 ( 
.A(n_3039),
.B(n_66),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_3002),
.B(n_2981),
.Y(n_3062)
);

INVx1_ASAP7_75t_SL g3063 ( 
.A(n_2992),
.Y(n_3063)
);

INVx2_ASAP7_75t_L g3064 ( 
.A(n_3036),
.Y(n_3064)
);

AND2x4_ASAP7_75t_L g3065 ( 
.A(n_3003),
.B(n_67),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2979),
.Y(n_3066)
);

INVx2_ASAP7_75t_L g3067 ( 
.A(n_3021),
.Y(n_3067)
);

OAI21xp33_ASAP7_75t_L g3068 ( 
.A1(n_3019),
.A2(n_67),
.B(n_68),
.Y(n_3068)
);

OR2x2_ASAP7_75t_L g3069 ( 
.A(n_3041),
.B(n_69),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_L g3070 ( 
.A(n_3038),
.B(n_69),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2982),
.Y(n_3071)
);

NAND2xp33_ASAP7_75t_SL g3072 ( 
.A(n_3031),
.B(n_71),
.Y(n_3072)
);

OR2x2_ASAP7_75t_L g3073 ( 
.A(n_3013),
.B(n_71),
.Y(n_3073)
);

INVx2_ASAP7_75t_L g3074 ( 
.A(n_3021),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_2998),
.B(n_72),
.Y(n_3075)
);

AOI211x1_ASAP7_75t_L g3076 ( 
.A1(n_3014),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_3076)
);

NOR3xp33_ASAP7_75t_SL g3077 ( 
.A(n_3016),
.B(n_73),
.C(n_74),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_3017),
.B(n_75),
.Y(n_3078)
);

NOR4xp25_ASAP7_75t_SL g3079 ( 
.A(n_2983),
.B(n_77),
.C(n_75),
.D(n_76),
.Y(n_3079)
);

INVx2_ASAP7_75t_L g3080 ( 
.A(n_2990),
.Y(n_3080)
);

OR2x2_ASAP7_75t_L g3081 ( 
.A(n_3032),
.B(n_3040),
.Y(n_3081)
);

AND2x2_ASAP7_75t_L g3082 ( 
.A(n_3000),
.B(n_76),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_3023),
.B(n_77),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2986),
.Y(n_3084)
);

AND2x2_ASAP7_75t_L g3085 ( 
.A(n_3004),
.B(n_78),
.Y(n_3085)
);

AND2x2_ASAP7_75t_L g3086 ( 
.A(n_3007),
.B(n_78),
.Y(n_3086)
);

INVxp67_ASAP7_75t_L g3087 ( 
.A(n_3025),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_3024),
.B(n_79),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2989),
.Y(n_3089)
);

OR2x6_ASAP7_75t_L g3090 ( 
.A(n_3022),
.B(n_79),
.Y(n_3090)
);

AOI22xp33_ASAP7_75t_L g3091 ( 
.A1(n_2996),
.A2(n_2993),
.B1(n_3027),
.B2(n_2991),
.Y(n_3091)
);

INVx3_ASAP7_75t_L g3092 ( 
.A(n_3034),
.Y(n_3092)
);

AND2x4_ASAP7_75t_SL g3093 ( 
.A(n_3035),
.B(n_80),
.Y(n_3093)
);

AND2x2_ASAP7_75t_L g3094 ( 
.A(n_3037),
.B(n_80),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_3042),
.B(n_81),
.Y(n_3095)
);

AND2x2_ASAP7_75t_L g3096 ( 
.A(n_3011),
.B(n_81),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2995),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_3001),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_3008),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_3010),
.Y(n_3100)
);

AOI22xp33_ASAP7_75t_L g3101 ( 
.A1(n_3012),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_3101)
);

BUFx2_ASAP7_75t_L g3102 ( 
.A(n_2994),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_3020),
.B(n_82),
.Y(n_3103)
);

OR2x2_ASAP7_75t_L g3104 ( 
.A(n_2997),
.B(n_83),
.Y(n_3104)
);

NAND2xp33_ASAP7_75t_SL g3105 ( 
.A(n_3006),
.B(n_84),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_3015),
.B(n_3018),
.Y(n_3106)
);

NOR3xp33_ASAP7_75t_SL g3107 ( 
.A(n_2994),
.B(n_85),
.C(n_86),
.Y(n_3107)
);

AND2x4_ASAP7_75t_SL g3108 ( 
.A(n_3029),
.B(n_86),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_3026),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_3029),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_3026),
.B(n_88),
.Y(n_3111)
);

INVx2_ASAP7_75t_L g3112 ( 
.A(n_3029),
.Y(n_3112)
);

NOR2xp33_ASAP7_75t_L g3113 ( 
.A(n_3029),
.B(n_88),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_3026),
.Y(n_3114)
);

OR2x2_ASAP7_75t_L g3115 ( 
.A(n_2999),
.B(n_89),
.Y(n_3115)
);

INVx2_ASAP7_75t_SL g3116 ( 
.A(n_3029),
.Y(n_3116)
);

INVx3_ASAP7_75t_L g3117 ( 
.A(n_3029),
.Y(n_3117)
);

AND2x2_ASAP7_75t_L g3118 ( 
.A(n_3029),
.B(n_93),
.Y(n_3118)
);

NOR2xp33_ASAP7_75t_R g3119 ( 
.A(n_3029),
.B(n_94),
.Y(n_3119)
);

NAND2x1_ASAP7_75t_L g3120 ( 
.A(n_3021),
.B(n_97),
.Y(n_3120)
);

AND2x2_ASAP7_75t_L g3121 ( 
.A(n_3029),
.B(n_97),
.Y(n_3121)
);

AND2x2_ASAP7_75t_L g3122 ( 
.A(n_3029),
.B(n_98),
.Y(n_3122)
);

INVxp67_ASAP7_75t_L g3123 ( 
.A(n_3026),
.Y(n_3123)
);

INVx2_ASAP7_75t_L g3124 ( 
.A(n_3029),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_3026),
.B(n_98),
.Y(n_3125)
);

NAND2xp33_ASAP7_75t_SL g3126 ( 
.A(n_2987),
.B(n_100),
.Y(n_3126)
);

NAND2xp33_ASAP7_75t_R g3127 ( 
.A(n_2980),
.B(n_101),
.Y(n_3127)
);

AND2x2_ASAP7_75t_L g3128 ( 
.A(n_3029),
.B(n_101),
.Y(n_3128)
);

AND2x2_ASAP7_75t_L g3129 ( 
.A(n_3029),
.B(n_102),
.Y(n_3129)
);

AND2x2_ASAP7_75t_L g3130 ( 
.A(n_3029),
.B(n_102),
.Y(n_3130)
);

AND2x2_ASAP7_75t_L g3131 ( 
.A(n_3029),
.B(n_104),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_L g3132 ( 
.A(n_3026),
.B(n_104),
.Y(n_3132)
);

AOI22xp33_ASAP7_75t_L g3133 ( 
.A1(n_2987),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_3133)
);

AND2x2_ASAP7_75t_L g3134 ( 
.A(n_3029),
.B(n_105),
.Y(n_3134)
);

AND2x2_ASAP7_75t_L g3135 ( 
.A(n_3029),
.B(n_108),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_3116),
.B(n_108),
.Y(n_3136)
);

OR2x2_ASAP7_75t_L g3137 ( 
.A(n_3046),
.B(n_109),
.Y(n_3137)
);

OR2x2_ASAP7_75t_L g3138 ( 
.A(n_3109),
.B(n_109),
.Y(n_3138)
);

HB1xp67_ASAP7_75t_L g3139 ( 
.A(n_3120),
.Y(n_3139)
);

INVx2_ASAP7_75t_L g3140 ( 
.A(n_3120),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_SL g3141 ( 
.A(n_3065),
.B(n_111),
.Y(n_3141)
);

INVxp67_ASAP7_75t_L g3142 ( 
.A(n_3047),
.Y(n_3142)
);

INVxp67_ASAP7_75t_L g3143 ( 
.A(n_3127),
.Y(n_3143)
);

AND2x2_ASAP7_75t_L g3144 ( 
.A(n_3063),
.B(n_111),
.Y(n_3144)
);

INVxp67_ASAP7_75t_L g3145 ( 
.A(n_3102),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_L g3146 ( 
.A(n_3117),
.B(n_112),
.Y(n_3146)
);

BUFx2_ASAP7_75t_L g3147 ( 
.A(n_3119),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_3114),
.Y(n_3148)
);

NOR2x1_ASAP7_75t_L g3149 ( 
.A(n_3115),
.B(n_112),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_L g3150 ( 
.A(n_3065),
.B(n_113),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_3092),
.Y(n_3151)
);

OR2x2_ASAP7_75t_L g3152 ( 
.A(n_3123),
.B(n_113),
.Y(n_3152)
);

HB1xp67_ASAP7_75t_L g3153 ( 
.A(n_3090),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_3055),
.B(n_114),
.Y(n_3154)
);

INVx2_ASAP7_75t_L g3155 ( 
.A(n_3108),
.Y(n_3155)
);

AND2x2_ASAP7_75t_SL g3156 ( 
.A(n_3062),
.B(n_114),
.Y(n_3156)
);

OR2x2_ASAP7_75t_L g3157 ( 
.A(n_3110),
.B(n_116),
.Y(n_3157)
);

AND2x2_ASAP7_75t_L g3158 ( 
.A(n_3112),
.B(n_117),
.Y(n_3158)
);

AND2x2_ASAP7_75t_L g3159 ( 
.A(n_3124),
.B(n_117),
.Y(n_3159)
);

OR2x2_ASAP7_75t_L g3160 ( 
.A(n_3064),
.B(n_118),
.Y(n_3160)
);

INVx2_ASAP7_75t_SL g3161 ( 
.A(n_3093),
.Y(n_3161)
);

AND2x2_ASAP7_75t_L g3162 ( 
.A(n_3080),
.B(n_119),
.Y(n_3162)
);

OR2x2_ASAP7_75t_L g3163 ( 
.A(n_3073),
.B(n_119),
.Y(n_3163)
);

NOR2xp67_ASAP7_75t_SL g3164 ( 
.A(n_3058),
.B(n_120),
.Y(n_3164)
);

NAND2x1_ASAP7_75t_L g3165 ( 
.A(n_3092),
.B(n_121),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_3078),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_L g3167 ( 
.A(n_3060),
.B(n_121),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_3053),
.B(n_122),
.Y(n_3168)
);

AND2x2_ASAP7_75t_L g3169 ( 
.A(n_3067),
.B(n_122),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_L g3170 ( 
.A(n_3118),
.B(n_123),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_3050),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_L g3172 ( 
.A(n_3121),
.B(n_124),
.Y(n_3172)
);

INVx2_ASAP7_75t_SL g3173 ( 
.A(n_3048),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_3122),
.Y(n_3174)
);

BUFx2_ASAP7_75t_SL g3175 ( 
.A(n_3048),
.Y(n_3175)
);

CKINVDCx16_ASAP7_75t_R g3176 ( 
.A(n_3126),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_3128),
.Y(n_3177)
);

AND2x2_ASAP7_75t_L g3178 ( 
.A(n_3074),
.B(n_3085),
.Y(n_3178)
);

AND2x2_ASAP7_75t_L g3179 ( 
.A(n_3082),
.B(n_124),
.Y(n_3179)
);

AND2x2_ASAP7_75t_L g3180 ( 
.A(n_3056),
.B(n_125),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_3129),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_3130),
.Y(n_3182)
);

INVx1_ASAP7_75t_SL g3183 ( 
.A(n_3131),
.Y(n_3183)
);

INVx1_ASAP7_75t_SL g3184 ( 
.A(n_3134),
.Y(n_3184)
);

OR2x2_ASAP7_75t_L g3185 ( 
.A(n_3043),
.B(n_127),
.Y(n_3185)
);

BUFx2_ASAP7_75t_L g3186 ( 
.A(n_3090),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_3135),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_3049),
.B(n_127),
.Y(n_3188)
);

NAND4xp25_ASAP7_75t_L g3189 ( 
.A(n_3091),
.B(n_131),
.C(n_129),
.D(n_130),
.Y(n_3189)
);

AND2x4_ASAP7_75t_L g3190 ( 
.A(n_3049),
.B(n_129),
.Y(n_3190)
);

BUFx2_ASAP7_75t_L g3191 ( 
.A(n_3061),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_3051),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_L g3193 ( 
.A(n_3076),
.B(n_132),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_3094),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_3113),
.B(n_133),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_3104),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_3096),
.Y(n_3197)
);

AND2x2_ASAP7_75t_L g3198 ( 
.A(n_3086),
.B(n_134),
.Y(n_3198)
);

NOR2x1_ASAP7_75t_L g3199 ( 
.A(n_3044),
.B(n_134),
.Y(n_3199)
);

INVx2_ASAP7_75t_L g3200 ( 
.A(n_3069),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_3075),
.Y(n_3201)
);

AND2x4_ASAP7_75t_SL g3202 ( 
.A(n_3107),
.B(n_135),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_3045),
.B(n_135),
.Y(n_3203)
);

NOR2x1_ASAP7_75t_L g3204 ( 
.A(n_3111),
.B(n_136),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_3052),
.B(n_136),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_L g3206 ( 
.A(n_3133),
.B(n_137),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_3068),
.B(n_138),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_3077),
.B(n_139),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_L g3209 ( 
.A(n_3087),
.B(n_139),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_3125),
.Y(n_3210)
);

INVx1_ASAP7_75t_SL g3211 ( 
.A(n_3105),
.Y(n_3211)
);

OR2x2_ASAP7_75t_L g3212 ( 
.A(n_3132),
.B(n_3081),
.Y(n_3212)
);

AND2x2_ASAP7_75t_L g3213 ( 
.A(n_3057),
.B(n_3088),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_3095),
.Y(n_3214)
);

OR2x6_ASAP7_75t_L g3215 ( 
.A(n_3083),
.B(n_141),
.Y(n_3215)
);

INVx1_ASAP7_75t_SL g3216 ( 
.A(n_3072),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_3054),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_3066),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_3071),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_3079),
.B(n_142),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_3103),
.B(n_143),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_3070),
.B(n_144),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_3059),
.B(n_3084),
.Y(n_3223)
);

AND2x4_ASAP7_75t_L g3224 ( 
.A(n_3099),
.B(n_145),
.Y(n_3224)
);

AND2x2_ASAP7_75t_L g3225 ( 
.A(n_3089),
.B(n_3106),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_3097),
.B(n_145),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_3098),
.Y(n_3227)
);

CKINVDCx20_ASAP7_75t_R g3228 ( 
.A(n_3100),
.Y(n_3228)
);

AND2x2_ASAP7_75t_L g3229 ( 
.A(n_3101),
.B(n_146),
.Y(n_3229)
);

HB1xp67_ASAP7_75t_L g3230 ( 
.A(n_3120),
.Y(n_3230)
);

HB1xp67_ASAP7_75t_L g3231 ( 
.A(n_3120),
.Y(n_3231)
);

AND2x2_ASAP7_75t_L g3232 ( 
.A(n_3063),
.B(n_146),
.Y(n_3232)
);

INVx2_ASAP7_75t_L g3233 ( 
.A(n_3120),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_3046),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_3046),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_L g3236 ( 
.A(n_3116),
.B(n_147),
.Y(n_3236)
);

AND2x2_ASAP7_75t_L g3237 ( 
.A(n_3063),
.B(n_147),
.Y(n_3237)
);

NAND4xp25_ASAP7_75t_L g3238 ( 
.A(n_3063),
.B(n_151),
.C(n_148),
.D(n_150),
.Y(n_3238)
);

NAND3xp33_ASAP7_75t_L g3239 ( 
.A(n_3091),
.B(n_150),
.C(n_151),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_L g3240 ( 
.A(n_3116),
.B(n_152),
.Y(n_3240)
);

NOR3xp33_ASAP7_75t_SL g3241 ( 
.A(n_3062),
.B(n_153),
.C(n_154),
.Y(n_3241)
);

INVx2_ASAP7_75t_L g3242 ( 
.A(n_3120),
.Y(n_3242)
);

AND2x2_ASAP7_75t_L g3243 ( 
.A(n_3063),
.B(n_153),
.Y(n_3243)
);

INVx2_ASAP7_75t_L g3244 ( 
.A(n_3120),
.Y(n_3244)
);

BUFx3_ASAP7_75t_L g3245 ( 
.A(n_3117),
.Y(n_3245)
);

INVx2_ASAP7_75t_SL g3246 ( 
.A(n_3120),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_3046),
.Y(n_3247)
);

CKINVDCx16_ASAP7_75t_R g3248 ( 
.A(n_3047),
.Y(n_3248)
);

NOR2xp33_ASAP7_75t_L g3249 ( 
.A(n_3063),
.B(n_154),
.Y(n_3249)
);

BUFx3_ASAP7_75t_L g3250 ( 
.A(n_3117),
.Y(n_3250)
);

OR2x2_ASAP7_75t_L g3251 ( 
.A(n_3046),
.B(n_155),
.Y(n_3251)
);

NAND2x1_ASAP7_75t_L g3252 ( 
.A(n_3117),
.B(n_155),
.Y(n_3252)
);

NAND2x1p5_ASAP7_75t_L g3253 ( 
.A(n_3120),
.B(n_156),
.Y(n_3253)
);

NAND3xp33_ASAP7_75t_L g3254 ( 
.A(n_3091),
.B(n_157),
.C(n_158),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_3046),
.Y(n_3255)
);

AND2x2_ASAP7_75t_L g3256 ( 
.A(n_3063),
.B(n_158),
.Y(n_3256)
);

AND2x2_ASAP7_75t_L g3257 ( 
.A(n_3063),
.B(n_159),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_3116),
.B(n_159),
.Y(n_3258)
);

OR2x2_ASAP7_75t_L g3259 ( 
.A(n_3046),
.B(n_160),
.Y(n_3259)
);

NOR2xp33_ASAP7_75t_L g3260 ( 
.A(n_3063),
.B(n_161),
.Y(n_3260)
);

AND2x2_ASAP7_75t_L g3261 ( 
.A(n_3063),
.B(n_161),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3046),
.Y(n_3262)
);

OR2x2_ASAP7_75t_L g3263 ( 
.A(n_3046),
.B(n_162),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_3046),
.Y(n_3264)
);

INVx3_ASAP7_75t_L g3265 ( 
.A(n_3117),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3046),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_3046),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_3046),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_3046),
.Y(n_3269)
);

INVx2_ASAP7_75t_SL g3270 ( 
.A(n_3120),
.Y(n_3270)
);

INVx2_ASAP7_75t_L g3271 ( 
.A(n_3120),
.Y(n_3271)
);

INVx2_ASAP7_75t_SL g3272 ( 
.A(n_3120),
.Y(n_3272)
);

AND2x4_ASAP7_75t_L g3273 ( 
.A(n_3116),
.B(n_163),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_SL g3274 ( 
.A(n_3065),
.B(n_163),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_3046),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_3046),
.Y(n_3276)
);

INVx3_ASAP7_75t_L g3277 ( 
.A(n_3117),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3046),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_3046),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_L g3280 ( 
.A(n_3116),
.B(n_164),
.Y(n_3280)
);

AND2x2_ASAP7_75t_L g3281 ( 
.A(n_3063),
.B(n_164),
.Y(n_3281)
);

INVx1_ASAP7_75t_SL g3282 ( 
.A(n_3119),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_3046),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_3046),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3046),
.Y(n_3285)
);

NAND2x1_ASAP7_75t_L g3286 ( 
.A(n_3117),
.B(n_165),
.Y(n_3286)
);

AOI22xp33_ASAP7_75t_L g3287 ( 
.A1(n_3060),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.Y(n_3287)
);

INVx2_ASAP7_75t_L g3288 ( 
.A(n_3120),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_L g3289 ( 
.A(n_3116),
.B(n_167),
.Y(n_3289)
);

NOR2x1_ASAP7_75t_L g3290 ( 
.A(n_3120),
.B(n_168),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_3116),
.B(n_169),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_3139),
.Y(n_3292)
);

AOI22xp5_ASAP7_75t_L g3293 ( 
.A1(n_3248),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_3293)
);

NOR3xp33_ASAP7_75t_SL g3294 ( 
.A(n_3176),
.B(n_171),
.C(n_173),
.Y(n_3294)
);

AOI211xp5_ASAP7_75t_L g3295 ( 
.A1(n_3239),
.A2(n_177),
.B(n_174),
.C(n_176),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_3246),
.B(n_179),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_3230),
.Y(n_3297)
);

INVx3_ASAP7_75t_L g3298 ( 
.A(n_3140),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_3231),
.Y(n_3299)
);

INVx1_ASAP7_75t_SL g3300 ( 
.A(n_3175),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_3153),
.Y(n_3301)
);

AOI322xp5_ASAP7_75t_L g3302 ( 
.A1(n_3142),
.A2(n_185),
.A3(n_183),
.B1(n_181),
.B2(n_179),
.C1(n_180),
.C2(n_182),
.Y(n_3302)
);

AOI22xp5_ASAP7_75t_L g3303 ( 
.A1(n_3216),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3186),
.Y(n_3304)
);

NAND2xp5_ASAP7_75t_L g3305 ( 
.A(n_3270),
.B(n_186),
.Y(n_3305)
);

OR2x2_ASAP7_75t_L g3306 ( 
.A(n_3173),
.B(n_186),
.Y(n_3306)
);

OAI22xp33_ASAP7_75t_SL g3307 ( 
.A1(n_3272),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_3233),
.B(n_188),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3147),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3165),
.Y(n_3310)
);

INVx1_ASAP7_75t_SL g3311 ( 
.A(n_3156),
.Y(n_3311)
);

OAI21xp5_ASAP7_75t_L g3312 ( 
.A1(n_3143),
.A2(n_189),
.B(n_190),
.Y(n_3312)
);

AND2x4_ASAP7_75t_L g3313 ( 
.A(n_3242),
.B(n_190),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_3165),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_3290),
.Y(n_3315)
);

NAND2x1_ASAP7_75t_L g3316 ( 
.A(n_3244),
.B(n_191),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_3137),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3251),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3259),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_L g3320 ( 
.A(n_3271),
.B(n_192),
.Y(n_3320)
);

AOI221xp5_ASAP7_75t_L g3321 ( 
.A1(n_3145),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.C(n_196),
.Y(n_3321)
);

AOI21xp33_ASAP7_75t_L g3322 ( 
.A1(n_3211),
.A2(n_193),
.B(n_195),
.Y(n_3322)
);

INVx1_ASAP7_75t_SL g3323 ( 
.A(n_3282),
.Y(n_3323)
);

OAI22xp33_ASAP7_75t_SL g3324 ( 
.A1(n_3288),
.A2(n_199),
.B1(n_196),
.B2(n_198),
.Y(n_3324)
);

XNOR2xp5_ASAP7_75t_L g3325 ( 
.A(n_3202),
.B(n_199),
.Y(n_3325)
);

AOI321xp33_ASAP7_75t_L g3326 ( 
.A1(n_3234),
.A2(n_202),
.A3(n_206),
.B1(n_200),
.B2(n_201),
.C(n_203),
.Y(n_3326)
);

A2O1A1Ixp33_ASAP7_75t_L g3327 ( 
.A1(n_3241),
.A2(n_203),
.B(n_200),
.C(n_201),
.Y(n_3327)
);

OAI322xp33_ASAP7_75t_L g3328 ( 
.A1(n_3235),
.A2(n_206),
.A3(n_208),
.B1(n_209),
.B2(n_210),
.C1(n_211),
.C2(n_214),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3263),
.Y(n_3329)
);

O2A1O1Ixp33_ASAP7_75t_L g3330 ( 
.A1(n_3220),
.A2(n_215),
.B(n_208),
.C(n_211),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3144),
.Y(n_3331)
);

OAI21xp33_ASAP7_75t_L g3332 ( 
.A1(n_3247),
.A2(n_216),
.B(n_217),
.Y(n_3332)
);

OAI21xp33_ASAP7_75t_L g3333 ( 
.A1(n_3255),
.A2(n_216),
.B(n_217),
.Y(n_3333)
);

INVx2_ASAP7_75t_L g3334 ( 
.A(n_3253),
.Y(n_3334)
);

OAI21xp5_ASAP7_75t_L g3335 ( 
.A1(n_3254),
.A2(n_218),
.B(n_219),
.Y(n_3335)
);

OR2x2_ASAP7_75t_L g3336 ( 
.A(n_3189),
.B(n_218),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3232),
.Y(n_3337)
);

AOI32xp33_ASAP7_75t_L g3338 ( 
.A1(n_3262),
.A2(n_221),
.A3(n_219),
.B1(n_220),
.B2(n_222),
.Y(n_3338)
);

AOI22xp5_ASAP7_75t_L g3339 ( 
.A1(n_3228),
.A2(n_224),
.B1(n_221),
.B2(n_223),
.Y(n_3339)
);

NAND3xp33_ASAP7_75t_L g3340 ( 
.A(n_3264),
.B(n_223),
.C(n_224),
.Y(n_3340)
);

INVx2_ASAP7_75t_L g3341 ( 
.A(n_3252),
.Y(n_3341)
);

INVxp67_ASAP7_75t_L g3342 ( 
.A(n_3149),
.Y(n_3342)
);

AOI21xp5_ASAP7_75t_L g3343 ( 
.A1(n_3203),
.A2(n_225),
.B(n_226),
.Y(n_3343)
);

OAI322xp33_ASAP7_75t_L g3344 ( 
.A1(n_3266),
.A2(n_227),
.A3(n_228),
.B1(n_229),
.B2(n_230),
.C1(n_231),
.C2(n_232),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_3237),
.Y(n_3345)
);

HB1xp67_ASAP7_75t_L g3346 ( 
.A(n_3286),
.Y(n_3346)
);

OAI22xp5_ASAP7_75t_L g3347 ( 
.A1(n_3267),
.A2(n_3268),
.B1(n_3275),
.B2(n_3269),
.Y(n_3347)
);

OAI21xp5_ASAP7_75t_L g3348 ( 
.A1(n_3199),
.A2(n_229),
.B(n_232),
.Y(n_3348)
);

OAI222xp33_ASAP7_75t_L g3349 ( 
.A1(n_3276),
.A2(n_3284),
.B1(n_3279),
.B2(n_3285),
.C1(n_3283),
.C2(n_3278),
.Y(n_3349)
);

OAI211xp5_ASAP7_75t_SL g3350 ( 
.A1(n_3223),
.A2(n_235),
.B(n_233),
.C(n_234),
.Y(n_3350)
);

AOI221xp5_ASAP7_75t_L g3351 ( 
.A1(n_3148),
.A2(n_238),
.B1(n_233),
.B2(n_237),
.C(n_240),
.Y(n_3351)
);

OAI21xp33_ASAP7_75t_L g3352 ( 
.A1(n_3245),
.A2(n_237),
.B(n_242),
.Y(n_3352)
);

AOI22xp5_ASAP7_75t_L g3353 ( 
.A1(n_3161),
.A2(n_245),
.B1(n_242),
.B2(n_243),
.Y(n_3353)
);

INVx1_ASAP7_75t_SL g3354 ( 
.A(n_3191),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_3265),
.B(n_243),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_3277),
.B(n_246),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3243),
.Y(n_3357)
);

AND2x2_ASAP7_75t_L g3358 ( 
.A(n_3256),
.B(n_246),
.Y(n_3358)
);

BUFx2_ASAP7_75t_L g3359 ( 
.A(n_3273),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3257),
.Y(n_3360)
);

AOI21xp33_ASAP7_75t_L g3361 ( 
.A1(n_3183),
.A2(n_247),
.B(n_250),
.Y(n_3361)
);

HB1xp67_ASAP7_75t_L g3362 ( 
.A(n_3273),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_3261),
.B(n_250),
.Y(n_3363)
);

AOI21xp5_ASAP7_75t_L g3364 ( 
.A1(n_3193),
.A2(n_251),
.B(n_252),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3281),
.Y(n_3365)
);

OR2x2_ASAP7_75t_L g3366 ( 
.A(n_3184),
.B(n_252),
.Y(n_3366)
);

A2O1A1Ixp33_ASAP7_75t_L g3367 ( 
.A1(n_3167),
.A2(n_258),
.B(n_256),
.C(n_257),
.Y(n_3367)
);

OR2x2_ASAP7_75t_L g3368 ( 
.A(n_3174),
.B(n_256),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_SL g3369 ( 
.A(n_3155),
.B(n_259),
.Y(n_3369)
);

OAI31xp33_ASAP7_75t_L g3370 ( 
.A1(n_3238),
.A2(n_261),
.A3(n_259),
.B(n_260),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_3250),
.Y(n_3371)
);

OAI21xp33_ASAP7_75t_SL g3372 ( 
.A1(n_3151),
.A2(n_261),
.B(n_262),
.Y(n_3372)
);

AND3x1_ASAP7_75t_L g3373 ( 
.A(n_3204),
.B(n_262),
.C(n_263),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3150),
.Y(n_3374)
);

AND2x2_ASAP7_75t_L g3375 ( 
.A(n_3178),
.B(n_264),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_3249),
.B(n_3260),
.Y(n_3376)
);

OAI21xp5_ASAP7_75t_SL g3377 ( 
.A1(n_3177),
.A2(n_264),
.B(n_265),
.Y(n_3377)
);

INVx2_ASAP7_75t_L g3378 ( 
.A(n_3190),
.Y(n_3378)
);

AOI22xp33_ASAP7_75t_L g3379 ( 
.A1(n_3181),
.A2(n_268),
.B1(n_266),
.B2(n_267),
.Y(n_3379)
);

OAI221xp5_ASAP7_75t_SL g3380 ( 
.A1(n_3171),
.A2(n_270),
.B1(n_268),
.B2(n_269),
.C(n_271),
.Y(n_3380)
);

NOR2xp33_ASAP7_75t_SL g3381 ( 
.A(n_3164),
.B(n_271),
.Y(n_3381)
);

OAI22xp5_ASAP7_75t_L g3382 ( 
.A1(n_3287),
.A2(n_3182),
.B1(n_3187),
.B2(n_3197),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_3179),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_3162),
.B(n_272),
.Y(n_3384)
);

AND2x2_ASAP7_75t_L g3385 ( 
.A(n_3194),
.B(n_272),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3190),
.Y(n_3386)
);

O2A1O1Ixp33_ASAP7_75t_L g3387 ( 
.A1(n_3205),
.A2(n_277),
.B(n_274),
.C(n_276),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_L g3388 ( 
.A(n_3169),
.B(n_274),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_3188),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_3198),
.Y(n_3390)
);

OAI22xp5_ASAP7_75t_L g3391 ( 
.A1(n_3208),
.A2(n_278),
.B1(n_276),
.B2(n_277),
.Y(n_3391)
);

AOI21xp33_ASAP7_75t_L g3392 ( 
.A1(n_3212),
.A2(n_278),
.B(n_279),
.Y(n_3392)
);

AOI22xp5_ASAP7_75t_L g3393 ( 
.A1(n_3229),
.A2(n_281),
.B1(n_279),
.B2(n_280),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_3158),
.B(n_3159),
.Y(n_3394)
);

OR2x2_ASAP7_75t_L g3395 ( 
.A(n_3200),
.B(n_280),
.Y(n_3395)
);

OAI21xp5_ASAP7_75t_L g3396 ( 
.A1(n_3141),
.A2(n_281),
.B(n_282),
.Y(n_3396)
);

OAI21xp33_ASAP7_75t_SL g3397 ( 
.A1(n_3192),
.A2(n_282),
.B(n_283),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3180),
.Y(n_3398)
);

OAI22xp5_ASAP7_75t_L g3399 ( 
.A1(n_3166),
.A2(n_287),
.B1(n_284),
.B2(n_286),
.Y(n_3399)
);

INVx1_ASAP7_75t_SL g3400 ( 
.A(n_3274),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_SL g3401 ( 
.A(n_3224),
.B(n_284),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3213),
.B(n_287),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_3168),
.Y(n_3403)
);

OAI21xp33_ASAP7_75t_L g3404 ( 
.A1(n_3210),
.A2(n_288),
.B(n_290),
.Y(n_3404)
);

OR2x2_ASAP7_75t_L g3405 ( 
.A(n_3152),
.B(n_288),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3170),
.Y(n_3406)
);

INVx2_ASAP7_75t_L g3407 ( 
.A(n_3157),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_3172),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_SL g3409 ( 
.A(n_3224),
.B(n_291),
.Y(n_3409)
);

AOI21xp5_ASAP7_75t_L g3410 ( 
.A1(n_3221),
.A2(n_292),
.B(n_293),
.Y(n_3410)
);

OAI33xp33_ASAP7_75t_L g3411 ( 
.A1(n_3217),
.A2(n_292),
.A3(n_294),
.B1(n_295),
.B2(n_296),
.B3(n_297),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_3163),
.Y(n_3412)
);

INVx2_ASAP7_75t_SL g3413 ( 
.A(n_3160),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_3138),
.Y(n_3414)
);

AOI21xp33_ASAP7_75t_L g3415 ( 
.A1(n_3196),
.A2(n_3214),
.B(n_3201),
.Y(n_3415)
);

INVx1_ASAP7_75t_SL g3416 ( 
.A(n_3185),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_3300),
.B(n_3225),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_SL g3418 ( 
.A(n_3373),
.B(n_3341),
.Y(n_3418)
);

OR2x2_ASAP7_75t_L g3419 ( 
.A(n_3359),
.B(n_3136),
.Y(n_3419)
);

NAND2x1_ASAP7_75t_L g3420 ( 
.A(n_3310),
.B(n_3215),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_3362),
.B(n_3236),
.Y(n_3421)
);

AND2x2_ASAP7_75t_L g3422 ( 
.A(n_3311),
.B(n_3215),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3315),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_3298),
.Y(n_3424)
);

NOR2xp33_ASAP7_75t_L g3425 ( 
.A(n_3342),
.B(n_3146),
.Y(n_3425)
);

AND2x2_ASAP7_75t_L g3426 ( 
.A(n_3323),
.B(n_3240),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3298),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_3292),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_3346),
.B(n_3258),
.Y(n_3429)
);

OR2x2_ASAP7_75t_L g3430 ( 
.A(n_3378),
.B(n_3280),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_3314),
.B(n_3289),
.Y(n_3431)
);

INVx5_ASAP7_75t_L g3432 ( 
.A(n_3313),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_3297),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3299),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_3386),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3325),
.B(n_3291),
.Y(n_3436)
);

AND2x2_ASAP7_75t_L g3437 ( 
.A(n_3304),
.B(n_3154),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_L g3438 ( 
.A(n_3334),
.B(n_3222),
.Y(n_3438)
);

AND2x2_ASAP7_75t_L g3439 ( 
.A(n_3301),
.B(n_3218),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3306),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_3313),
.Y(n_3441)
);

NAND2xp33_ASAP7_75t_L g3442 ( 
.A(n_3294),
.B(n_3195),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_3296),
.Y(n_3443)
);

OR2x2_ASAP7_75t_L g3444 ( 
.A(n_3354),
.B(n_3209),
.Y(n_3444)
);

INVx1_ASAP7_75t_SL g3445 ( 
.A(n_3400),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3305),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_3358),
.Y(n_3447)
);

AND2x2_ASAP7_75t_L g3448 ( 
.A(n_3371),
.B(n_3309),
.Y(n_3448)
);

BUFx2_ASAP7_75t_SL g3449 ( 
.A(n_3413),
.Y(n_3449)
);

INVx2_ASAP7_75t_L g3450 ( 
.A(n_3316),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_L g3451 ( 
.A(n_3375),
.B(n_3331),
.Y(n_3451)
);

AND2x4_ASAP7_75t_SL g3452 ( 
.A(n_3398),
.B(n_3219),
.Y(n_3452)
);

AND2x2_ASAP7_75t_L g3453 ( 
.A(n_3337),
.B(n_3227),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_L g3454 ( 
.A(n_3345),
.B(n_3226),
.Y(n_3454)
);

INVx1_ASAP7_75t_SL g3455 ( 
.A(n_3366),
.Y(n_3455)
);

OAI21xp5_ASAP7_75t_SL g3456 ( 
.A1(n_3349),
.A2(n_3347),
.B(n_3330),
.Y(n_3456)
);

NAND2xp33_ASAP7_75t_L g3457 ( 
.A(n_3327),
.B(n_3207),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3308),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_L g3459 ( 
.A(n_3357),
.B(n_3360),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3320),
.Y(n_3460)
);

AND2x2_ASAP7_75t_L g3461 ( 
.A(n_3365),
.B(n_3206),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_3363),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_3383),
.B(n_294),
.Y(n_3463)
);

INVx2_ASAP7_75t_L g3464 ( 
.A(n_3405),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_L g3465 ( 
.A(n_3390),
.B(n_295),
.Y(n_3465)
);

NOR2xp33_ASAP7_75t_L g3466 ( 
.A(n_3381),
.B(n_298),
.Y(n_3466)
);

INVx1_ASAP7_75t_L g3467 ( 
.A(n_3385),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_SL g3468 ( 
.A(n_3307),
.B(n_298),
.Y(n_3468)
);

NOR2xp33_ASAP7_75t_L g3469 ( 
.A(n_3397),
.B(n_299),
.Y(n_3469)
);

NAND3xp33_ASAP7_75t_L g3470 ( 
.A(n_3372),
.B(n_300),
.C(n_301),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_3370),
.B(n_300),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3368),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_SL g3473 ( 
.A(n_3324),
.B(n_301),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3317),
.B(n_302),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3355),
.Y(n_3475)
);

OR2x2_ASAP7_75t_L g3476 ( 
.A(n_3394),
.B(n_3318),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3356),
.Y(n_3477)
);

AND2x2_ASAP7_75t_L g3478 ( 
.A(n_3407),
.B(n_302),
.Y(n_3478)
);

INVxp67_ASAP7_75t_L g3479 ( 
.A(n_3401),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3384),
.Y(n_3480)
);

AND2x2_ASAP7_75t_L g3481 ( 
.A(n_3319),
.B(n_304),
.Y(n_3481)
);

AND2x2_ASAP7_75t_L g3482 ( 
.A(n_3329),
.B(n_304),
.Y(n_3482)
);

HB1xp67_ASAP7_75t_L g3483 ( 
.A(n_3409),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3364),
.B(n_305),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_3338),
.B(n_305),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3395),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3303),
.B(n_306),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_3412),
.B(n_307),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3388),
.Y(n_3489)
);

NOR2x1_ASAP7_75t_L g3490 ( 
.A(n_3340),
.B(n_3377),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3402),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_3369),
.Y(n_3492)
);

A2O1A1Ixp33_ASAP7_75t_L g3493 ( 
.A1(n_3387),
.A2(n_309),
.B(n_307),
.C(n_308),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_L g3494 ( 
.A(n_3416),
.B(n_310),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3414),
.Y(n_3495)
);

AND2x2_ASAP7_75t_L g3496 ( 
.A(n_3348),
.B(n_311),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3410),
.B(n_311),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_3382),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_L g3499 ( 
.A(n_3343),
.B(n_312),
.Y(n_3499)
);

OA21x2_ASAP7_75t_L g3500 ( 
.A1(n_3376),
.A2(n_312),
.B(n_313),
.Y(n_3500)
);

AND2x2_ASAP7_75t_L g3501 ( 
.A(n_3312),
.B(n_313),
.Y(n_3501)
);

NAND2x1_ASAP7_75t_L g3502 ( 
.A(n_3403),
.B(n_314),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_3393),
.B(n_315),
.Y(n_3503)
);

AND2x2_ASAP7_75t_L g3504 ( 
.A(n_3374),
.B(n_316),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3295),
.B(n_316),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_3353),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_3332),
.B(n_317),
.Y(n_3507)
);

INVx2_ASAP7_75t_L g3508 ( 
.A(n_3389),
.Y(n_3508)
);

INVx1_ASAP7_75t_SL g3509 ( 
.A(n_3336),
.Y(n_3509)
);

AND2x2_ASAP7_75t_L g3510 ( 
.A(n_3406),
.B(n_317),
.Y(n_3510)
);

INVx2_ASAP7_75t_SL g3511 ( 
.A(n_3408),
.Y(n_3511)
);

OR2x2_ASAP7_75t_L g3512 ( 
.A(n_3335),
.B(n_3391),
.Y(n_3512)
);

HB1xp67_ASAP7_75t_L g3513 ( 
.A(n_3396),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_3333),
.B(n_318),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_SL g3515 ( 
.A(n_3326),
.B(n_318),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3352),
.Y(n_3516)
);

AND2x2_ASAP7_75t_L g3517 ( 
.A(n_3322),
.B(n_319),
.Y(n_3517)
);

AOI21xp5_ASAP7_75t_L g3518 ( 
.A1(n_3415),
.A2(n_320),
.B(n_321),
.Y(n_3518)
);

INVx1_ASAP7_75t_L g3519 ( 
.A(n_3293),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_3367),
.B(n_320),
.Y(n_3520)
);

INVx3_ASAP7_75t_L g3521 ( 
.A(n_3361),
.Y(n_3521)
);

INVx2_ASAP7_75t_L g3522 ( 
.A(n_3339),
.Y(n_3522)
);

AOI21xp5_ASAP7_75t_L g3523 ( 
.A1(n_3392),
.A2(n_321),
.B(n_322),
.Y(n_3523)
);

NOR2xp33_ASAP7_75t_L g3524 ( 
.A(n_3404),
.B(n_322),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3399),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_3328),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_L g3527 ( 
.A(n_3302),
.B(n_323),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_3344),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_3321),
.B(n_324),
.Y(n_3529)
);

AND2x2_ASAP7_75t_L g3530 ( 
.A(n_3379),
.B(n_3351),
.Y(n_3530)
);

INVxp67_ASAP7_75t_L g3531 ( 
.A(n_3411),
.Y(n_3531)
);

NOR2xp33_ASAP7_75t_L g3532 ( 
.A(n_3350),
.B(n_325),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3380),
.Y(n_3533)
);

AND2x2_ASAP7_75t_L g3534 ( 
.A(n_3300),
.B(n_325),
.Y(n_3534)
);

AND2x2_ASAP7_75t_L g3535 ( 
.A(n_3300),
.B(n_326),
.Y(n_3535)
);

OR2x2_ASAP7_75t_L g3536 ( 
.A(n_3359),
.B(n_326),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3359),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_3359),
.Y(n_3538)
);

INVxp67_ASAP7_75t_L g3539 ( 
.A(n_3362),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_3359),
.Y(n_3540)
);

OR2x2_ASAP7_75t_L g3541 ( 
.A(n_3359),
.B(n_328),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_3359),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_L g3543 ( 
.A(n_3300),
.B(n_329),
.Y(n_3543)
);

AND2x2_ASAP7_75t_L g3544 ( 
.A(n_3300),
.B(n_331),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3359),
.Y(n_3545)
);

INVx2_ASAP7_75t_L g3546 ( 
.A(n_3359),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3359),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_L g3548 ( 
.A(n_3300),
.B(n_331),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_3359),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3359),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3359),
.Y(n_3551)
);

AND2x2_ASAP7_75t_L g3552 ( 
.A(n_3300),
.B(n_332),
.Y(n_3552)
);

AND2x2_ASAP7_75t_L g3553 ( 
.A(n_3300),
.B(n_332),
.Y(n_3553)
);

OR2x2_ASAP7_75t_L g3554 ( 
.A(n_3359),
.B(n_333),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_L g3555 ( 
.A(n_3300),
.B(n_334),
.Y(n_3555)
);

AND2x4_ASAP7_75t_SL g3556 ( 
.A(n_3341),
.B(n_334),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_L g3557 ( 
.A(n_3300),
.B(n_335),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3359),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_3300),
.B(n_335),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3359),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_L g3561 ( 
.A(n_3300),
.B(n_336),
.Y(n_3561)
);

AND2x4_ASAP7_75t_L g3562 ( 
.A(n_3359),
.B(n_337),
.Y(n_3562)
);

AND2x2_ASAP7_75t_L g3563 ( 
.A(n_3300),
.B(n_338),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3359),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3359),
.Y(n_3565)
);

NOR2xp67_ASAP7_75t_SL g3566 ( 
.A(n_3362),
.B(n_338),
.Y(n_3566)
);

AND2x2_ASAP7_75t_L g3567 ( 
.A(n_3300),
.B(n_339),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_3300),
.B(n_339),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_L g3569 ( 
.A(n_3300),
.B(n_340),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_3359),
.Y(n_3570)
);

AND2x2_ASAP7_75t_L g3571 ( 
.A(n_3300),
.B(n_340),
.Y(n_3571)
);

INVx1_ASAP7_75t_SL g3572 ( 
.A(n_3359),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3300),
.B(n_341),
.Y(n_3573)
);

AND2x2_ASAP7_75t_L g3574 ( 
.A(n_3300),
.B(n_342),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3432),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3432),
.Y(n_3576)
);

OR2x2_ASAP7_75t_L g3577 ( 
.A(n_3572),
.B(n_3449),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_SL g3578 ( 
.A(n_3432),
.B(n_342),
.Y(n_3578)
);

OR2x2_ASAP7_75t_L g3579 ( 
.A(n_3540),
.B(n_343),
.Y(n_3579)
);

NOR3xp33_ASAP7_75t_SL g3580 ( 
.A(n_3456),
.B(n_345),
.C(n_346),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_3536),
.Y(n_3581)
);

O2A1O1Ixp33_ASAP7_75t_SL g3582 ( 
.A1(n_3420),
.A2(n_347),
.B(n_345),
.C(n_346),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3541),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3554),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3537),
.Y(n_3585)
);

INVx1_ASAP7_75t_SL g3586 ( 
.A(n_3556),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3538),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3542),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_L g3589 ( 
.A(n_3546),
.B(n_349),
.Y(n_3589)
);

INVx2_ASAP7_75t_L g3590 ( 
.A(n_3450),
.Y(n_3590)
);

INVx1_ASAP7_75t_SL g3591 ( 
.A(n_3422),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_3545),
.B(n_349),
.Y(n_3592)
);

NOR2x1_ASAP7_75t_L g3593 ( 
.A(n_3470),
.B(n_3502),
.Y(n_3593)
);

INVx1_ASAP7_75t_SL g3594 ( 
.A(n_3452),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3547),
.Y(n_3595)
);

XNOR2xp5_ASAP7_75t_L g3596 ( 
.A(n_3445),
.B(n_350),
.Y(n_3596)
);

OAI21xp5_ASAP7_75t_SL g3597 ( 
.A1(n_3539),
.A2(n_351),
.B(n_352),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_SL g3598 ( 
.A(n_3562),
.B(n_351),
.Y(n_3598)
);

NOR2xp33_ASAP7_75t_R g3599 ( 
.A(n_3549),
.B(n_353),
.Y(n_3599)
);

INVxp33_ASAP7_75t_L g3600 ( 
.A(n_3566),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3550),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3551),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_3558),
.Y(n_3603)
);

OAI21xp5_ASAP7_75t_SL g3604 ( 
.A1(n_3560),
.A2(n_353),
.B(n_354),
.Y(n_3604)
);

NOR3xp33_ASAP7_75t_SL g3605 ( 
.A(n_3418),
.B(n_354),
.C(n_356),
.Y(n_3605)
);

NOR3xp33_ASAP7_75t_L g3606 ( 
.A(n_3417),
.B(n_356),
.C(n_357),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3564),
.B(n_359),
.Y(n_3607)
);

HB1xp67_ASAP7_75t_L g3608 ( 
.A(n_3500),
.Y(n_3608)
);

AND2x2_ASAP7_75t_L g3609 ( 
.A(n_3565),
.B(n_359),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_L g3610 ( 
.A(n_3570),
.B(n_3562),
.Y(n_3610)
);

XNOR2xp5_ASAP7_75t_L g3611 ( 
.A(n_3448),
.B(n_360),
.Y(n_3611)
);

AND2x2_ASAP7_75t_L g3612 ( 
.A(n_3534),
.B(n_360),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_3441),
.B(n_362),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3535),
.Y(n_3614)
);

INVxp67_ASAP7_75t_L g3615 ( 
.A(n_3469),
.Y(n_3615)
);

NAND2xp5_ASAP7_75t_L g3616 ( 
.A(n_3544),
.B(n_3552),
.Y(n_3616)
);

INVx2_ASAP7_75t_L g3617 ( 
.A(n_3553),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_L g3618 ( 
.A(n_3563),
.B(n_363),
.Y(n_3618)
);

AOI21xp5_ASAP7_75t_L g3619 ( 
.A1(n_3515),
.A2(n_3442),
.B(n_3421),
.Y(n_3619)
);

XNOR2x2_ASAP7_75t_L g3620 ( 
.A(n_3527),
.B(n_364),
.Y(n_3620)
);

AOI21xp33_ASAP7_75t_L g3621 ( 
.A1(n_3479),
.A2(n_365),
.B(n_366),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_L g3622 ( 
.A(n_3567),
.B(n_367),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3571),
.Y(n_3623)
);

AND2x2_ASAP7_75t_L g3624 ( 
.A(n_3574),
.B(n_368),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_3500),
.Y(n_3625)
);

NOR2xp33_ASAP7_75t_L g3626 ( 
.A(n_3531),
.B(n_368),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_3424),
.B(n_369),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3427),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_L g3629 ( 
.A(n_3435),
.B(n_369),
.Y(n_3629)
);

NOR2xp33_ASAP7_75t_L g3630 ( 
.A(n_3526),
.B(n_3528),
.Y(n_3630)
);

AND2x2_ASAP7_75t_L g3631 ( 
.A(n_3426),
.B(n_370),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3419),
.Y(n_3632)
);

A2O1A1Ixp33_ASAP7_75t_SL g3633 ( 
.A1(n_3498),
.A2(n_373),
.B(n_371),
.C(n_372),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_SL g3634 ( 
.A(n_3455),
.B(n_371),
.Y(n_3634)
);

NAND2xp5_ASAP7_75t_L g3635 ( 
.A(n_3447),
.B(n_372),
.Y(n_3635)
);

OR2x2_ASAP7_75t_L g3636 ( 
.A(n_3543),
.B(n_374),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_SL g3637 ( 
.A(n_3440),
.B(n_375),
.Y(n_3637)
);

INVxp67_ASAP7_75t_SL g3638 ( 
.A(n_3483),
.Y(n_3638)
);

INVxp33_ASAP7_75t_L g3639 ( 
.A(n_3532),
.Y(n_3639)
);

INVx1_ASAP7_75t_SL g3640 ( 
.A(n_3481),
.Y(n_3640)
);

NAND2xp5_ASAP7_75t_SL g3641 ( 
.A(n_3464),
.B(n_375),
.Y(n_3641)
);

AND2x2_ASAP7_75t_L g3642 ( 
.A(n_3437),
.B(n_376),
.Y(n_3642)
);

NAND2xp5_ASAP7_75t_L g3643 ( 
.A(n_3482),
.B(n_377),
.Y(n_3643)
);

NOR2x1_ASAP7_75t_L g3644 ( 
.A(n_3444),
.B(n_379),
.Y(n_3644)
);

AND2x4_ASAP7_75t_L g3645 ( 
.A(n_3478),
.B(n_379),
.Y(n_3645)
);

AND2x2_ASAP7_75t_L g3646 ( 
.A(n_3467),
.B(n_380),
.Y(n_3646)
);

HB1xp67_ASAP7_75t_L g3647 ( 
.A(n_3513),
.Y(n_3647)
);

NAND3xp33_ASAP7_75t_L g3648 ( 
.A(n_3518),
.B(n_381),
.C(n_382),
.Y(n_3648)
);

INVxp67_ASAP7_75t_L g3649 ( 
.A(n_3466),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3548),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3555),
.Y(n_3651)
);

AND2x2_ASAP7_75t_L g3652 ( 
.A(n_3490),
.B(n_381),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_3439),
.B(n_3428),
.Y(n_3653)
);

OR2x2_ASAP7_75t_L g3654 ( 
.A(n_3573),
.B(n_382),
.Y(n_3654)
);

NAND3xp33_ASAP7_75t_SL g3655 ( 
.A(n_3468),
.B(n_384),
.C(n_385),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_3557),
.Y(n_3656)
);

NAND4xp25_ASAP7_75t_L g3657 ( 
.A(n_3533),
.B(n_387),
.C(n_384),
.D(n_386),
.Y(n_3657)
);

HB1xp67_ASAP7_75t_L g3658 ( 
.A(n_3559),
.Y(n_3658)
);

AND2x2_ASAP7_75t_L g3659 ( 
.A(n_3496),
.B(n_388),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3561),
.Y(n_3660)
);

AND2x2_ASAP7_75t_L g3661 ( 
.A(n_3492),
.B(n_388),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3568),
.Y(n_3662)
);

O2A1O1Ixp33_ASAP7_75t_L g3663 ( 
.A1(n_3493),
.A2(n_3473),
.B(n_3520),
.C(n_3457),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_L g3664 ( 
.A(n_3433),
.B(n_389),
.Y(n_3664)
);

NOR2xp33_ASAP7_75t_L g3665 ( 
.A(n_3569),
.B(n_389),
.Y(n_3665)
);

INVxp67_ASAP7_75t_L g3666 ( 
.A(n_3425),
.Y(n_3666)
);

NAND2xp5_ASAP7_75t_L g3667 ( 
.A(n_3434),
.B(n_390),
.Y(n_3667)
);

AND2x2_ASAP7_75t_L g3668 ( 
.A(n_3501),
.B(n_390),
.Y(n_3668)
);

OR2x2_ASAP7_75t_L g3669 ( 
.A(n_3430),
.B(n_391),
.Y(n_3669)
);

AND2x2_ASAP7_75t_L g3670 ( 
.A(n_3461),
.B(n_393),
.Y(n_3670)
);

NOR4xp25_ASAP7_75t_L g3671 ( 
.A(n_3663),
.B(n_3423),
.C(n_3509),
.D(n_3429),
.Y(n_3671)
);

NAND3xp33_ASAP7_75t_L g3672 ( 
.A(n_3605),
.B(n_3525),
.C(n_3516),
.Y(n_3672)
);

NOR3xp33_ASAP7_75t_L g3673 ( 
.A(n_3626),
.B(n_3459),
.C(n_3436),
.Y(n_3673)
);

AOI21xp5_ASAP7_75t_L g3674 ( 
.A1(n_3575),
.A2(n_3431),
.B(n_3451),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_L g3675 ( 
.A(n_3586),
.B(n_3453),
.Y(n_3675)
);

AOI21xp33_ASAP7_75t_SL g3676 ( 
.A1(n_3577),
.A2(n_3476),
.B(n_3472),
.Y(n_3676)
);

NOR3xp33_ASAP7_75t_L g3677 ( 
.A(n_3591),
.B(n_3438),
.C(n_3521),
.Y(n_3677)
);

NOR2xp33_ASAP7_75t_L g3678 ( 
.A(n_3600),
.B(n_3594),
.Y(n_3678)
);

AOI22xp5_ASAP7_75t_L g3679 ( 
.A1(n_3630),
.A2(n_3519),
.B1(n_3506),
.B2(n_3530),
.Y(n_3679)
);

NAND3xp33_ASAP7_75t_SL g3680 ( 
.A(n_3640),
.B(n_3523),
.C(n_3486),
.Y(n_3680)
);

OAI211xp5_ASAP7_75t_SL g3681 ( 
.A1(n_3580),
.A2(n_3615),
.B(n_3619),
.C(n_3666),
.Y(n_3681)
);

NAND4xp25_ASAP7_75t_L g3682 ( 
.A(n_3616),
.B(n_3512),
.C(n_3522),
.D(n_3454),
.Y(n_3682)
);

AND4x1_ASAP7_75t_L g3683 ( 
.A(n_3644),
.B(n_3524),
.C(n_3485),
.D(n_3495),
.Y(n_3683)
);

NAND3xp33_ASAP7_75t_L g3684 ( 
.A(n_3608),
.B(n_3508),
.C(n_3521),
.Y(n_3684)
);

NOR2xp33_ASAP7_75t_SL g3685 ( 
.A(n_3593),
.B(n_3638),
.Y(n_3685)
);

OAI21xp5_ASAP7_75t_L g3686 ( 
.A1(n_3648),
.A2(n_3494),
.B(n_3511),
.Y(n_3686)
);

NAND3xp33_ASAP7_75t_L g3687 ( 
.A(n_3625),
.B(n_3446),
.C(n_3443),
.Y(n_3687)
);

NAND3x1_ASAP7_75t_L g3688 ( 
.A(n_3576),
.B(n_3465),
.C(n_3463),
.Y(n_3688)
);

NAND2xp33_ASAP7_75t_L g3689 ( 
.A(n_3599),
.B(n_3647),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3596),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_L g3691 ( 
.A(n_3590),
.B(n_3504),
.Y(n_3691)
);

AOI21xp5_ASAP7_75t_L g3692 ( 
.A1(n_3578),
.A2(n_3484),
.B(n_3497),
.Y(n_3692)
);

NOR2xp33_ASAP7_75t_L g3693 ( 
.A(n_3610),
.B(n_3471),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_L g3694 ( 
.A(n_3612),
.B(n_3517),
.Y(n_3694)
);

NOR2xp33_ASAP7_75t_L g3695 ( 
.A(n_3639),
.B(n_3499),
.Y(n_3695)
);

NAND3xp33_ASAP7_75t_SL g3696 ( 
.A(n_3606),
.B(n_3488),
.C(n_3474),
.Y(n_3696)
);

NOR2x1_ASAP7_75t_L g3697 ( 
.A(n_3657),
.B(n_3487),
.Y(n_3697)
);

NOR2xp33_ASAP7_75t_L g3698 ( 
.A(n_3604),
.B(n_3507),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3611),
.Y(n_3699)
);

O2A1O1Ixp33_ASAP7_75t_SL g3700 ( 
.A1(n_3633),
.A2(n_3505),
.B(n_3514),
.C(n_3503),
.Y(n_3700)
);

NOR2xp33_ASAP7_75t_L g3701 ( 
.A(n_3614),
.B(n_3529),
.Y(n_3701)
);

NOR3xp33_ASAP7_75t_L g3702 ( 
.A(n_3655),
.B(n_3460),
.C(n_3458),
.Y(n_3702)
);

AOI321xp33_ASAP7_75t_L g3703 ( 
.A1(n_3585),
.A2(n_3491),
.A3(n_3462),
.B1(n_3489),
.B2(n_3480),
.C(n_3477),
.Y(n_3703)
);

NOR2xp33_ASAP7_75t_L g3704 ( 
.A(n_3623),
.B(n_3597),
.Y(n_3704)
);

NAND4xp25_ASAP7_75t_L g3705 ( 
.A(n_3587),
.B(n_3475),
.C(n_3510),
.D(n_396),
.Y(n_3705)
);

NAND4xp75_ASAP7_75t_L g3706 ( 
.A(n_3588),
.B(n_396),
.C(n_393),
.D(n_394),
.Y(n_3706)
);

NOR3xp33_ASAP7_75t_L g3707 ( 
.A(n_3632),
.B(n_394),
.C(n_397),
.Y(n_3707)
);

AOI211xp5_ASAP7_75t_L g3708 ( 
.A1(n_3582),
.A2(n_400),
.B(n_398),
.C(n_399),
.Y(n_3708)
);

NOR2xp33_ASAP7_75t_L g3709 ( 
.A(n_3617),
.B(n_398),
.Y(n_3709)
);

INVx2_ASAP7_75t_L g3710 ( 
.A(n_3645),
.Y(n_3710)
);

NOR3xp33_ASAP7_75t_L g3711 ( 
.A(n_3649),
.B(n_399),
.C(n_400),
.Y(n_3711)
);

O2A1O1Ixp33_ASAP7_75t_L g3712 ( 
.A1(n_3652),
.A2(n_405),
.B(n_401),
.C(n_404),
.Y(n_3712)
);

O2A1O1Ixp33_ASAP7_75t_SL g3713 ( 
.A1(n_3653),
.A2(n_407),
.B(n_401),
.C(n_406),
.Y(n_3713)
);

NAND2xp5_ASAP7_75t_L g3714 ( 
.A(n_3624),
.B(n_406),
.Y(n_3714)
);

OAI21xp33_ASAP7_75t_L g3715 ( 
.A1(n_3595),
.A2(n_407),
.B(n_408),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_3631),
.B(n_408),
.Y(n_3716)
);

INVx2_ASAP7_75t_SL g3717 ( 
.A(n_3645),
.Y(n_3717)
);

O2A1O1Ixp33_ASAP7_75t_L g3718 ( 
.A1(n_3634),
.A2(n_409),
.B(n_410),
.C(n_411),
.Y(n_3718)
);

OAI211xp5_ASAP7_75t_SL g3719 ( 
.A1(n_3601),
.A2(n_409),
.B(n_412),
.C(n_413),
.Y(n_3719)
);

OAI21xp5_ASAP7_75t_L g3720 ( 
.A1(n_3648),
.A2(n_414),
.B(n_415),
.Y(n_3720)
);

NOR2x1_ASAP7_75t_L g3721 ( 
.A(n_3598),
.B(n_415),
.Y(n_3721)
);

AOI211xp5_ASAP7_75t_L g3722 ( 
.A1(n_3602),
.A2(n_416),
.B(n_417),
.C(n_418),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_SL g3723 ( 
.A(n_3581),
.B(n_3583),
.Y(n_3723)
);

NAND2xp5_ASAP7_75t_SL g3724 ( 
.A(n_3584),
.B(n_416),
.Y(n_3724)
);

AOI221x1_ASAP7_75t_L g3725 ( 
.A1(n_3603),
.A2(n_417),
.B1(n_418),
.B2(n_419),
.C(n_420),
.Y(n_3725)
);

OAI21xp5_ASAP7_75t_SL g3726 ( 
.A1(n_3609),
.A2(n_3628),
.B(n_3670),
.Y(n_3726)
);

NAND3xp33_ASAP7_75t_L g3727 ( 
.A(n_3589),
.B(n_419),
.C(n_420),
.Y(n_3727)
);

NAND3xp33_ASAP7_75t_L g3728 ( 
.A(n_3592),
.B(n_421),
.C(n_422),
.Y(n_3728)
);

NOR2xp33_ASAP7_75t_L g3729 ( 
.A(n_3618),
.B(n_421),
.Y(n_3729)
);

INVxp67_ASAP7_75t_L g3730 ( 
.A(n_3642),
.Y(n_3730)
);

O2A1O1Ixp33_ASAP7_75t_L g3731 ( 
.A1(n_3664),
.A2(n_423),
.B(n_424),
.C(n_425),
.Y(n_3731)
);

NAND3xp33_ASAP7_75t_SL g3732 ( 
.A(n_3669),
.B(n_423),
.C(n_424),
.Y(n_3732)
);

NAND3xp33_ASAP7_75t_L g3733 ( 
.A(n_3607),
.B(n_425),
.C(n_426),
.Y(n_3733)
);

AOI22xp33_ASAP7_75t_L g3734 ( 
.A1(n_3677),
.A2(n_3650),
.B1(n_3656),
.B2(n_3651),
.Y(n_3734)
);

OAI22xp33_ASAP7_75t_L g3735 ( 
.A1(n_3685),
.A2(n_3613),
.B1(n_3635),
.B2(n_3579),
.Y(n_3735)
);

OAI211xp5_ASAP7_75t_L g3736 ( 
.A1(n_3679),
.A2(n_3658),
.B(n_3629),
.C(n_3667),
.Y(n_3736)
);

NAND3xp33_ASAP7_75t_L g3737 ( 
.A(n_3708),
.B(n_3627),
.C(n_3660),
.Y(n_3737)
);

AOI21xp33_ASAP7_75t_SL g3738 ( 
.A1(n_3717),
.A2(n_3684),
.B(n_3671),
.Y(n_3738)
);

XNOR2x1_ASAP7_75t_L g3739 ( 
.A(n_3697),
.B(n_3620),
.Y(n_3739)
);

NOR3xp33_ASAP7_75t_L g3740 ( 
.A(n_3681),
.B(n_3662),
.C(n_3641),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3710),
.B(n_3646),
.Y(n_3741)
);

OAI21xp33_ASAP7_75t_L g3742 ( 
.A1(n_3678),
.A2(n_3661),
.B(n_3665),
.Y(n_3742)
);

OAI322xp33_ASAP7_75t_L g3743 ( 
.A1(n_3675),
.A2(n_3637),
.A3(n_3654),
.B1(n_3636),
.B2(n_3622),
.C1(n_3643),
.C2(n_3659),
.Y(n_3743)
);

AOI22xp5_ASAP7_75t_L g3744 ( 
.A1(n_3673),
.A2(n_3668),
.B1(n_3621),
.B2(n_428),
.Y(n_3744)
);

NAND3xp33_ASAP7_75t_SL g3745 ( 
.A(n_3676),
.B(n_426),
.C(n_427),
.Y(n_3745)
);

NOR2x1_ASAP7_75t_L g3746 ( 
.A(n_3706),
.B(n_429),
.Y(n_3746)
);

OAI211xp5_ASAP7_75t_L g3747 ( 
.A1(n_3726),
.A2(n_3686),
.B(n_3674),
.C(n_3721),
.Y(n_3747)
);

NOR3xp33_ASAP7_75t_L g3748 ( 
.A(n_3680),
.B(n_429),
.C(n_430),
.Y(n_3748)
);

AOI211xp5_ASAP7_75t_L g3749 ( 
.A1(n_3689),
.A2(n_431),
.B(n_432),
.C(n_433),
.Y(n_3749)
);

NAND5xp2_ASAP7_75t_L g3750 ( 
.A(n_3703),
.B(n_432),
.C(n_433),
.D(n_437),
.E(n_438),
.Y(n_3750)
);

NOR3xp33_ASAP7_75t_SL g3751 ( 
.A(n_3672),
.B(n_438),
.C(n_440),
.Y(n_3751)
);

NAND2xp5_ASAP7_75t_SL g3752 ( 
.A(n_3720),
.B(n_441),
.Y(n_3752)
);

AOI222xp33_ASAP7_75t_L g3753 ( 
.A1(n_3687),
.A2(n_442),
.B1(n_443),
.B2(n_444),
.C1(n_445),
.C2(n_448),
.Y(n_3753)
);

AOI22xp5_ASAP7_75t_L g3754 ( 
.A1(n_3704),
.A2(n_443),
.B1(n_445),
.B2(n_448),
.Y(n_3754)
);

NOR3xp33_ASAP7_75t_SL g3755 ( 
.A(n_3682),
.B(n_450),
.C(n_451),
.Y(n_3755)
);

NAND4xp25_ASAP7_75t_L g3756 ( 
.A(n_3693),
.B(n_452),
.C(n_453),
.D(n_454),
.Y(n_3756)
);

AOI22xp5_ASAP7_75t_L g3757 ( 
.A1(n_3698),
.A2(n_3690),
.B1(n_3702),
.B2(n_3730),
.Y(n_3757)
);

XNOR2xp5_ASAP7_75t_L g3758 ( 
.A(n_3683),
.B(n_452),
.Y(n_3758)
);

NAND4xp75_ASAP7_75t_L g3759 ( 
.A(n_3723),
.B(n_455),
.C(n_456),
.D(n_457),
.Y(n_3759)
);

AOI22xp33_ASAP7_75t_L g3760 ( 
.A1(n_3699),
.A2(n_458),
.B1(n_459),
.B2(n_460),
.Y(n_3760)
);

BUFx6f_ASAP7_75t_L g3761 ( 
.A(n_3691),
.Y(n_3761)
);

AOI22xp5_ASAP7_75t_L g3762 ( 
.A1(n_3701),
.A2(n_458),
.B1(n_461),
.B2(n_462),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_SL g3763 ( 
.A(n_3712),
.B(n_461),
.Y(n_3763)
);

NAND3xp33_ASAP7_75t_L g3764 ( 
.A(n_3725),
.B(n_462),
.C(n_463),
.Y(n_3764)
);

OAI21xp33_ASAP7_75t_SL g3765 ( 
.A1(n_3705),
.A2(n_465),
.B(n_466),
.Y(n_3765)
);

NOR3x1_ASAP7_75t_L g3766 ( 
.A(n_3732),
.B(n_465),
.C(n_466),
.Y(n_3766)
);

O2A1O1Ixp5_ASAP7_75t_L g3767 ( 
.A1(n_3692),
.A2(n_467),
.B(n_468),
.C(n_471),
.Y(n_3767)
);

O2A1O1Ixp33_ASAP7_75t_SL g3768 ( 
.A1(n_3716),
.A2(n_3724),
.B(n_3714),
.C(n_3694),
.Y(n_3768)
);

NAND3xp33_ASAP7_75t_L g3769 ( 
.A(n_3718),
.B(n_468),
.C(n_471),
.Y(n_3769)
);

NOR2xp67_ASAP7_75t_L g3770 ( 
.A(n_3728),
.B(n_3733),
.Y(n_3770)
);

NOR2xp33_ASAP7_75t_SL g3771 ( 
.A(n_3764),
.B(n_3715),
.Y(n_3771)
);

AOI21xp5_ASAP7_75t_L g3772 ( 
.A1(n_3747),
.A2(n_3700),
.B(n_3713),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3758),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3741),
.Y(n_3774)
);

AOI21xp5_ASAP7_75t_L g3775 ( 
.A1(n_3739),
.A2(n_3731),
.B(n_3696),
.Y(n_3775)
);

AND2x2_ASAP7_75t_L g3776 ( 
.A(n_3755),
.B(n_3729),
.Y(n_3776)
);

AOI22xp5_ASAP7_75t_L g3777 ( 
.A1(n_3740),
.A2(n_3695),
.B1(n_3688),
.B2(n_3707),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3759),
.Y(n_3778)
);

AOI222xp33_ASAP7_75t_L g3779 ( 
.A1(n_3745),
.A2(n_3719),
.B1(n_3727),
.B2(n_3709),
.C1(n_3711),
.C2(n_3722),
.Y(n_3779)
);

AND2x2_ASAP7_75t_L g3780 ( 
.A(n_3751),
.B(n_472),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3746),
.Y(n_3781)
);

AOI221xp5_ASAP7_75t_L g3782 ( 
.A1(n_3738),
.A2(n_473),
.B1(n_474),
.B2(n_476),
.C(n_477),
.Y(n_3782)
);

AOI22xp5_ASAP7_75t_L g3783 ( 
.A1(n_3748),
.A2(n_473),
.B1(n_474),
.B2(n_478),
.Y(n_3783)
);

OAI22xp5_ASAP7_75t_L g3784 ( 
.A1(n_3734),
.A2(n_478),
.B1(n_479),
.B2(n_480),
.Y(n_3784)
);

NOR2xp33_ASAP7_75t_L g3785 ( 
.A(n_3750),
.B(n_480),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_L g3786 ( 
.A(n_3753),
.B(n_481),
.Y(n_3786)
);

NOR2x1_ASAP7_75t_L g3787 ( 
.A(n_3756),
.B(n_482),
.Y(n_3787)
);

OAI221xp5_ASAP7_75t_L g3788 ( 
.A1(n_3757),
.A2(n_482),
.B1(n_483),
.B2(n_484),
.C(n_486),
.Y(n_3788)
);

O2A1O1Ixp33_ASAP7_75t_L g3789 ( 
.A1(n_3767),
.A2(n_483),
.B(n_484),
.C(n_486),
.Y(n_3789)
);

HB1xp67_ASAP7_75t_L g3790 ( 
.A(n_3781),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_L g3791 ( 
.A(n_3785),
.B(n_3749),
.Y(n_3791)
);

AND2x4_ASAP7_75t_L g3792 ( 
.A(n_3774),
.B(n_3761),
.Y(n_3792)
);

AND2x2_ASAP7_75t_L g3793 ( 
.A(n_3780),
.B(n_3766),
.Y(n_3793)
);

AND2x2_ASAP7_75t_L g3794 ( 
.A(n_3776),
.B(n_3761),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_SL g3795 ( 
.A(n_3782),
.B(n_3761),
.Y(n_3795)
);

NOR3x1_ASAP7_75t_L g3796 ( 
.A(n_3788),
.B(n_3769),
.C(n_3737),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3787),
.Y(n_3797)
);

AO22x2_ASAP7_75t_SL g3798 ( 
.A1(n_3773),
.A2(n_3736),
.B1(n_3765),
.B2(n_3742),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3786),
.Y(n_3799)
);

NAND3xp33_ASAP7_75t_SL g3800 ( 
.A(n_3772),
.B(n_3744),
.C(n_3763),
.Y(n_3800)
);

NOR3x1_ASAP7_75t_L g3801 ( 
.A(n_3778),
.B(n_3752),
.C(n_3743),
.Y(n_3801)
);

NOR3x2_ASAP7_75t_L g3802 ( 
.A(n_3777),
.B(n_3735),
.C(n_3768),
.Y(n_3802)
);

NOR2x1_ASAP7_75t_L g3803 ( 
.A(n_3800),
.B(n_3784),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3790),
.B(n_3779),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3798),
.Y(n_3805)
);

INVx2_ASAP7_75t_L g3806 ( 
.A(n_3794),
.Y(n_3806)
);

NAND2xp5_ASAP7_75t_L g3807 ( 
.A(n_3792),
.B(n_3775),
.Y(n_3807)
);

NOR3xp33_ASAP7_75t_L g3808 ( 
.A(n_3795),
.B(n_3789),
.C(n_3770),
.Y(n_3808)
);

NOR2xp33_ASAP7_75t_R g3809 ( 
.A(n_3797),
.B(n_3771),
.Y(n_3809)
);

NOR2x1_ASAP7_75t_L g3810 ( 
.A(n_3793),
.B(n_3754),
.Y(n_3810)
);

AND3x2_ASAP7_75t_L g3811 ( 
.A(n_3799),
.B(n_3791),
.C(n_3802),
.Y(n_3811)
);

AOI211xp5_ASAP7_75t_L g3812 ( 
.A1(n_3801),
.A2(n_3783),
.B(n_3762),
.C(n_3760),
.Y(n_3812)
);

AND2x4_ASAP7_75t_L g3813 ( 
.A(n_3806),
.B(n_3796),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3805),
.Y(n_3814)
);

OA22x2_ASAP7_75t_L g3815 ( 
.A1(n_3811),
.A2(n_487),
.B1(n_488),
.B2(n_489),
.Y(n_3815)
);

XNOR2x1_ASAP7_75t_L g3816 ( 
.A(n_3803),
.B(n_490),
.Y(n_3816)
);

XNOR2xp5_ASAP7_75t_L g3817 ( 
.A(n_3816),
.B(n_3812),
.Y(n_3817)
);

AOI21xp5_ASAP7_75t_L g3818 ( 
.A1(n_3814),
.A2(n_3804),
.B(n_3807),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3815),
.Y(n_3819)
);

OAI211xp5_ASAP7_75t_SL g3820 ( 
.A1(n_3818),
.A2(n_3810),
.B(n_3808),
.C(n_3809),
.Y(n_3820)
);

XNOR2xp5_ASAP7_75t_L g3821 ( 
.A(n_3820),
.B(n_3817),
.Y(n_3821)
);

XNOR2x1_ASAP7_75t_L g3822 ( 
.A(n_3821),
.B(n_3813),
.Y(n_3822)
);

NOR2x1p5_ASAP7_75t_L g3823 ( 
.A(n_3822),
.B(n_3819),
.Y(n_3823)
);

INVx1_ASAP7_75t_L g3824 ( 
.A(n_3823),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_SL g3825 ( 
.A(n_3824),
.B(n_490),
.Y(n_3825)
);

AOI21xp5_ASAP7_75t_L g3826 ( 
.A1(n_3825),
.A2(n_491),
.B(n_492),
.Y(n_3826)
);

INVx2_ASAP7_75t_L g3827 ( 
.A(n_3826),
.Y(n_3827)
);

OR2x6_ASAP7_75t_L g3828 ( 
.A(n_3827),
.B(n_491),
.Y(n_3828)
);

AOI221xp5_ASAP7_75t_L g3829 ( 
.A1(n_3828),
.A2(n_492),
.B1(n_493),
.B2(n_494),
.C(n_496),
.Y(n_3829)
);

AOI211xp5_ASAP7_75t_L g3830 ( 
.A1(n_3829),
.A2(n_493),
.B(n_498),
.C(n_499),
.Y(n_3830)
);


endmodule