module fake_jpeg_5854_n_252 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_252);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx9p33_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_17),
.B(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_42),
.Y(n_71)
);

INVx2_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_14),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_34),
.A2(n_18),
.B1(n_25),
.B2(n_14),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_18),
.B1(n_32),
.B2(n_19),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_32),
.A2(n_23),
.B(n_20),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_51),
.A2(n_25),
.B(n_24),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_53),
.A2(n_43),
.B1(n_45),
.B2(n_36),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_18),
.B1(n_17),
.B2(n_19),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_57),
.A2(n_64),
.B1(n_45),
.B2(n_41),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_58),
.B(n_68),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_66),
.B(n_69),
.C(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_70),
.Y(n_74)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_63),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_37),
.A2(n_26),
.B1(n_11),
.B2(n_23),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_48),
.A2(n_33),
.B1(n_26),
.B2(n_31),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

AO22x1_ASAP7_75t_L g69 ( 
.A1(n_48),
.A2(n_31),
.B1(n_28),
.B2(n_33),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_28),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_76),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_51),
.B1(n_48),
.B2(n_46),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_79),
.B1(n_84),
.B2(n_89),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_33),
.Y(n_109)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_40),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_84),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_59),
.A2(n_43),
.B1(n_41),
.B2(n_49),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_82),
.A2(n_65),
.B1(n_54),
.B2(n_88),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_87),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_43),
.B1(n_40),
.B2(n_37),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_85),
.B(n_56),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_60),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_60),
.A2(n_36),
.B1(n_47),
.B2(n_50),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_66),
.A2(n_47),
.B1(n_31),
.B2(n_28),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_68),
.B1(n_63),
.B2(n_58),
.Y(n_108)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_67),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_54),
.B(n_30),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_92),
.A2(n_93),
.B(n_94),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_87),
.A2(n_61),
.B1(n_47),
.B2(n_56),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_107),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_62),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_104),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_101),
.Y(n_117)
);

AO22x1_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_39),
.B1(n_52),
.B2(n_50),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_SL g113 ( 
.A1(n_102),
.A2(n_110),
.B(n_80),
.C(n_52),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_74),
.B(n_62),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_104),
.A2(n_108),
.B1(n_86),
.B2(n_85),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_74),
.B(n_76),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_105),
.B(n_106),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_75),
.A2(n_89),
.B(n_79),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_77),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_SL g111 ( 
.A1(n_109),
.A2(n_82),
.B(n_90),
.Y(n_111)
);

AO21x2_ASAP7_75t_L g110 ( 
.A1(n_77),
.A2(n_52),
.B(n_50),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_111),
.A2(n_130),
.B1(n_52),
.B2(n_23),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_102),
.B1(n_110),
.B2(n_108),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_97),
.B(n_92),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_114),
.B(n_115),
.Y(n_151)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_118),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_88),
.Y(n_119)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_88),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_120),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_81),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_121),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_81),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_122),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_75),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_125),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_80),
.Y(n_125)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_86),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_55),
.B(n_39),
.Y(n_146)
);

CKINVDCx12_ASAP7_75t_R g130 ( 
.A(n_110),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_103),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_114),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_106),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_137),
.C(n_143),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_98),
.C(n_100),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_140),
.A2(n_141),
.B1(n_144),
.B2(n_122),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_128),
.A2(n_98),
.B1(n_109),
.B2(n_102),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_109),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_110),
.B1(n_91),
.B2(n_50),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_145),
.A2(n_146),
.B(n_112),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_39),
.C(n_20),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_149),
.C(n_152),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_127),
.A2(n_39),
.B1(n_20),
.B2(n_16),
.Y(n_148)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_16),
.C(n_15),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_16),
.C(n_15),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_149),
.B(n_119),
.Y(n_154)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_155),
.A2(n_166),
.B(n_145),
.Y(n_188)
);

AOI22x1_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_126),
.B1(n_113),
.B2(n_130),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_159),
.B1(n_142),
.B2(n_113),
.Y(n_180)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_158),
.Y(n_181)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_L g159 ( 
.A1(n_142),
.A2(n_126),
.B1(n_113),
.B2(n_117),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_146),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_160),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_132),
.B(n_120),
.Y(n_161)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_169),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_164),
.C(n_151),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_121),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_135),
.Y(n_165)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_129),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_173),
.Y(n_176)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_143),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_L g175 ( 
.A1(n_166),
.A2(n_133),
.B(n_147),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_168),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_164),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_180),
.A2(n_188),
.B1(n_156),
.B2(n_174),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_133),
.B1(n_152),
.B2(n_132),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_182),
.A2(n_159),
.B1(n_113),
.B2(n_112),
.Y(n_203)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_191),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_139),
.C(n_117),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_167),
.C(n_179),
.Y(n_196)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_178),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_205),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_196),
.C(n_201),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_200),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_195),
.A2(n_198),
.B1(n_184),
.B2(n_197),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_187),
.A2(n_174),
.B1(n_168),
.B2(n_116),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_163),
.C(n_173),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_204),
.C(n_206),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_171),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_182),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_203),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_15),
.C(n_2),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_1),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_1),
.C(n_3),
.Y(n_206)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_208),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_196),
.A2(n_185),
.B1(n_189),
.B2(n_188),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_210),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_204),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_206),
.B(n_186),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_213),
.A2(n_7),
.B(n_8),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_185),
.C(n_181),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_217),
.C(n_200),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_191),
.C(n_183),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_218),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_224),
.C(n_226),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_220),
.Y(n_230)
);

OAI21x1_ASAP7_75t_SL g222 ( 
.A1(n_216),
.A2(n_3),
.B(n_4),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_222),
.A2(n_223),
.B(n_225),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_217),
.B(n_5),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_214),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_224)
);

AOI21x1_ASAP7_75t_SL g225 ( 
.A1(n_214),
.A2(n_5),
.B(n_6),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_5),
.C(n_6),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_8),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_233),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_207),
.Y(n_232)
);

INVxp33_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_219),
.A2(n_211),
.B(n_215),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_228),
.A2(n_211),
.B(n_9),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_236),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_226),
.A2(n_8),
.B(n_9),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_224),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_239),
.B(n_9),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_235),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_241),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_229),
.B(n_225),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_237),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_244),
.B(n_245),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_10),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_246),
.A2(n_242),
.B(n_10),
.Y(n_248)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_248),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_247),
.A2(n_243),
.B1(n_242),
.B2(n_10),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_249),
.A2(n_250),
.B(n_10),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_67),
.Y(n_252)
);


endmodule