module fake_netlist_1_5704_n_547 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_547);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_547;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_445;
wire n_398;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx3_ASAP7_75t_L g79 ( .A(n_29), .Y(n_79) );
INVxp67_ASAP7_75t_L g80 ( .A(n_78), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_41), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_35), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_60), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_17), .Y(n_84) );
CKINVDCx20_ASAP7_75t_R g85 ( .A(n_32), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_75), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_63), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_12), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_12), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_69), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_77), .Y(n_91) );
CKINVDCx16_ASAP7_75t_R g92 ( .A(n_14), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_62), .Y(n_93) );
BUFx3_ASAP7_75t_L g94 ( .A(n_61), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_45), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_67), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_22), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_46), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_20), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_74), .Y(n_100) );
BUFx3_ASAP7_75t_L g101 ( .A(n_37), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_52), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_10), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_72), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_25), .Y(n_105) );
INVxp33_ASAP7_75t_L g106 ( .A(n_2), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_40), .Y(n_107) );
INVxp33_ASAP7_75t_SL g108 ( .A(n_6), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_11), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_10), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_31), .Y(n_111) );
INVxp33_ASAP7_75t_L g112 ( .A(n_47), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_53), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_64), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_8), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_13), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_81), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_79), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_92), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_81), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_79), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_103), .B(n_0), .Y(n_122) );
INVx3_ASAP7_75t_L g123 ( .A(n_79), .Y(n_123) );
INVxp67_ASAP7_75t_SL g124 ( .A(n_106), .Y(n_124) );
NAND2xp33_ASAP7_75t_L g125 ( .A(n_112), .B(n_76), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_84), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_84), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_110), .B(n_0), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_86), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_89), .B(n_1), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_88), .B(n_1), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_109), .Y(n_132) );
AND2x6_ASAP7_75t_L g133 ( .A(n_94), .B(n_34), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_86), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_89), .B(n_2), .Y(n_135) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_87), .A2(n_36), .B(n_71), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_94), .Y(n_137) );
OR2x2_ASAP7_75t_L g138 ( .A(n_88), .B(n_3), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_87), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_136), .Y(n_140) );
BUFx3_ASAP7_75t_L g141 ( .A(n_133), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_121), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_118), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_123), .B(n_82), .Y(n_144) );
INVx2_ASAP7_75t_SL g145 ( .A(n_123), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_121), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_118), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_117), .B(n_91), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_123), .B(n_115), .Y(n_149) );
BUFx3_ASAP7_75t_L g150 ( .A(n_133), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_121), .Y(n_151) );
INVx4_ASAP7_75t_L g152 ( .A(n_133), .Y(n_152) );
INVx4_ASAP7_75t_L g153 ( .A(n_133), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_123), .B(n_83), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_118), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_118), .Y(n_156) );
INVx4_ASAP7_75t_L g157 ( .A(n_133), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_117), .B(n_97), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_118), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_135), .B(n_120), .Y(n_160) );
OAI22xp5_ASAP7_75t_L g161 ( .A1(n_138), .A2(n_116), .B1(n_110), .B2(n_108), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_120), .B(n_100), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_118), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_137), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g165 ( .A1(n_160), .A2(n_135), .B1(n_130), .B2(n_129), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_160), .B(n_124), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_152), .B(n_135), .Y(n_167) );
INVx5_ASAP7_75t_L g168 ( .A(n_152), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_141), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_148), .B(n_119), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_143), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_160), .B(n_129), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_160), .A2(n_135), .B1(n_130), .B2(n_139), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_160), .B(n_134), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_142), .Y(n_175) );
OR2x2_ASAP7_75t_L g176 ( .A(n_161), .B(n_119), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_141), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_142), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_143), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_161), .B(n_134), .Y(n_180) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_149), .A2(n_139), .B1(n_131), .B2(n_128), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_149), .B(n_138), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_149), .B(n_131), .Y(n_183) );
BUFx3_ASAP7_75t_L g184 ( .A(n_141), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_149), .B(n_91), .Y(n_185) );
INVx3_ASAP7_75t_L g186 ( .A(n_149), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_145), .B(n_93), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_158), .B(n_122), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_143), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_146), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_152), .B(n_93), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_152), .B(n_96), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_158), .B(n_116), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_145), .Y(n_194) );
NAND2x1p5_ASAP7_75t_L g195 ( .A(n_152), .B(n_136), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_153), .B(n_96), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_155), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_180), .A2(n_145), .B1(n_162), .B2(n_154), .Y(n_198) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_193), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_188), .B(n_162), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_175), .Y(n_201) );
NAND3xp33_ASAP7_75t_L g202 ( .A(n_170), .B(n_125), .C(n_144), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_175), .Y(n_203) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_193), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_168), .B(n_153), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_176), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_188), .B(n_146), .Y(n_207) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_178), .A2(n_144), .B(n_154), .Y(n_208) );
BUFx3_ASAP7_75t_L g209 ( .A(n_169), .Y(n_209) );
NAND2xp33_ASAP7_75t_L g210 ( .A(n_168), .B(n_133), .Y(n_210) );
BUFx4f_ASAP7_75t_L g211 ( .A(n_186), .Y(n_211) );
BUFx2_ASAP7_75t_L g212 ( .A(n_186), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_169), .Y(n_213) );
BUFx3_ASAP7_75t_L g214 ( .A(n_169), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_178), .Y(n_215) );
NAND3xp33_ASAP7_75t_L g216 ( .A(n_181), .B(n_157), .C(n_153), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_167), .A2(n_153), .B(n_157), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g218 ( .A1(n_166), .A2(n_172), .B(n_174), .C(n_183), .Y(n_218) );
NOR2x1_ASAP7_75t_L g219 ( .A(n_186), .B(n_151), .Y(n_219) );
BUFx4f_ASAP7_75t_L g220 ( .A(n_186), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_165), .A2(n_85), .B1(n_95), .B2(n_151), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_182), .B(n_153), .Y(n_222) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_184), .Y(n_223) );
BUFx2_ASAP7_75t_L g224 ( .A(n_176), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_182), .B(n_105), .Y(n_225) );
BUFx3_ASAP7_75t_L g226 ( .A(n_184), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_190), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_190), .Y(n_228) );
INVx3_ASAP7_75t_L g229 ( .A(n_184), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_197), .Y(n_230) );
OAI21x1_ASAP7_75t_L g231 ( .A1(n_201), .A2(n_195), .B(n_136), .Y(n_231) );
OAI21x1_ASAP7_75t_L g232 ( .A1(n_201), .A2(n_195), .B(n_136), .Y(n_232) );
OAI21x1_ASAP7_75t_L g233 ( .A1(n_201), .A2(n_195), .B(n_164), .Y(n_233) );
BUFx2_ASAP7_75t_L g234 ( .A(n_207), .Y(n_234) );
AND2x4_ASAP7_75t_SL g235 ( .A(n_207), .B(n_165), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_203), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_203), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_200), .B(n_172), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_203), .B(n_173), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_221), .Y(n_240) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_228), .A2(n_164), .B(n_126), .Y(n_241) );
BUFx12f_ASAP7_75t_L g242 ( .A(n_224), .Y(n_242) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_228), .A2(n_111), .B(n_113), .Y(n_243) );
OAI21x1_ASAP7_75t_L g244 ( .A1(n_215), .A2(n_164), .B(n_163), .Y(n_244) );
OAI21x1_ASAP7_75t_L g245 ( .A1(n_215), .A2(n_155), .B(n_163), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_208), .B(n_173), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_227), .Y(n_247) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_227), .A2(n_111), .B(n_113), .Y(n_248) );
OAI222xp33_ASAP7_75t_L g249 ( .A1(n_224), .A2(n_132), .B1(n_115), .B2(n_90), .C1(n_185), .C2(n_126), .Y(n_249) );
OAI21x1_ASAP7_75t_L g250 ( .A1(n_217), .A2(n_163), .B(n_155), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_208), .B(n_166), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_230), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_230), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_218), .A2(n_126), .B(n_127), .C(n_194), .Y(n_254) );
OAI21x1_ASAP7_75t_L g255 ( .A1(n_230), .A2(n_156), .B(n_159), .Y(n_255) );
AOI21xp33_ASAP7_75t_SL g256 ( .A1(n_206), .A2(n_105), .B(n_114), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_208), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_240), .A2(n_204), .B1(n_199), .B2(n_202), .Y(n_258) );
OAI21x1_ASAP7_75t_L g259 ( .A1(n_233), .A2(n_229), .B(n_205), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_257), .A2(n_210), .B(n_208), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_234), .Y(n_261) );
OAI21xp5_ASAP7_75t_L g262 ( .A1(n_254), .A2(n_198), .B(n_216), .Y(n_262) );
AOI21x1_ASAP7_75t_L g263 ( .A1(n_257), .A2(n_127), .B(n_187), .Y(n_263) );
AOI221xp5_ASAP7_75t_L g264 ( .A1(n_249), .A2(n_225), .B1(n_198), .B2(n_212), .C(n_222), .Y(n_264) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_251), .A2(n_127), .B(n_222), .C(n_219), .Y(n_265) );
AOI221xp5_ASAP7_75t_L g266 ( .A1(n_249), .A2(n_212), .B1(n_211), .B2(n_220), .C(n_90), .Y(n_266) );
OR2x2_ASAP7_75t_L g267 ( .A(n_234), .B(n_114), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g268 ( .A1(n_240), .A2(n_211), .B1(n_220), .B2(n_214), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_234), .B(n_238), .Y(n_269) );
AO21x2_ASAP7_75t_L g270 ( .A1(n_254), .A2(n_107), .B(n_98), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_236), .A2(n_157), .B(n_192), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_237), .Y(n_272) );
AOI22xp33_ASAP7_75t_SL g273 ( .A1(n_242), .A2(n_220), .B1(n_211), .B2(n_209), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_235), .A2(n_219), .B1(n_211), .B2(n_220), .Y(n_274) );
AOI221xp5_ASAP7_75t_L g275 ( .A1(n_238), .A2(n_99), .B1(n_102), .B2(n_104), .C(n_80), .Y(n_275) );
OAI22xp5_ASAP7_75t_L g276 ( .A1(n_235), .A2(n_226), .B1(n_214), .B2(n_209), .Y(n_276) );
OAI221xp5_ASAP7_75t_L g277 ( .A1(n_256), .A2(n_194), .B1(n_229), .B2(n_214), .C(n_226), .Y(n_277) );
OR2x6_ASAP7_75t_L g278 ( .A(n_246), .B(n_213), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_252), .Y(n_279) );
INVx1_ASAP7_75t_SL g280 ( .A(n_242), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_272), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_269), .B(n_246), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_279), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_278), .B(n_237), .Y(n_284) );
BUFx2_ASAP7_75t_L g285 ( .A(n_278), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_279), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_278), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_261), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_278), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_258), .B(n_246), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_258), .B(n_251), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_259), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_267), .B(n_251), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_265), .B(n_236), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_259), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_265), .Y(n_296) );
INVx2_ASAP7_75t_SL g297 ( .A(n_276), .Y(n_297) );
BUFx3_ASAP7_75t_L g298 ( .A(n_280), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_263), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_274), .B(n_236), .Y(n_300) );
BUFx2_ASAP7_75t_L g301 ( .A(n_270), .Y(n_301) );
OAI21xp5_ASAP7_75t_L g302 ( .A1(n_262), .A2(n_239), .B(n_248), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_291), .B(n_248), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_291), .B(n_248), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_281), .Y(n_305) );
INVx5_ASAP7_75t_SL g306 ( .A(n_284), .Y(n_306) );
BUFx2_ASAP7_75t_L g307 ( .A(n_285), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_281), .Y(n_308) );
OAI21x1_ASAP7_75t_L g309 ( .A1(n_299), .A2(n_260), .B(n_233), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_292), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_282), .B(n_248), .Y(n_311) );
BUFx3_ASAP7_75t_L g312 ( .A(n_284), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_290), .B(n_243), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_282), .B(n_248), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_290), .B(n_248), .Y(n_315) );
INVx5_ASAP7_75t_L g316 ( .A(n_284), .Y(n_316) );
NAND3xp33_ASAP7_75t_L g317 ( .A(n_296), .B(n_275), .C(n_264), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_294), .B(n_243), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_292), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_283), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_283), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_286), .B(n_243), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_286), .B(n_243), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_287), .B(n_241), .Y(n_324) );
INVx2_ASAP7_75t_SL g325 ( .A(n_284), .Y(n_325) );
AO21x2_ASAP7_75t_L g326 ( .A1(n_302), .A2(n_270), .B(n_233), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_293), .B(n_243), .Y(n_327) );
AOI221xp5_ASAP7_75t_L g328 ( .A1(n_296), .A2(n_266), .B1(n_235), .B2(n_256), .C(n_238), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_288), .Y(n_329) );
AND2x4_ASAP7_75t_L g330 ( .A(n_287), .B(n_241), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_288), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_287), .B(n_241), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_316), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_325), .B(n_289), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_318), .B(n_289), .Y(n_335) );
OAI22xp5_ASAP7_75t_SL g336 ( .A1(n_316), .A2(n_298), .B1(n_242), .B2(n_273), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_325), .B(n_289), .Y(n_337) );
NAND3x1_ASAP7_75t_SL g338 ( .A(n_328), .B(n_302), .C(n_294), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_305), .B(n_293), .Y(n_339) );
NAND2x1_ASAP7_75t_L g340 ( .A(n_320), .B(n_297), .Y(n_340) );
OAI21x1_ASAP7_75t_L g341 ( .A1(n_309), .A2(n_299), .B(n_292), .Y(n_341) );
AND2x4_ASAP7_75t_L g342 ( .A(n_325), .B(n_297), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_312), .B(n_285), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_305), .B(n_298), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_318), .B(n_300), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_310), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_308), .B(n_298), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_318), .B(n_300), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_315), .B(n_301), .Y(n_349) );
OAI21xp5_ASAP7_75t_SL g350 ( .A1(n_328), .A2(n_268), .B(n_274), .Y(n_350) );
INVx2_ASAP7_75t_SL g351 ( .A(n_316), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_320), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_321), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_308), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_310), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_321), .Y(n_356) );
BUFx3_ASAP7_75t_L g357 ( .A(n_316), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_315), .B(n_301), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_329), .B(n_331), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_329), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_312), .B(n_297), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_315), .B(n_295), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_331), .B(n_235), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_310), .Y(n_364) );
OAI31xp33_ASAP7_75t_L g365 ( .A1(n_317), .A2(n_101), .A3(n_239), .B(n_247), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_303), .B(n_295), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_322), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_316), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_322), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_303), .B(n_295), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_304), .B(n_299), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_304), .B(n_243), .Y(n_372) );
INVx1_ASAP7_75t_SL g373 ( .A(n_316), .Y(n_373) );
INVxp67_ASAP7_75t_L g374 ( .A(n_311), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_312), .B(n_241), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_323), .Y(n_376) );
AND2x4_ASAP7_75t_L g377 ( .A(n_368), .B(n_316), .Y(n_377) );
AND2x2_ASAP7_75t_SL g378 ( .A(n_342), .B(n_307), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_376), .B(n_311), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_344), .B(n_317), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_376), .B(n_314), .Y(n_381) );
NOR2x1_ASAP7_75t_L g382 ( .A(n_368), .B(n_327), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_336), .A2(n_314), .B1(n_327), .B2(n_330), .Y(n_383) );
O2A1O1Ixp33_ASAP7_75t_L g384 ( .A1(n_365), .A2(n_323), .B(n_247), .C(n_101), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_352), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_374), .B(n_307), .Y(n_386) );
BUFx2_ASAP7_75t_L g387 ( .A(n_368), .Y(n_387) );
O2A1O1Ixp33_ASAP7_75t_L g388 ( .A1(n_350), .A2(n_347), .B(n_340), .C(n_351), .Y(n_388) );
AOI21xp5_ASAP7_75t_L g389 ( .A1(n_340), .A2(n_313), .B(n_326), .Y(n_389) );
OR2x6_ASAP7_75t_L g390 ( .A(n_351), .B(n_324), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_339), .B(n_313), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_352), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_353), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_367), .B(n_306), .Y(n_394) );
OAI21xp5_ASAP7_75t_L g395 ( .A1(n_375), .A2(n_309), .B(n_330), .Y(n_395) );
NOR3xp33_ASAP7_75t_L g396 ( .A(n_338), .B(n_277), .C(n_332), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_369), .B(n_345), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_346), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_353), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_335), .B(n_306), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_346), .Y(n_401) );
OAI22xp33_ASAP7_75t_L g402 ( .A1(n_361), .A2(n_332), .B1(n_330), .B2(n_324), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_356), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_349), .B(n_306), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_345), .B(n_324), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_348), .B(n_324), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_348), .B(n_330), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_354), .B(n_332), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_355), .Y(n_409) );
XNOR2x2_ASAP7_75t_L g410 ( .A(n_333), .B(n_309), .Y(n_410) );
OAI31xp33_ASAP7_75t_L g411 ( .A1(n_373), .A2(n_332), .A3(n_319), .B(n_253), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_360), .B(n_306), .Y(n_412) );
INVx1_ASAP7_75t_SL g413 ( .A(n_357), .Y(n_413) );
INVx1_ASAP7_75t_SL g414 ( .A(n_357), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_356), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_349), .B(n_306), .Y(n_416) );
OAI21xp33_ASAP7_75t_L g417 ( .A1(n_358), .A2(n_137), .B(n_319), .Y(n_417) );
INVx1_ASAP7_75t_SL g418 ( .A(n_371), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_358), .B(n_326), .Y(n_419) );
NAND2xp67_ASAP7_75t_L g420 ( .A(n_371), .B(n_319), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_359), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_361), .A2(n_253), .B1(n_252), .B2(n_137), .Y(n_422) );
INVx2_ASAP7_75t_SL g423 ( .A(n_343), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_335), .B(n_326), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_362), .B(n_326), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_372), .B(n_3), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_362), .B(n_4), .Y(n_427) );
INVx1_ASAP7_75t_SL g428 ( .A(n_343), .Y(n_428) );
OAI32xp33_ASAP7_75t_L g429 ( .A1(n_418), .A2(n_337), .A3(n_334), .B1(n_372), .B2(n_363), .Y(n_429) );
AOI221x1_ASAP7_75t_L g430 ( .A1(n_396), .A2(n_375), .B1(n_342), .B2(n_355), .C(n_364), .Y(n_430) );
OAI21xp5_ASAP7_75t_L g431 ( .A1(n_384), .A2(n_375), .B(n_342), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_380), .B(n_370), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_380), .B(n_370), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_421), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_396), .A2(n_366), .B1(n_334), .B2(n_337), .Y(n_435) );
OAI322xp33_ASAP7_75t_L g436 ( .A1(n_391), .A2(n_366), .A3(n_137), .B1(n_364), .B2(n_338), .C1(n_8), .C2(n_9), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_400), .B(n_341), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_385), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g439 ( .A1(n_417), .A2(n_341), .B(n_253), .Y(n_439) );
NAND2xp33_ASAP7_75t_R g440 ( .A(n_387), .B(n_377), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_391), .B(n_137), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_397), .B(n_137), .Y(n_442) );
AOI321xp33_ASAP7_75t_L g443 ( .A1(n_388), .A2(n_4), .A3(n_5), .B1(n_6), .B2(n_7), .C(n_9), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_383), .A2(n_241), .B1(n_133), .B2(n_252), .Y(n_444) );
NAND2xp33_ASAP7_75t_SL g445 ( .A(n_383), .B(n_5), .Y(n_445) );
INVx2_ASAP7_75t_SL g446 ( .A(n_423), .Y(n_446) );
AOI221xp5_ASAP7_75t_L g447 ( .A1(n_388), .A2(n_156), .B1(n_159), .B2(n_13), .C(n_14), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_382), .A2(n_250), .B1(n_231), .B2(n_232), .Y(n_448) );
OAI21xp33_ASAP7_75t_L g449 ( .A1(n_420), .A2(n_250), .B(n_231), .Y(n_449) );
AND2x4_ASAP7_75t_L g450 ( .A(n_377), .B(n_7), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_392), .Y(n_451) );
INVx4_ASAP7_75t_L g452 ( .A(n_390), .Y(n_452) );
AOI31xp33_ASAP7_75t_L g453 ( .A1(n_427), .A2(n_11), .A3(n_15), .B(n_16), .Y(n_453) );
AOI321xp33_ASAP7_75t_L g454 ( .A1(n_426), .A2(n_15), .A3(n_16), .B1(n_271), .B2(n_191), .C(n_196), .Y(n_454) );
A2O1A1Ixp33_ASAP7_75t_L g455 ( .A1(n_384), .A2(n_232), .B(n_231), .C(n_245), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_393), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_401), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_403), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_378), .A2(n_133), .B1(n_140), .B2(n_250), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_425), .B(n_232), .Y(n_460) );
OAI221xp5_ASAP7_75t_L g461 ( .A1(n_411), .A2(n_140), .B1(n_229), .B2(n_209), .C(n_226), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_378), .A2(n_140), .B1(n_244), .B2(n_245), .Y(n_462) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_389), .A2(n_244), .B(n_245), .Y(n_463) );
INVxp67_ASAP7_75t_L g464 ( .A(n_386), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_379), .B(n_140), .Y(n_465) );
AOI21xp33_ASAP7_75t_SL g466 ( .A1(n_402), .A2(n_390), .B(n_404), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_390), .A2(n_140), .B1(n_244), .B2(n_229), .Y(n_467) );
OAI21xp33_ASAP7_75t_L g468 ( .A1(n_419), .A2(n_140), .B(n_147), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_416), .A2(n_140), .B1(n_213), .B2(n_223), .Y(n_469) );
AOI222xp33_ASAP7_75t_L g470 ( .A1(n_424), .A2(n_147), .B1(n_255), .B2(n_213), .C1(n_223), .C2(n_197), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_381), .B(n_255), .Y(n_471) );
OAI22xp33_ASAP7_75t_L g472 ( .A1(n_413), .A2(n_223), .B1(n_213), .B2(n_147), .Y(n_472) );
NAND2x1_ASAP7_75t_SL g473 ( .A(n_401), .B(n_147), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_434), .Y(n_474) );
INVx1_ASAP7_75t_SL g475 ( .A(n_446), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_442), .Y(n_476) );
OAI222xp33_ASAP7_75t_L g477 ( .A1(n_452), .A2(n_414), .B1(n_428), .B2(n_402), .C1(n_394), .C2(n_405), .Y(n_477) );
OAI21xp33_ASAP7_75t_L g478 ( .A1(n_466), .A2(n_406), .B(n_407), .Y(n_478) );
OAI21xp5_ASAP7_75t_SL g479 ( .A1(n_453), .A2(n_395), .B(n_410), .Y(n_479) );
OAI221xp5_ASAP7_75t_L g480 ( .A1(n_443), .A2(n_412), .B1(n_408), .B2(n_415), .C(n_399), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_445), .A2(n_422), .B(n_409), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_457), .Y(n_482) );
AOI211xp5_ASAP7_75t_L g483 ( .A1(n_429), .A2(n_409), .B(n_398), .C(n_255), .Y(n_483) );
NAND2x1_ASAP7_75t_L g484 ( .A(n_452), .B(n_398), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_450), .B(n_223), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_437), .B(n_18), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_438), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_435), .A2(n_223), .B1(n_213), .B2(n_147), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g489 ( .A1(n_447), .A2(n_157), .B(n_21), .Y(n_489) );
INVx2_ASAP7_75t_SL g490 ( .A(n_473), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_451), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_432), .B(n_19), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_433), .B(n_23), .Y(n_493) );
NOR2x1_ASAP7_75t_L g494 ( .A(n_450), .B(n_223), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_456), .Y(n_495) );
XOR2x2_ASAP7_75t_L g496 ( .A(n_440), .B(n_24), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_441), .B(n_26), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_458), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_464), .B(n_27), .Y(n_499) );
OAI22xp33_ASAP7_75t_L g500 ( .A1(n_430), .A2(n_213), .B1(n_30), .B2(n_33), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_436), .B(n_28), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_465), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_460), .B(n_38), .Y(n_503) );
AOI21xp33_ASAP7_75t_L g504 ( .A1(n_479), .A2(n_501), .B(n_490), .Y(n_504) );
OAI211xp5_ASAP7_75t_SL g505 ( .A1(n_478), .A2(n_431), .B(n_454), .C(n_444), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_475), .A2(n_462), .B1(n_461), .B2(n_455), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_481), .A2(n_459), .B(n_468), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_483), .A2(n_471), .B1(n_467), .B2(n_448), .Y(n_508) );
AOI21xp33_ASAP7_75t_L g509 ( .A1(n_501), .A2(n_500), .B(n_492), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_500), .A2(n_439), .B(n_449), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_495), .Y(n_511) );
NAND5xp2_ASAP7_75t_L g512 ( .A(n_489), .B(n_470), .C(n_448), .D(n_469), .E(n_472), .Y(n_512) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_488), .B(n_463), .C(n_157), .Y(n_513) );
NOR3xp33_ASAP7_75t_L g514 ( .A(n_477), .B(n_463), .C(n_197), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_495), .Y(n_515) );
OAI21xp5_ASAP7_75t_SL g516 ( .A1(n_477), .A2(n_39), .B(n_42), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_496), .B(n_150), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_484), .A2(n_150), .B1(n_44), .B2(n_48), .Y(n_518) );
NOR2x1_ASAP7_75t_L g519 ( .A(n_494), .B(n_43), .Y(n_519) );
AOI221xp5_ASAP7_75t_L g520 ( .A1(n_480), .A2(n_189), .B1(n_179), .B2(n_171), .C(n_150), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_474), .B(n_49), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_504), .A2(n_485), .B(n_476), .C(n_486), .Y(n_522) );
OAI211xp5_ASAP7_75t_L g523 ( .A1(n_516), .A2(n_485), .B(n_499), .C(n_493), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_509), .A2(n_498), .B(n_491), .C(n_487), .Y(n_524) );
OAI221xp5_ASAP7_75t_L g525 ( .A1(n_505), .A2(n_502), .B1(n_482), .B2(n_503), .C(n_497), .Y(n_525) );
AOI221x1_ASAP7_75t_L g526 ( .A1(n_514), .A2(n_482), .B1(n_51), .B2(n_54), .C(n_55), .Y(n_526) );
AOI221xp5_ASAP7_75t_L g527 ( .A1(n_508), .A2(n_189), .B1(n_179), .B2(n_171), .C(n_58), .Y(n_527) );
BUFx2_ASAP7_75t_L g528 ( .A(n_519), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_520), .A2(n_189), .B1(n_179), .B2(n_171), .Y(n_529) );
AOI211xp5_ASAP7_75t_L g530 ( .A1(n_507), .A2(n_50), .B(n_56), .C(n_57), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_510), .A2(n_59), .B(n_65), .Y(n_531) );
NAND4xp75_ASAP7_75t_L g532 ( .A(n_531), .B(n_510), .C(n_517), .D(n_521), .Y(n_532) );
NOR3x1_ASAP7_75t_L g533 ( .A(n_525), .B(n_506), .C(n_513), .Y(n_533) );
OAI21xp5_ASAP7_75t_SL g534 ( .A1(n_522), .A2(n_518), .B(n_512), .Y(n_534) );
NAND4xp75_ASAP7_75t_L g535 ( .A(n_526), .B(n_511), .C(n_515), .D(n_70), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_524), .A2(n_66), .B(n_68), .Y(n_536) );
OR4x2_ASAP7_75t_L g537 ( .A(n_534), .B(n_528), .C(n_523), .D(n_530), .Y(n_537) );
AO22x2_ASAP7_75t_L g538 ( .A1(n_532), .A2(n_527), .B1(n_529), .B2(n_73), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_533), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_539), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_538), .Y(n_541) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_540), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_541), .A2(n_538), .B1(n_537), .B2(n_536), .Y(n_543) );
OAI22xp5_ASAP7_75t_SL g544 ( .A1(n_543), .A2(n_535), .B1(n_168), .B2(n_177), .Y(n_544) );
OAI21x1_ASAP7_75t_L g545 ( .A1(n_544), .A2(n_542), .B(n_168), .Y(n_545) );
OAI221xp5_ASAP7_75t_R g546 ( .A1(n_545), .A2(n_168), .B1(n_177), .B2(n_543), .C(n_539), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_546), .A2(n_168), .B1(n_177), .B2(n_539), .Y(n_547) );
endmodule