module real_aes_16114_n_344 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_344);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_344;
wire n_476;
wire n_887;
wire n_599;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1346;
wire n_1383;
wire n_552;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1250;
wire n_1284;
wire n_1095;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_346;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_1499;
wire n_399;
wire n_700;
wire n_948;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_1404;
wire n_733;
wire n_658;
wire n_1856;
wire n_676;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_1403;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_1840;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1175;
wire n_1170;
wire n_778;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1827;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_1802;
wire n_727;
wire n_397;
wire n_1056;
wire n_1855;
wire n_1083;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_1226;
wire n_1790;
wire n_525;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_1343;
wire n_719;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_1851;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_1826;
wire n_1836;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_1484;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI221xp5_ASAP7_75t_L g1081 ( .A1(n_0), .A2(n_103), .B1(n_465), .B2(n_1059), .C(n_1082), .Y(n_1081) );
AOI22xp33_ASAP7_75t_SL g1103 ( .A1(n_0), .A2(n_225), .B1(n_1104), .B2(n_1106), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g1577 ( .A1(n_1), .A2(n_86), .B1(n_1544), .B2(n_1549), .Y(n_1577) );
AOI22xp33_ASAP7_75t_L g1283 ( .A1(n_2), .A2(n_265), .B1(n_511), .B2(n_1008), .Y(n_1283) );
AOI22xp33_ASAP7_75t_L g1296 ( .A1(n_2), .A2(n_235), .B1(n_406), .B2(n_1297), .Y(n_1296) );
INVx1_ASAP7_75t_L g359 ( .A(n_3), .Y(n_359) );
AND2x2_ASAP7_75t_L g387 ( .A(n_3), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g400 ( .A(n_3), .B(n_242), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_3), .B(n_369), .Y(n_432) );
INVx1_ASAP7_75t_L g445 ( .A(n_4), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_4), .A2(n_78), .B1(n_473), .B2(n_485), .Y(n_472) );
INVx1_ASAP7_75t_L g947 ( .A(n_5), .Y(n_947) );
AOI22xp5_ASAP7_75t_L g968 ( .A1(n_5), .A2(n_12), .B1(n_969), .B2(n_970), .Y(n_968) );
OAI22xp5_ASAP7_75t_L g899 ( .A1(n_6), .A2(n_256), .B1(n_900), .B2(n_901), .Y(n_899) );
OAI22xp33_ASAP7_75t_L g913 ( .A1(n_6), .A2(n_256), .B1(n_914), .B2(n_916), .Y(n_913) );
INVx1_ASAP7_75t_L g997 ( .A(n_7), .Y(n_997) );
OAI221xp5_ASAP7_75t_L g1034 ( .A1(n_7), .A2(n_143), .B1(n_1035), .B2(n_1039), .C(n_1043), .Y(n_1034) );
INVx1_ASAP7_75t_L g1247 ( .A(n_8), .Y(n_1247) );
INVx1_ASAP7_75t_L g1071 ( .A(n_9), .Y(n_1071) );
OAI22xp33_ASAP7_75t_L g1112 ( .A1(n_9), .A2(n_92), .B1(n_1015), .B2(n_1113), .Y(n_1112) );
INVx1_ASAP7_75t_L g380 ( .A(n_10), .Y(n_380) );
INVx1_ASAP7_75t_L g1139 ( .A(n_11), .Y(n_1139) );
OA222x2_ASAP7_75t_L g1153 ( .A1(n_11), .A2(n_145), .B1(n_169), .B2(n_394), .C1(n_721), .C2(n_1154), .Y(n_1153) );
INVx1_ASAP7_75t_L g956 ( .A(n_12), .Y(n_956) );
INVxp67_ASAP7_75t_SL g1236 ( .A(n_13), .Y(n_1236) );
AOI22xp33_ASAP7_75t_L g1266 ( .A1(n_13), .A2(n_116), .B1(n_499), .B2(n_1129), .Y(n_1266) );
AOI22xp33_ASAP7_75t_L g1824 ( .A1(n_14), .A2(n_29), .B1(n_499), .B2(n_1825), .Y(n_1824) );
INVx1_ASAP7_75t_L g1857 ( .A(n_14), .Y(n_1857) );
INVx1_ASAP7_75t_L g1234 ( .A(n_15), .Y(n_1234) );
AOI22xp33_ASAP7_75t_L g1267 ( .A1(n_15), .A2(n_162), .B1(n_506), .B2(n_534), .Y(n_1267) );
AOI22xp33_ASAP7_75t_SL g1284 ( .A1(n_16), .A2(n_196), .B1(n_1002), .B2(n_1101), .Y(n_1284) );
AOI221xp5_ASAP7_75t_L g1295 ( .A1(n_16), .A2(n_113), .B1(n_570), .B2(n_1065), .C(n_1160), .Y(n_1295) );
INVx1_ASAP7_75t_L g895 ( .A(n_17), .Y(n_895) );
OAI221xp5_ASAP7_75t_L g1765 ( .A1(n_18), .A2(n_335), .B1(n_485), .B2(n_492), .C(n_1343), .Y(n_1765) );
OAI21xp33_ASAP7_75t_SL g1793 ( .A1(n_18), .A2(n_434), .B(n_721), .Y(n_1793) );
AOI22xp33_ASAP7_75t_L g1466 ( .A1(n_19), .A2(n_69), .B1(n_652), .B2(n_1130), .Y(n_1466) );
AOI221xp5_ASAP7_75t_L g1483 ( .A1(n_19), .A2(n_307), .B1(n_463), .B2(n_970), .C(n_1484), .Y(n_1483) );
AOI221xp5_ASAP7_75t_L g1058 ( .A1(n_20), .A2(n_91), .B1(n_1059), .B2(n_1061), .C(n_1064), .Y(n_1058) );
AOI22xp33_ASAP7_75t_SL g1111 ( .A1(n_20), .A2(n_187), .B1(n_499), .B2(n_1102), .Y(n_1111) );
INVx2_ASAP7_75t_L g482 ( .A(n_21), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_22), .A2(n_162), .B1(n_406), .B2(n_426), .Y(n_1244) );
AOI22xp5_ASAP7_75t_L g1268 ( .A1(n_22), .A2(n_305), .B1(n_506), .B2(n_524), .Y(n_1268) );
CKINVDCx5p33_ASAP7_75t_R g1378 ( .A(n_23), .Y(n_1378) );
INVx1_ASAP7_75t_L g850 ( .A(n_24), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g1131 ( .A1(n_25), .A2(n_172), .B1(n_1127), .B2(n_1132), .Y(n_1131) );
INVxp67_ASAP7_75t_SL g1168 ( .A(n_25), .Y(n_1168) );
OAI22xp33_ASAP7_75t_L g1776 ( .A1(n_26), .A2(n_280), .B1(n_1506), .B2(n_1507), .Y(n_1776) );
INVx1_ASAP7_75t_L g1792 ( .A(n_26), .Y(n_1792) );
OAI211xp5_ASAP7_75t_L g893 ( .A1(n_27), .A2(n_781), .B(n_817), .C(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g912 ( .A(n_27), .Y(n_912) );
CKINVDCx5p33_ASAP7_75t_R g1455 ( .A(n_28), .Y(n_1455) );
AOI221xp5_ASAP7_75t_L g1838 ( .A1(n_29), .A2(n_43), .B1(n_428), .B2(n_1297), .C(n_1839), .Y(n_1838) );
INVx1_ASAP7_75t_L g1328 ( .A(n_30), .Y(n_1328) );
AOI221xp5_ASAP7_75t_L g1345 ( .A1(n_30), .A2(n_141), .B1(n_652), .B2(n_1346), .C(n_1348), .Y(n_1345) );
INVx1_ASAP7_75t_L g690 ( .A(n_31), .Y(n_690) );
AOI221x1_ASAP7_75t_SL g697 ( .A1(n_31), .A2(n_185), .B1(n_406), .B2(n_588), .C(n_698), .Y(n_697) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_32), .Y(n_354) );
AND2x2_ASAP7_75t_L g1545 ( .A(n_32), .B(n_352), .Y(n_1545) );
OA22x2_ASAP7_75t_L g728 ( .A1(n_33), .A2(n_729), .B1(n_842), .B2(n_843), .Y(n_728) );
INVxp67_ASAP7_75t_L g843 ( .A(n_33), .Y(n_843) );
INVx1_ASAP7_75t_L g863 ( .A(n_34), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g1195 ( .A1(n_35), .A2(n_215), .B1(n_1110), .B2(n_1135), .Y(n_1195) );
AOI22xp5_ASAP7_75t_L g1216 ( .A1(n_35), .A2(n_289), .B1(n_428), .B2(n_575), .Y(n_1216) );
INVx1_ASAP7_75t_L g682 ( .A(n_36), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_36), .A2(n_173), .B1(n_423), .B2(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g770 ( .A(n_37), .Y(n_770) );
INVx1_ASAP7_75t_L g1404 ( .A(n_38), .Y(n_1404) );
OAI22xp5_ASAP7_75t_L g1447 ( .A1(n_38), .A2(n_63), .B1(n_718), .B2(n_1448), .Y(n_1447) );
AOI22xp33_ASAP7_75t_L g1826 ( .A1(n_39), .A2(n_195), .B1(n_1417), .B2(n_1468), .Y(n_1826) );
INVx1_ASAP7_75t_L g1842 ( .A(n_39), .Y(n_1842) );
INVx1_ASAP7_75t_L g1336 ( .A(n_40), .Y(n_1336) );
OAI22xp33_ASAP7_75t_L g1342 ( .A1(n_40), .A2(n_51), .B1(n_485), .B2(n_1343), .Y(n_1342) );
AOI22xp33_ASAP7_75t_L g1576 ( .A1(n_41), .A2(n_68), .B1(n_1552), .B2(n_1561), .Y(n_1576) );
AOI22xp33_ASAP7_75t_L g1282 ( .A1(n_42), .A2(n_235), .B1(n_511), .B2(n_1008), .Y(n_1282) );
AOI221xp5_ASAP7_75t_L g1292 ( .A1(n_42), .A2(n_265), .B1(n_590), .B2(n_1060), .C(n_1063), .Y(n_1292) );
AOI22xp33_ASAP7_75t_SL g1828 ( .A1(n_43), .A2(n_308), .B1(n_499), .B2(n_1829), .Y(n_1828) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_44), .A2(n_555), .B1(n_556), .B2(n_557), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_44), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g678 ( .A(n_45), .Y(n_678) );
AOI22xp33_ASAP7_75t_SL g1126 ( .A1(n_46), .A2(n_263), .B1(n_1099), .B2(n_1127), .Y(n_1126) );
INVxp67_ASAP7_75t_SL g1162 ( .A(n_46), .Y(n_1162) );
INVxp67_ASAP7_75t_SL g1238 ( .A(n_47), .Y(n_1238) );
AOI22xp33_ASAP7_75t_SL g1269 ( .A1(n_47), .A2(n_88), .B1(n_499), .B2(n_1129), .Y(n_1269) );
OAI22xp5_ASAP7_75t_L g1366 ( .A1(n_48), .A2(n_932), .B1(n_1367), .B2(n_1370), .Y(n_1366) );
INVx1_ASAP7_75t_L g1384 ( .A(n_48), .Y(n_1384) );
CKINVDCx5p33_ASAP7_75t_R g1276 ( .A(n_49), .Y(n_1276) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_50), .A2(n_181), .B1(n_406), .B2(n_427), .Y(n_592) );
INVx1_ASAP7_75t_L g643 ( .A(n_50), .Y(n_643) );
OAI221xp5_ASAP7_75t_L g1332 ( .A1(n_51), .A2(n_300), .B1(n_434), .B2(n_716), .C(n_718), .Y(n_1332) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_52), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g1827 ( .A1(n_53), .A2(n_65), .B1(n_652), .B2(n_1132), .Y(n_1827) );
INVx1_ASAP7_75t_L g1841 ( .A(n_53), .Y(n_1841) );
AOI221xp5_ASAP7_75t_L g1420 ( .A1(n_54), .A2(n_321), .B1(n_509), .B2(n_519), .C(n_1421), .Y(n_1420) );
AOI22xp33_ASAP7_75t_L g1427 ( .A1(n_54), .A2(n_167), .B1(n_463), .B2(n_1061), .Y(n_1427) );
INVx1_ASAP7_75t_L g1286 ( .A(n_55), .Y(n_1286) );
INVx1_ASAP7_75t_L g946 ( .A(n_56), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_56), .A2(n_176), .B1(n_422), .B2(n_969), .Y(n_974) );
OAI22xp5_ASAP7_75t_L g1401 ( .A1(n_57), .A2(n_186), .B1(n_930), .B2(n_932), .Y(n_1401) );
CKINVDCx5p33_ASAP7_75t_R g1432 ( .A(n_57), .Y(n_1432) );
CKINVDCx5p33_ASAP7_75t_R g1819 ( .A(n_58), .Y(n_1819) );
AOI22xp5_ASAP7_75t_L g1560 ( .A1(n_59), .A2(n_107), .B1(n_1552), .B2(n_1561), .Y(n_1560) );
CKINVDCx5p33_ASAP7_75t_R g1323 ( .A(n_60), .Y(n_1323) );
AOI22xp5_ASAP7_75t_L g1568 ( .A1(n_61), .A2(n_245), .B1(n_1552), .B2(n_1561), .Y(n_1568) );
INVx1_ASAP7_75t_L g1372 ( .A(n_62), .Y(n_1372) );
AOI22xp33_ASAP7_75t_L g1392 ( .A1(n_62), .A2(n_66), .B1(n_427), .B2(n_456), .Y(n_1392) );
INVx1_ASAP7_75t_L g1424 ( .A(n_63), .Y(n_1424) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_64), .A2(n_207), .B1(n_426), .B2(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g637 ( .A(n_64), .Y(n_637) );
INVx1_ASAP7_75t_L g1861 ( .A(n_65), .Y(n_1861) );
AOI221xp5_ASAP7_75t_L g1361 ( .A1(n_66), .A2(n_328), .B1(n_506), .B2(n_1136), .C(n_1362), .Y(n_1361) );
INVxp67_ASAP7_75t_SL g1334 ( .A(n_67), .Y(n_1334) );
OAI22xp5_ASAP7_75t_L g1349 ( .A1(n_67), .A2(n_932), .B1(n_1350), .B2(n_1351), .Y(n_1349) );
AOI22xp33_ASAP7_75t_SL g1481 ( .A1(n_69), .A2(n_144), .B1(n_568), .B2(n_976), .Y(n_1481) );
AOI21xp33_ASAP7_75t_L g1777 ( .A1(n_70), .A2(n_1778), .B(n_1781), .Y(n_1777) );
AOI221xp5_ASAP7_75t_L g1802 ( .A1(n_70), .A2(n_104), .B1(n_1059), .B2(n_1803), .C(n_1804), .Y(n_1802) );
INVx1_ASAP7_75t_L g1177 ( .A(n_71), .Y(n_1177) );
INVx1_ASAP7_75t_L g1405 ( .A(n_72), .Y(n_1405) );
OAI21xp33_ASAP7_75t_L g1446 ( .A1(n_72), .A2(n_434), .B(n_721), .Y(n_1446) );
OAI22xp5_ASAP7_75t_L g1848 ( .A1(n_73), .A2(n_293), .B1(n_700), .B2(n_710), .Y(n_1848) );
INVx1_ASAP7_75t_L g1863 ( .A(n_73), .Y(n_1863) );
CKINVDCx5p33_ASAP7_75t_R g1186 ( .A(n_74), .Y(n_1186) );
AOI22xp33_ASAP7_75t_L g1583 ( .A1(n_75), .A2(n_230), .B1(n_1552), .B2(n_1561), .Y(n_1583) );
INVx1_ASAP7_75t_L g1338 ( .A(n_76), .Y(n_1338) );
OAI222xp33_ASAP7_75t_L g1341 ( .A1(n_76), .A2(n_286), .B1(n_300), .B2(n_609), .C1(n_675), .C2(n_812), .Y(n_1341) );
AOI22xp5_ASAP7_75t_L g1543 ( .A1(n_77), .A2(n_240), .B1(n_1544), .B2(n_1549), .Y(n_1543) );
INVx1_ASAP7_75t_L g410 ( .A(n_78), .Y(n_410) );
OAI22xp33_ASAP7_75t_L g759 ( .A1(n_79), .A2(n_177), .B1(n_760), .B2(n_762), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g828 ( .A1(n_79), .A2(n_177), .B1(n_829), .B2(n_833), .Y(n_828) );
AOI22xp5_ASAP7_75t_L g1551 ( .A1(n_80), .A2(n_99), .B1(n_1552), .B2(n_1554), .Y(n_1551) );
AO22x1_ASAP7_75t_L g1574 ( .A1(n_81), .A2(n_246), .B1(n_1544), .B2(n_1549), .Y(n_1574) );
OAI221xp5_ASAP7_75t_L g560 ( .A1(n_82), .A2(n_122), .B1(n_561), .B2(n_563), .C(n_567), .Y(n_560) );
INVx1_ASAP7_75t_L g606 ( .A(n_82), .Y(n_606) );
CKINVDCx5p33_ASAP7_75t_R g1410 ( .A(n_83), .Y(n_1410) );
AOI22xp33_ASAP7_75t_SL g1011 ( .A1(n_84), .A2(n_340), .B1(n_499), .B2(n_1002), .Y(n_1011) );
AOI221xp5_ASAP7_75t_L g1023 ( .A1(n_84), .A2(n_191), .B1(n_588), .B2(n_589), .C(n_1024), .Y(n_1023) );
CKINVDCx5p33_ASAP7_75t_R g1254 ( .A(n_85), .Y(n_1254) );
XOR2xp5_ASAP7_75t_L g1272 ( .A(n_86), .B(n_1273), .Y(n_1272) );
INVx1_ASAP7_75t_L g793 ( .A(n_87), .Y(n_793) );
AOI221xp5_ASAP7_75t_L g1241 ( .A1(n_88), .A2(n_116), .B1(n_594), .B2(n_969), .C(n_1242), .Y(n_1241) );
OAI22xp5_ASAP7_75t_L g1086 ( .A1(n_89), .A2(n_192), .B1(n_1087), .B2(n_1088), .Y(n_1086) );
INVx1_ASAP7_75t_L g571 ( .A(n_90), .Y(n_571) );
OAI221xp5_ASAP7_75t_SL g619 ( .A1(n_90), .A2(n_119), .B1(n_488), .B2(n_620), .C(n_621), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_91), .A2(n_264), .B1(n_1098), .B2(n_1102), .Y(n_1097) );
INVx1_ASAP7_75t_L g1069 ( .A(n_92), .Y(n_1069) );
AOI221xp5_ASAP7_75t_L g1508 ( .A1(n_93), .A2(n_316), .B1(n_652), .B2(n_1414), .C(n_1509), .Y(n_1508) );
INVx1_ASAP7_75t_L g1533 ( .A(n_93), .Y(n_1533) );
OAI22xp5_ASAP7_75t_L g1766 ( .A1(n_94), .A2(n_200), .B1(n_930), .B2(n_932), .Y(n_1766) );
INVxp67_ASAP7_75t_SL g1801 ( .A(n_94), .Y(n_1801) );
INVx1_ASAP7_75t_L g1300 ( .A(n_95), .Y(n_1300) );
AOI221xp5_ASAP7_75t_L g1134 ( .A1(n_96), .A2(n_112), .B1(n_509), .B2(n_519), .C(n_1135), .Y(n_1134) );
AOI22xp33_ASAP7_75t_SL g1169 ( .A1(n_96), .A2(n_263), .B1(n_427), .B2(n_428), .Y(n_1169) );
AOI222xp33_ASAP7_75t_L g1782 ( .A1(n_97), .A2(n_149), .B1(n_325), .B2(n_507), .C1(n_526), .C2(n_681), .Y(n_1782) );
INVx1_ASAP7_75t_L g1805 ( .A(n_97), .Y(n_1805) );
CKINVDCx5p33_ASAP7_75t_R g1324 ( .A(n_98), .Y(n_1324) );
AOI22xp33_ASAP7_75t_L g1810 ( .A1(n_99), .A2(n_1811), .B1(n_1814), .B2(n_1866), .Y(n_1810) );
INVx1_ASAP7_75t_L g1865 ( .A(n_99), .Y(n_1865) );
OAI22xp33_ASAP7_75t_L g1379 ( .A1(n_100), .A2(n_146), .B1(n_485), .B2(n_1343), .Y(n_1379) );
OAI22xp5_ASAP7_75t_L g1393 ( .A1(n_100), .A2(n_284), .B1(n_716), .B2(n_718), .Y(n_1393) );
INVx1_ASAP7_75t_L g796 ( .A(n_101), .Y(n_796) );
CKINVDCx5p33_ASAP7_75t_R g1329 ( .A(n_102), .Y(n_1329) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_103), .A2(n_267), .B1(n_1108), .B2(n_1110), .Y(n_1107) );
AOI221xp5_ASAP7_75t_L g1768 ( .A1(n_104), .A2(n_214), .B1(n_1769), .B2(n_1771), .C(n_1773), .Y(n_1768) );
INVx1_ASAP7_75t_L g352 ( .A(n_105), .Y(n_352) );
INVx1_ASAP7_75t_L g1369 ( .A(n_106), .Y(n_1369) );
AOI22xp33_ASAP7_75t_L g1389 ( .A1(n_106), .A2(n_328), .B1(n_406), .B2(n_427), .Y(n_1389) );
INVx1_ASAP7_75t_L g1335 ( .A(n_108), .Y(n_1335) );
AO221x2_ASAP7_75t_L g1661 ( .A1(n_109), .A2(n_324), .B1(n_1544), .B2(n_1549), .C(n_1662), .Y(n_1661) );
AOI221xp5_ASAP7_75t_L g593 ( .A1(n_110), .A2(n_150), .B1(n_588), .B2(n_589), .C(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g630 ( .A(n_110), .Y(n_630) );
INVx1_ASAP7_75t_L g1764 ( .A(n_111), .Y(n_1764) );
OAI21xp33_ASAP7_75t_L g1789 ( .A1(n_111), .A2(n_720), .B(n_1790), .Y(n_1789) );
AOI221xp5_ASAP7_75t_L g1159 ( .A1(n_112), .A2(n_155), .B1(n_589), .B2(n_1160), .C(n_1161), .Y(n_1159) );
AOI22xp33_ASAP7_75t_L g1279 ( .A1(n_113), .A2(n_241), .B1(n_1280), .B2(n_1281), .Y(n_1279) );
INVx1_ASAP7_75t_L g855 ( .A(n_114), .Y(n_855) );
INVx1_ASAP7_75t_L g954 ( .A(n_115), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_115), .A2(n_159), .B1(n_406), .B2(n_427), .Y(n_971) );
XOR2x2_ASAP7_75t_L g1490 ( .A(n_117), .B(n_1491), .Y(n_1490) );
CKINVDCx5p33_ASAP7_75t_R g1835 ( .A(n_118), .Y(n_1835) );
INVx1_ASAP7_75t_L g583 ( .A(n_119), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g943 ( .A(n_120), .Y(n_943) );
INVx1_ASAP7_75t_L g656 ( .A(n_121), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_121), .A2(n_238), .B1(n_716), .B2(n_718), .Y(n_715) );
INVx1_ASAP7_75t_L g600 ( .A(n_122), .Y(n_600) );
INVx1_ASAP7_75t_L g1504 ( .A(n_123), .Y(n_1504) );
INVx1_ASAP7_75t_L g1511 ( .A(n_124), .Y(n_1511) );
XOR2x2_ASAP7_75t_L g982 ( .A(n_125), .B(n_983), .Y(n_982) );
OAI221xp5_ASAP7_75t_L g929 ( .A1(n_126), .A2(n_277), .B1(n_930), .B2(n_932), .C(n_934), .Y(n_929) );
INVx1_ASAP7_75t_L g980 ( .A(n_126), .Y(n_980) );
AOI22xp5_ASAP7_75t_L g1173 ( .A1(n_127), .A2(n_1174), .B1(n_1175), .B2(n_1222), .Y(n_1173) );
INVx1_ASAP7_75t_L g1222 ( .A(n_127), .Y(n_1222) );
INVx1_ASAP7_75t_L g1510 ( .A(n_128), .Y(n_1510) );
INVx1_ASAP7_75t_L g577 ( .A(n_129), .Y(n_577) );
OAI21xp33_ASAP7_75t_L g615 ( .A1(n_129), .A2(n_616), .B(n_618), .Y(n_615) );
CKINVDCx5p33_ASAP7_75t_R g1456 ( .A(n_130), .Y(n_1456) );
CKINVDCx5p33_ASAP7_75t_R g1364 ( .A(n_131), .Y(n_1364) );
OAI22xp5_ASAP7_75t_L g1505 ( .A1(n_132), .A2(n_189), .B1(n_1506), .B2(n_1507), .Y(n_1505) );
OAI22xp5_ASAP7_75t_L g1520 ( .A1(n_132), .A2(n_273), .B1(n_441), .B2(n_447), .Y(n_1520) );
AOI22xp33_ASAP7_75t_SL g425 ( .A1(n_133), .A2(n_247), .B1(n_426), .B2(n_428), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g518 ( .A1(n_133), .A2(n_323), .B1(n_499), .B2(n_509), .C(n_519), .Y(n_518) );
OAI22xp33_ASAP7_75t_L g903 ( .A1(n_134), .A2(n_311), .B1(n_904), .B2(n_905), .Y(n_903) );
OAI22xp5_ASAP7_75t_L g907 ( .A1(n_134), .A2(n_311), .B1(n_740), .B2(n_908), .Y(n_907) );
CKINVDCx5p33_ASAP7_75t_R g987 ( .A(n_135), .Y(n_987) );
OAI211xp5_ASAP7_75t_SL g1239 ( .A1(n_136), .A2(n_1056), .B(n_1240), .C(n_1245), .Y(n_1239) );
INVx1_ASAP7_75t_L g1263 ( .A(n_136), .Y(n_1263) );
AOI22xp33_ASAP7_75t_SL g1462 ( .A1(n_137), .A2(n_294), .B1(n_1463), .B2(n_1465), .Y(n_1462) );
AOI22xp33_ASAP7_75t_L g1485 ( .A1(n_137), .A2(n_282), .B1(n_568), .B2(n_976), .Y(n_1485) );
OAI22xp5_ASAP7_75t_L g1496 ( .A1(n_138), .A2(n_211), .B1(n_930), .B2(n_932), .Y(n_1496) );
INVxp67_ASAP7_75t_SL g1518 ( .A(n_138), .Y(n_1518) );
AO22x1_ASAP7_75t_L g1565 ( .A1(n_139), .A2(n_329), .B1(n_1544), .B2(n_1549), .Y(n_1565) );
OAI222xp33_ASAP7_75t_L g1229 ( .A1(n_140), .A2(n_258), .B1(n_1040), .B2(n_1230), .C1(n_1231), .C2(n_1235), .Y(n_1229) );
INVx1_ASAP7_75t_L g1257 ( .A(n_140), .Y(n_1257) );
INVx1_ASAP7_75t_L g1312 ( .A(n_141), .Y(n_1312) );
XNOR2x1_ASAP7_75t_L g1225 ( .A(n_142), .B(n_1226), .Y(n_1225) );
INVx1_ASAP7_75t_L g995 ( .A(n_143), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g1467 ( .A1(n_144), .A2(n_307), .B1(n_526), .B2(n_1468), .Y(n_1467) );
INVx1_ASAP7_75t_L g1149 ( .A(n_145), .Y(n_1149) );
INVx1_ASAP7_75t_L g1385 ( .A(n_146), .Y(n_1385) );
AOI221xp5_ASAP7_75t_SL g587 ( .A1(n_147), .A2(n_304), .B1(n_588), .B2(n_589), .C(n_590), .Y(n_587) );
INVx1_ASAP7_75t_L g640 ( .A(n_147), .Y(n_640) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_148), .Y(n_585) );
INVx1_ASAP7_75t_L g1799 ( .A(n_149), .Y(n_1799) );
INVx1_ASAP7_75t_L g644 ( .A(n_150), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_151), .A2(n_298), .B1(n_511), .B2(n_1005), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_151), .A2(n_253), .B1(n_1026), .B2(n_1027), .Y(n_1025) );
INVx1_ASAP7_75t_L g1411 ( .A(n_152), .Y(n_1411) );
AOI22xp33_ASAP7_75t_SL g1428 ( .A1(n_152), .A2(n_163), .B1(n_1429), .B2(n_1430), .Y(n_1428) );
INVx1_ASAP7_75t_L g938 ( .A(n_153), .Y(n_938) );
OAI22xp5_ASAP7_75t_L g966 ( .A1(n_153), .A2(n_318), .B1(n_441), .B2(n_447), .Y(n_966) );
CKINVDCx5p33_ASAP7_75t_R g669 ( .A(n_154), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g1128 ( .A1(n_155), .A2(n_178), .B1(n_516), .B2(n_1129), .C(n_1130), .Y(n_1128) );
AO22x1_ASAP7_75t_L g1572 ( .A1(n_156), .A2(n_330), .B1(n_1552), .B2(n_1573), .Y(n_1572) );
CKINVDCx16_ASAP7_75t_R g1663 ( .A(n_157), .Y(n_1663) );
INVxp67_ASAP7_75t_SL g1181 ( .A(n_158), .Y(n_1181) );
OAI221xp5_ASAP7_75t_L g1196 ( .A1(n_158), .A2(n_492), .B1(n_930), .B2(n_1197), .C(n_1202), .Y(n_1196) );
INVx1_ASAP7_75t_L g949 ( .A(n_159), .Y(n_949) );
AOI21xp5_ASAP7_75t_L g1194 ( .A1(n_160), .A2(n_516), .B(n_1108), .Y(n_1194) );
INVx1_ASAP7_75t_L g1211 ( .A(n_160), .Y(n_1211) );
INVx1_ASAP7_75t_L g1201 ( .A(n_161), .Y(n_1201) );
AOI22xp33_ASAP7_75t_SL g1213 ( .A1(n_161), .A2(n_215), .B1(n_596), .B2(n_1026), .Y(n_1213) );
INVx1_ASAP7_75t_L g1419 ( .A(n_163), .Y(n_1419) );
INVx1_ASAP7_75t_L g1275 ( .A(n_164), .Y(n_1275) );
OAI221xp5_ASAP7_75t_L g1495 ( .A1(n_165), .A2(n_273), .B1(n_485), .B2(n_492), .C(n_1343), .Y(n_1495) );
INVxp67_ASAP7_75t_SL g1516 ( .A(n_165), .Y(n_1516) );
INVx1_ASAP7_75t_L g1374 ( .A(n_166), .Y(n_1374) );
AOI221xp5_ASAP7_75t_L g1412 ( .A1(n_167), .A2(n_297), .B1(n_516), .B2(n_1413), .C(n_1414), .Y(n_1412) );
INVx1_ASAP7_75t_L g896 ( .A(n_168), .Y(n_896) );
OAI211xp5_ASAP7_75t_L g909 ( .A1(n_168), .A2(n_747), .B(n_869), .C(n_910), .Y(n_909) );
OAI221xp5_ASAP7_75t_L g1143 ( .A1(n_169), .A2(n_171), .B1(n_683), .B2(n_1144), .C(n_1145), .Y(n_1143) );
INVx1_ASAP7_75t_L g1246 ( .A(n_170), .Y(n_1246) );
INVxp67_ASAP7_75t_SL g1156 ( .A(n_171), .Y(n_1156) );
INVxp33_ASAP7_75t_SL g1163 ( .A(n_172), .Y(n_1163) );
INVx1_ASAP7_75t_L g672 ( .A(n_173), .Y(n_672) );
INVx2_ASAP7_75t_L g1547 ( .A(n_174), .Y(n_1547) );
AND2x2_ASAP7_75t_L g1550 ( .A(n_174), .B(n_1548), .Y(n_1550) );
AND2x2_ASAP7_75t_L g1555 ( .A(n_174), .B(n_291), .Y(n_1555) );
INVx1_ASAP7_75t_L g1287 ( .A(n_175), .Y(n_1287) );
INVx1_ASAP7_75t_L g953 ( .A(n_176), .Y(n_953) );
INVx1_ASAP7_75t_L g1166 ( .A(n_178), .Y(n_1166) );
INVx1_ASAP7_75t_L g981 ( .A(n_179), .Y(n_981) );
OAI21xp33_ASAP7_75t_L g393 ( .A1(n_180), .A2(n_394), .B(n_401), .Y(n_393) );
OAI221xp5_ASAP7_75t_L g532 ( .A1(n_180), .A2(n_275), .B1(n_533), .B2(n_535), .C(n_539), .Y(n_532) );
INVx1_ASAP7_75t_L g629 ( .A(n_181), .Y(n_629) );
OAI21xp5_ASAP7_75t_SL g1399 ( .A1(n_182), .A2(n_927), .B(n_1400), .Y(n_1399) );
INVx1_ASAP7_75t_L g1423 ( .A(n_182), .Y(n_1423) );
INVx1_ASAP7_75t_L g853 ( .A(n_183), .Y(n_853) );
CKINVDCx5p33_ASAP7_75t_R g666 ( .A(n_184), .Y(n_666) );
INVx1_ASAP7_75t_L g676 ( .A(n_185), .Y(n_676) );
INVx1_ASAP7_75t_L g1440 ( .A(n_186), .Y(n_1440) );
INVxp67_ASAP7_75t_SL g1080 ( .A(n_187), .Y(n_1080) );
CKINVDCx5p33_ASAP7_75t_R g1460 ( .A(n_188), .Y(n_1460) );
OAI211xp5_ASAP7_75t_L g1513 ( .A1(n_189), .A2(n_927), .B(n_1514), .C(n_1517), .Y(n_1513) );
INVx1_ASAP7_75t_L g1148 ( .A(n_190), .Y(n_1148) );
OAI22xp5_ASAP7_75t_L g1170 ( .A1(n_190), .A2(n_227), .B1(n_441), .B2(n_447), .Y(n_1170) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_191), .A2(n_201), .B1(n_499), .B2(n_1002), .Y(n_1001) );
OAI211xp5_ASAP7_75t_L g1055 ( .A1(n_192), .A2(n_1056), .B(n_1057), .C(n_1068), .Y(n_1055) );
CKINVDCx5p33_ASAP7_75t_R g1204 ( .A(n_193), .Y(n_1204) );
AOI22xp33_ASAP7_75t_SL g417 ( .A1(n_194), .A2(n_313), .B1(n_418), .B2(n_422), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g508 ( .A1(n_194), .A2(n_222), .B1(n_509), .B2(n_511), .C(n_516), .Y(n_508) );
INVx1_ASAP7_75t_L g1859 ( .A(n_195), .Y(n_1859) );
AOI22xp33_ASAP7_75t_L g1293 ( .A1(n_196), .A2(n_241), .B1(n_426), .B2(n_428), .Y(n_1293) );
AOI22xp33_ASAP7_75t_SL g1469 ( .A1(n_197), .A2(n_282), .B1(n_602), .B2(n_1465), .Y(n_1469) );
AOI221xp5_ASAP7_75t_L g1477 ( .A1(n_197), .A2(n_294), .B1(n_1059), .B2(n_1065), .C(n_1478), .Y(n_1477) );
INVx2_ASAP7_75t_L g484 ( .A(n_198), .Y(n_484) );
INVx1_ASAP7_75t_L g522 ( .A(n_198), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_198), .B(n_482), .Y(n_531) );
OAI211xp5_ASAP7_75t_L g1402 ( .A1(n_199), .A2(n_492), .B(n_543), .C(n_1403), .Y(n_1402) );
CKINVDCx5p33_ASAP7_75t_R g1445 ( .A(n_199), .Y(n_1445) );
INVxp67_ASAP7_75t_SL g1785 ( .A(n_200), .Y(n_1785) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_201), .A2(n_340), .B1(n_426), .B2(n_1027), .Y(n_1046) );
XOR2xp5_ASAP7_75t_L g646 ( .A(n_202), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g1305 ( .A(n_203), .Y(n_1305) );
OAI221xp5_ASAP7_75t_SL g1074 ( .A1(n_204), .A2(n_292), .B1(n_1039), .B2(n_1075), .C(n_1076), .Y(n_1074) );
INVx1_ASAP7_75t_L g1092 ( .A(n_204), .Y(n_1092) );
INVx1_ASAP7_75t_L g957 ( .A(n_205), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_205), .A2(n_314), .B1(n_568), .B2(n_976), .Y(n_975) );
OAI22xp33_ASAP7_75t_L g657 ( .A1(n_206), .A2(n_303), .B1(n_658), .B2(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g724 ( .A(n_206), .Y(n_724) );
INVx1_ASAP7_75t_L g641 ( .A(n_207), .Y(n_641) );
INVx1_ASAP7_75t_L g780 ( .A(n_208), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g1473 ( .A(n_209), .Y(n_1473) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_210), .A2(n_322), .B1(n_426), .B2(n_454), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_210), .A2(n_247), .B1(n_499), .B2(n_506), .Y(n_498) );
INVxp67_ASAP7_75t_SL g1515 ( .A(n_211), .Y(n_1515) );
OAI22xp5_ASAP7_75t_L g988 ( .A1(n_212), .A2(n_296), .B1(n_989), .B2(n_990), .Y(n_988) );
OAI211xp5_ASAP7_75t_L g1019 ( .A1(n_212), .A2(n_1020), .B(n_1022), .C(n_1029), .Y(n_1019) );
BUFx3_ASAP7_75t_L g490 ( .A(n_213), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g1795 ( .A(n_214), .B(n_1796), .Y(n_1795) );
OAI21xp5_ASAP7_75t_SL g1488 ( .A1(n_216), .A2(n_1087), .B(n_1489), .Y(n_1488) );
AOI22xp33_ASAP7_75t_L g1584 ( .A1(n_217), .A2(n_224), .B1(n_1544), .B2(n_1549), .Y(n_1584) );
INVx1_ASAP7_75t_L g1774 ( .A(n_218), .Y(n_1774) );
INVx1_ASAP7_75t_L g402 ( .A(n_219), .Y(n_402) );
OAI221xp5_ASAP7_75t_L g1375 ( .A1(n_220), .A2(n_284), .B1(n_1193), .B2(n_1376), .C(n_1377), .Y(n_1375) );
OAI211xp5_ASAP7_75t_L g1382 ( .A1(n_220), .A2(n_547), .B(n_1383), .C(n_1386), .Y(n_1382) );
CKINVDCx5p33_ASAP7_75t_R g1363 ( .A(n_221), .Y(n_1363) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_222), .A2(n_323), .B1(n_463), .B2(n_465), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g1249 ( .A1(n_223), .A2(n_989), .B(n_1250), .Y(n_1249) );
XOR2xp5_ASAP7_75t_L g1052 ( .A(n_224), .B(n_1053), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_225), .A2(n_267), .B1(n_454), .B2(n_1067), .Y(n_1066) );
OAI22xp33_ASAP7_75t_L g1012 ( .A1(n_226), .A2(n_334), .B1(n_1013), .B2(n_1015), .Y(n_1012) );
INVx1_ASAP7_75t_L g1030 ( .A(n_226), .Y(n_1030) );
INVx1_ASAP7_75t_L g1138 ( .A(n_227), .Y(n_1138) );
OAI211xp5_ASAP7_75t_SL g744 ( .A1(n_228), .A2(n_745), .B(n_747), .C(n_749), .Y(n_744) );
INVx1_ASAP7_75t_L g824 ( .A(n_228), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g1085 ( .A(n_229), .Y(n_1085) );
CKINVDCx5p33_ASAP7_75t_R g1180 ( .A(n_231), .Y(n_1180) );
INVx1_ASAP7_75t_L g1502 ( .A(n_232), .Y(n_1502) );
INVx1_ASAP7_75t_L g758 ( .A(n_233), .Y(n_758) );
OAI211xp5_ASAP7_75t_SL g815 ( .A1(n_233), .A2(n_816), .B(n_817), .C(n_820), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g1319 ( .A(n_234), .Y(n_1319) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_236), .A2(n_253), .B1(n_511), .B2(n_1008), .Y(n_1007) );
INVx1_ASAP7_75t_L g1044 ( .A(n_236), .Y(n_1044) );
OAI211xp5_ASAP7_75t_L g940 ( .A1(n_237), .A2(n_492), .B(n_545), .C(n_941), .Y(n_940) );
INVxp33_ASAP7_75t_SL g965 ( .A(n_237), .Y(n_965) );
OAI221xp5_ASAP7_75t_L g662 ( .A1(n_238), .A2(n_255), .B1(n_488), .B2(n_620), .C(n_631), .Y(n_662) );
INVx1_ASAP7_75t_L g1494 ( .A(n_239), .Y(n_1494) );
BUFx3_ASAP7_75t_L g369 ( .A(n_242), .Y(n_369) );
INVx1_ASAP7_75t_L g388 ( .A(n_242), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g1665 ( .A(n_243), .Y(n_1665) );
AOI22xp5_ASAP7_75t_L g1567 ( .A1(n_244), .A2(n_259), .B1(n_1544), .B2(n_1549), .Y(n_1567) );
NOR2xp33_ASAP7_75t_L g1218 ( .A(n_248), .B(n_1219), .Y(n_1218) );
CKINVDCx5p33_ASAP7_75t_R g686 ( .A(n_249), .Y(n_686) );
INVxp67_ASAP7_75t_SL g376 ( .A(n_250), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_251), .Y(n_569) );
INVx1_ASAP7_75t_L g1188 ( .A(n_252), .Y(n_1188) );
CKINVDCx5p33_ASAP7_75t_R g1371 ( .A(n_254), .Y(n_1371) );
OA222x2_ASAP7_75t_L g719 ( .A1(n_255), .A2(n_272), .B1(n_326), .B2(n_394), .C1(n_720), .C2(n_721), .Y(n_719) );
INVx1_ASAP7_75t_L g868 ( .A(n_257), .Y(n_868) );
INVx1_ASAP7_75t_L g1260 ( .A(n_258), .Y(n_1260) );
OAI21xp5_ASAP7_75t_L g1301 ( .A1(n_260), .A2(n_1087), .B(n_1302), .Y(n_1301) );
INVx1_ASAP7_75t_L g1775 ( .A(n_261), .Y(n_1775) );
CKINVDCx5p33_ASAP7_75t_R g1200 ( .A(n_262), .Y(n_1200) );
INVxp67_ASAP7_75t_SL g1078 ( .A(n_264), .Y(n_1078) );
AOI211xp5_ASAP7_75t_L g1498 ( .A1(n_266), .A2(n_509), .B(n_1499), .C(n_1501), .Y(n_1498) );
INVx1_ASAP7_75t_L g1529 ( .A(n_266), .Y(n_1529) );
CKINVDCx5p33_ASAP7_75t_R g1836 ( .A(n_268), .Y(n_1836) );
AOI22xp5_ASAP7_75t_L g1559 ( .A1(n_269), .A2(n_333), .B1(n_1544), .B2(n_1549), .Y(n_1559) );
AO22x1_ASAP7_75t_L g1564 ( .A1(n_270), .A2(n_278), .B1(n_1552), .B2(n_1561), .Y(n_1564) );
INVx1_ASAP7_75t_L g479 ( .A(n_271), .Y(n_479) );
INVx1_ASAP7_75t_L g505 ( .A(n_271), .Y(n_505) );
INVx1_ASAP7_75t_L g661 ( .A(n_272), .Y(n_661) );
INVx1_ASAP7_75t_L g451 ( .A(n_274), .Y(n_451) );
INVxp67_ASAP7_75t_SL g551 ( .A(n_275), .Y(n_551) );
CKINVDCx5p33_ASAP7_75t_R g1317 ( .A(n_276), .Y(n_1317) );
INVxp67_ASAP7_75t_SL g963 ( .A(n_277), .Y(n_963) );
INVx1_ASAP7_75t_L g783 ( .A(n_279), .Y(n_783) );
INVxp67_ASAP7_75t_SL g1788 ( .A(n_280), .Y(n_1788) );
INVx1_ASAP7_75t_L g861 ( .A(n_281), .Y(n_861) );
INVx1_ASAP7_75t_L g786 ( .A(n_283), .Y(n_786) );
INVx1_ASAP7_75t_L g1146 ( .A(n_285), .Y(n_1146) );
NOR2xp33_ASAP7_75t_L g1151 ( .A(n_285), .B(n_927), .Y(n_1151) );
INVx1_ASAP7_75t_L g1354 ( .A(n_286), .Y(n_1354) );
CKINVDCx5p33_ASAP7_75t_R g1474 ( .A(n_287), .Y(n_1474) );
INVx1_ASAP7_75t_L g775 ( .A(n_288), .Y(n_775) );
INVx1_ASAP7_75t_L g1205 ( .A(n_289), .Y(n_1205) );
CKINVDCx5p33_ASAP7_75t_R g1831 ( .A(n_290), .Y(n_1831) );
INVx1_ASAP7_75t_L g1548 ( .A(n_291), .Y(n_1548) );
AND2x2_ASAP7_75t_L g1553 ( .A(n_291), .B(n_1547), .Y(n_1553) );
INVx1_ASAP7_75t_L g1094 ( .A(n_292), .Y(n_1094) );
INVx1_ASAP7_75t_L g1820 ( .A(n_293), .Y(n_1820) );
OAI22xp33_ASAP7_75t_L g737 ( .A1(n_295), .A2(n_343), .B1(n_738), .B2(n_741), .Y(n_737) );
OAI22xp33_ASAP7_75t_L g836 ( .A1(n_295), .A2(n_343), .B1(n_361), .B2(n_837), .Y(n_836) );
AOI221xp5_ASAP7_75t_SL g1433 ( .A1(n_297), .A2(n_299), .B1(n_1061), .B2(n_1434), .C(n_1435), .Y(n_1433) );
AOI21xp33_ASAP7_75t_L g1045 ( .A1(n_298), .A2(n_588), .B(n_590), .Y(n_1045) );
INVx1_ASAP7_75t_L g1418 ( .A(n_299), .Y(n_1418) );
OAI22xp5_ASAP7_75t_L g1396 ( .A1(n_301), .A2(n_1397), .B1(n_1398), .B2(n_1449), .Y(n_1396) );
INVx1_ASAP7_75t_L g1449 ( .A(n_301), .Y(n_1449) );
INVx1_ASAP7_75t_L g857 ( .A(n_302), .Y(n_857) );
INVx1_ASAP7_75t_L g723 ( .A(n_303), .Y(n_723) );
INVx1_ASAP7_75t_L g633 ( .A(n_304), .Y(n_633) );
INVx1_ASAP7_75t_L g1233 ( .A(n_305), .Y(n_1233) );
INVx1_ASAP7_75t_L g1500 ( .A(n_306), .Y(n_1500) );
AOI211xp5_ASAP7_75t_SL g1855 ( .A1(n_308), .A2(n_422), .B(n_1856), .C(n_1858), .Y(n_1855) );
INVx1_ASAP7_75t_L g1299 ( .A(n_309), .Y(n_1299) );
XNOR2xp5_ASAP7_75t_L g1759 ( .A(n_310), .B(n_1760), .Y(n_1759) );
INVx1_ASAP7_75t_L g1189 ( .A(n_312), .Y(n_1189) );
OAI221xp5_ASAP7_75t_L g1214 ( .A1(n_312), .A2(n_703), .B1(n_721), .B2(n_1215), .C(n_1217), .Y(n_1214) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_313), .A2(n_322), .B1(n_506), .B2(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g950 ( .A(n_314), .Y(n_950) );
INVx1_ASAP7_75t_L g754 ( .A(n_315), .Y(n_754) );
INVx1_ASAP7_75t_L g1524 ( .A(n_316), .Y(n_1524) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_317), .Y(n_365) );
INVx1_ASAP7_75t_L g942 ( .A(n_318), .Y(n_942) );
CKINVDCx5p33_ASAP7_75t_R g1459 ( .A(n_319), .Y(n_1459) );
CKINVDCx5p33_ASAP7_75t_R g1368 ( .A(n_320), .Y(n_1368) );
INVx1_ASAP7_75t_L g1436 ( .A(n_321), .Y(n_1436) );
AOI21xp33_ASAP7_75t_L g1800 ( .A1(n_325), .A2(n_570), .B(n_872), .Y(n_1800) );
INVx1_ASAP7_75t_L g653 ( .A(n_326), .Y(n_653) );
CKINVDCx5p33_ASAP7_75t_R g1314 ( .A(n_327), .Y(n_1314) );
INVx1_ASAP7_75t_L g1171 ( .A(n_329), .Y(n_1171) );
XOR2xp5_ASAP7_75t_L g1452 ( .A(n_331), .B(n_1453), .Y(n_1452) );
INVx1_ASAP7_75t_L g385 ( .A(n_332), .Y(n_385) );
INVx1_ASAP7_75t_L g398 ( .A(n_332), .Y(n_398) );
INVx2_ASAP7_75t_L g431 ( .A(n_332), .Y(n_431) );
XOR2x2_ASAP7_75t_L g844 ( .A(n_333), .B(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g1032 ( .A(n_334), .Y(n_1032) );
INVx1_ASAP7_75t_L g1791 ( .A(n_335), .Y(n_1791) );
INVx1_ASAP7_75t_L g1357 ( .A(n_336), .Y(n_1357) );
CKINVDCx5p33_ASAP7_75t_R g1191 ( .A(n_337), .Y(n_1191) );
OAI21xp33_ASAP7_75t_SL g926 ( .A1(n_338), .A2(n_927), .B(n_928), .Y(n_926) );
INVx1_ASAP7_75t_L g935 ( .A(n_338), .Y(n_935) );
INVx1_ASAP7_75t_L g870 ( .A(n_339), .Y(n_870) );
CKINVDCx5p33_ASAP7_75t_R g1822 ( .A(n_341), .Y(n_1822) );
INVx1_ASAP7_75t_L g778 ( .A(n_342), .Y(n_778) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_370), .B(n_1535), .Y(n_344) );
INVx2_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_355), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g1813 ( .A(n_349), .B(n_358), .Y(n_1813) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g1809 ( .A(n_351), .B(n_354), .Y(n_1809) );
INVx1_ASAP7_75t_L g1869 ( .A(n_351), .Y(n_1869) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g1871 ( .A(n_354), .B(n_1869), .Y(n_1871) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_357), .B(n_360), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x4_ASAP7_75t_L g840 ( .A(n_358), .B(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x4_ASAP7_75t_L g458 ( .A(n_359), .B(n_369), .Y(n_458) );
AND2x4_ASAP7_75t_L g591 ( .A(n_359), .B(n_368), .Y(n_591) );
INVx1_ASAP7_75t_L g904 ( .A(n_360), .Y(n_904) );
AND2x4_ASAP7_75t_SL g1812 ( .A(n_360), .B(n_1813), .Y(n_1812) );
INVx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x6_ASAP7_75t_L g361 ( .A(n_362), .B(n_367), .Y(n_361) );
INVx1_ASAP7_75t_L g774 ( .A(n_362), .Y(n_774) );
OR2x6_ASAP7_75t_L g831 ( .A(n_362), .B(n_832), .Y(n_831) );
BUFx4f_ASAP7_75t_L g1313 ( .A(n_362), .Y(n_1313) );
INVxp67_ASAP7_75t_L g1327 ( .A(n_362), .Y(n_1327) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx4f_ASAP7_75t_L g562 ( .A(n_363), .Y(n_562) );
INVx3_ASAP7_75t_L g700 ( .A(n_363), .Y(n_700) );
INVx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVx2_ASAP7_75t_L g390 ( .A(n_365), .Y(n_390) );
INVx2_ASAP7_75t_L g409 ( .A(n_365), .Y(n_409) );
NAND2x1_ASAP7_75t_L g414 ( .A(n_365), .B(n_366), .Y(n_414) );
AND2x2_ASAP7_75t_L g420 ( .A(n_365), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g424 ( .A(n_365), .B(n_366), .Y(n_424) );
INVx1_ASAP7_75t_L g450 ( .A(n_365), .Y(n_450) );
INVx1_ASAP7_75t_L g391 ( .A(n_366), .Y(n_391) );
AND2x2_ASAP7_75t_L g408 ( .A(n_366), .B(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g421 ( .A(n_366), .Y(n_421) );
BUFx2_ASAP7_75t_L g444 ( .A(n_366), .Y(n_444) );
OR2x2_ASAP7_75t_L g566 ( .A(n_366), .B(n_390), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_366), .B(n_409), .Y(n_711) );
INVxp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g819 ( .A(n_368), .Y(n_819) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g823 ( .A(n_369), .Y(n_823) );
AND2x4_ASAP7_75t_L g827 ( .A(n_369), .B(n_449), .Y(n_827) );
XNOR2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_1116), .Y(n_370) );
XNOR2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_920), .Y(n_371) );
XOR2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_726), .Y(n_372) );
OAI22xp33_ASAP7_75t_SL g373 ( .A1(n_374), .A2(n_375), .B1(n_553), .B2(n_725), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI21x1_ASAP7_75t_SL g375 ( .A1(n_376), .A2(n_377), .B(n_552), .Y(n_375) );
NAND4xp25_ASAP7_75t_L g552 ( .A(n_376), .B(n_379), .C(n_392), .D(n_468), .Y(n_552) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND3xp33_ASAP7_75t_L g378 ( .A(n_379), .B(n_392), .C(n_468), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_380), .A2(n_451), .B1(n_540), .B2(n_541), .Y(n_539) );
AOI22xp33_ASAP7_75t_SL g722 ( .A1(n_381), .A2(n_548), .B1(n_723), .B2(n_724), .Y(n_722) );
INVx3_ASAP7_75t_L g927 ( .A(n_381), .Y(n_927) );
AOI222xp33_ASAP7_75t_L g1176 ( .A1(n_381), .A2(n_548), .B1(n_1177), .B2(n_1178), .C1(n_1180), .C2(n_1181), .Y(n_1176) );
NAND2xp5_ASAP7_75t_L g1337 ( .A(n_381), .B(n_1338), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g1381 ( .A(n_381), .B(n_1378), .Y(n_1381) );
AOI211xp5_ASAP7_75t_L g1787 ( .A1(n_381), .A2(n_1788), .B(n_1789), .C(n_1793), .Y(n_1787) );
AND2x4_ASAP7_75t_L g381 ( .A(n_382), .B(n_386), .Y(n_381) );
AND2x4_ASAP7_75t_L g548 ( .A(n_382), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g447 ( .A(n_383), .B(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g718 ( .A(n_383), .B(n_448), .Y(n_718) );
INVx1_ASAP7_75t_L g841 ( .A(n_383), .Y(n_841) );
INVxp67_ASAP7_75t_L g991 ( .A(n_383), .Y(n_991) );
BUFx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g461 ( .A(n_384), .Y(n_461) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx6f_ASAP7_75t_L g1031 ( .A(n_386), .Y(n_1031) );
AND2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_387), .B(n_398), .Y(n_405) );
AND2x2_ASAP7_75t_L g549 ( .A(n_387), .B(n_550), .Y(n_549) );
BUFx2_ASAP7_75t_L g572 ( .A(n_387), .Y(n_572) );
AND2x4_ASAP7_75t_L g1021 ( .A(n_387), .B(n_456), .Y(n_1021) );
AND2x4_ASAP7_75t_L g1033 ( .A(n_387), .B(n_550), .Y(n_1033) );
AND2x4_ASAP7_75t_SL g1038 ( .A(n_387), .B(n_423), .Y(n_1038) );
HB1xp67_ASAP7_75t_L g832 ( .A(n_388), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_389), .B(n_400), .Y(n_399) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_389), .Y(n_427) );
INVx3_ASAP7_75t_L g714 ( .A(n_389), .Y(n_714) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
HB1xp67_ASAP7_75t_L g1853 ( .A(n_390), .Y(n_1853) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_393), .B(n_415), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x4_ASAP7_75t_L g986 ( .A(n_396), .B(n_616), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g1220 ( .A(n_396), .B(n_1221), .Y(n_1220) );
OR2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_399), .Y(n_396) );
AND2x4_ASAP7_75t_L g622 ( .A(n_397), .B(n_480), .Y(n_622) );
INVx1_ASAP7_75t_L g978 ( .A(n_397), .Y(n_978) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g809 ( .A(n_398), .Y(n_809) );
INVx1_ASAP7_75t_L g979 ( .A(n_399), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_400), .B(n_431), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_400), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g579 ( .A(n_400), .Y(n_579) );
AND2x2_ASAP7_75t_L g581 ( .A(n_400), .B(n_582), .Y(n_581) );
AND2x6_ASAP7_75t_L g1028 ( .A(n_400), .B(n_423), .Y(n_1028) );
HB1xp67_ASAP7_75t_L g1854 ( .A(n_400), .Y(n_1854) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B1(n_410), .B2(n_411), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_402), .A2(n_528), .B1(n_532), .B2(n_542), .Y(n_527) );
INVx1_ASAP7_75t_L g720 ( .A(n_403), .Y(n_720) );
AOI21xp33_ASAP7_75t_L g964 ( .A1(n_403), .A2(n_965), .B(n_966), .Y(n_964) );
INVxp67_ASAP7_75t_L g1154 ( .A(n_403), .Y(n_1154) );
INVx1_ASAP7_75t_L g1179 ( .A(n_403), .Y(n_1179) );
AOI222xp33_ASAP7_75t_L g1333 ( .A1(n_403), .A2(n_411), .B1(n_977), .B2(n_1334), .C1(n_1335), .C2(n_1336), .Y(n_1333) );
AOI211xp5_ASAP7_75t_L g1444 ( .A1(n_403), .A2(n_1445), .B(n_1446), .C(n_1447), .Y(n_1444) );
AOI222xp33_ASAP7_75t_L g1514 ( .A1(n_403), .A2(n_411), .B1(n_977), .B2(n_1494), .C1(n_1515), .C2(n_1516), .Y(n_1514) );
AND2x4_ASAP7_75t_L g403 ( .A(n_404), .B(n_406), .Y(n_403) );
AOI332xp33_ASAP7_75t_L g1383 ( .A1(n_404), .A2(n_406), .A3(n_411), .B1(n_978), .B2(n_979), .B3(n_1374), .C1(n_1384), .C2(n_1385), .Y(n_1383) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OR2x2_ASAP7_75t_L g412 ( .A(n_405), .B(n_413), .Y(n_412) );
OR2x2_ASAP7_75t_L g721 ( .A(n_405), .B(n_413), .Y(n_721) );
INVx3_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx3_ASAP7_75t_L g428 ( .A(n_408), .Y(n_428) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_408), .Y(n_456) );
BUFx3_ASAP7_75t_L g568 ( .A(n_408), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g961 ( .A1(n_411), .A2(n_433), .B(n_943), .Y(n_961) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx3_ASAP7_75t_L g701 ( .A(n_413), .Y(n_701) );
INVx2_ASAP7_75t_SL g785 ( .A(n_413), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g1850 ( .A(n_413), .B(n_1851), .Y(n_1850) );
BUFx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_414), .Y(n_435) );
NAND3xp33_ASAP7_75t_SL g415 ( .A(n_416), .B(n_439), .C(n_452), .Y(n_415) );
AOI31xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_425), .A3(n_429), .B(n_433), .Y(n_416) );
INVx2_ASAP7_75t_L g464 ( .A(n_418), .Y(n_464) );
HB1xp67_ASAP7_75t_L g1434 ( .A(n_418), .Y(n_1434) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g1160 ( .A(n_419), .Y(n_1160) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_420), .Y(n_550) );
AND2x4_ASAP7_75t_L g838 ( .A(n_420), .B(n_832), .Y(n_838) );
BUFx3_ASAP7_75t_L g1060 ( .A(n_420), .Y(n_1060) );
BUFx3_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx3_ASAP7_75t_L g570 ( .A(n_423), .Y(n_570) );
BUFx3_ASAP7_75t_L g589 ( .A(n_423), .Y(n_589) );
AND2x2_ASAP7_75t_L g818 ( .A(n_423), .B(n_819), .Y(n_818) );
BUFx3_ASAP7_75t_L g970 ( .A(n_423), .Y(n_970) );
BUFx6f_ASAP7_75t_L g1063 ( .A(n_423), .Y(n_1063) );
INVx1_ASAP7_75t_L g1243 ( .A(n_423), .Y(n_1243) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g467 ( .A(n_424), .Y(n_467) );
HB1xp67_ASAP7_75t_L g1067 ( .A(n_426), .Y(n_1067) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx3_ASAP7_75t_L g576 ( .A(n_427), .Y(n_576) );
A2O1A1Ixp33_ASAP7_75t_L g1849 ( .A1(n_427), .A2(n_1822), .B(n_1850), .C(n_1854), .Y(n_1849) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_429), .Y(n_696) );
INVx2_ASAP7_75t_L g768 ( .A(n_429), .Y(n_768) );
INVx2_ASAP7_75t_L g872 ( .A(n_429), .Y(n_872) );
INVx4_ASAP7_75t_L g973 ( .A(n_429), .Y(n_973) );
INVx2_ASAP7_75t_L g1310 ( .A(n_429), .Y(n_1310) );
AND2x4_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
INVx1_ASAP7_75t_L g597 ( .A(n_430), .Y(n_597) );
OR2x2_ASAP7_75t_L g645 ( .A(n_430), .B(n_521), .Y(n_645) );
OR2x6_ASAP7_75t_L g1010 ( .A(n_430), .B(n_521), .Y(n_1010) );
BUFx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g469 ( .A(n_431), .Y(n_469) );
NOR3xp33_ASAP7_75t_L g1386 ( .A(n_433), .B(n_1387), .C(n_1393), .Y(n_1386) );
OR3x1_ASAP7_75t_L g1519 ( .A(n_433), .B(n_1520), .C(n_1521), .Y(n_1519) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_434), .Y(n_433) );
OAI21xp5_ASAP7_75t_L g702 ( .A1(n_434), .A2(n_703), .B(n_704), .Y(n_702) );
OAI21xp5_ASAP7_75t_L g1164 ( .A1(n_434), .A2(n_767), .B(n_1165), .Y(n_1164) );
OAI21xp5_ASAP7_75t_SL g1207 ( .A1(n_434), .A2(n_1208), .B(n_1210), .Y(n_1207) );
OR2x6_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
BUFx6f_ASAP7_75t_L g781 ( .A(n_435), .Y(n_781) );
INVx4_ASAP7_75t_L g883 ( .A(n_435), .Y(n_883) );
BUFx4f_ASAP7_75t_L g888 ( .A(n_435), .Y(n_888) );
BUFx4f_ASAP7_75t_L g1212 ( .A(n_435), .Y(n_1212) );
BUFx4f_ASAP7_75t_L g1232 ( .A(n_435), .Y(n_1232) );
BUFx4f_ASAP7_75t_L g1523 ( .A(n_435), .Y(n_1523) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2x2_ASAP7_75t_L g441 ( .A(n_437), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI22xp33_ASAP7_75t_SL g439 ( .A1(n_440), .A2(n_445), .B1(n_446), .B2(n_451), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g1217 ( .A1(n_440), .A2(n_446), .B1(n_1186), .B2(n_1188), .Y(n_1217) );
AOI22xp5_ASAP7_75t_L g1790 ( .A1(n_440), .A2(n_446), .B1(n_1791), .B2(n_1792), .Y(n_1790) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_SL g717 ( .A(n_441), .Y(n_717) );
HB1xp67_ASAP7_75t_L g1448 ( .A(n_441), .Y(n_1448) );
INVx2_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
BUFx2_ASAP7_75t_L g582 ( .A(n_444), .Y(n_582) );
AND2x4_ASAP7_75t_L g822 ( .A(n_444), .B(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g1042 ( .A(n_444), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g1851 ( .A1(n_444), .A2(n_1819), .B1(n_1835), .B2(n_1852), .Y(n_1851) );
INVx2_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
AND2x4_ASAP7_75t_L g989 ( .A(n_447), .B(n_612), .Y(n_989) );
AND2x4_ASAP7_75t_L g1087 ( .A(n_447), .B(n_612), .Y(n_1087) );
INVx1_ASAP7_75t_L g584 ( .A(n_448), .Y(n_584) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NAND3xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_457), .C(n_462), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx2_ASAP7_75t_L g596 ( .A(n_456), .Y(n_596) );
HB1xp67_ASAP7_75t_L g1027 ( .A(n_456), .Y(n_1027) );
CKINVDCx5p33_ASAP7_75t_R g703 ( .A(n_457), .Y(n_703) );
AOI332xp33_ASAP7_75t_L g967 ( .A1(n_457), .A2(n_968), .A3(n_971), .B1(n_972), .B2(n_974), .B3(n_975), .C1(n_977), .C2(n_980), .Y(n_967) );
AOI211xp5_ASAP7_75t_L g1158 ( .A1(n_457), .A2(n_1159), .B(n_1164), .C(n_1170), .Y(n_1158) );
AOI322xp5_ASAP7_75t_L g1426 ( .A1(n_457), .A2(n_977), .A3(n_1427), .B1(n_1428), .B2(n_1432), .C1(n_1433), .C2(n_1438), .Y(n_1426) );
AOI322xp5_ASAP7_75t_L g1794 ( .A1(n_457), .A2(n_977), .A3(n_1795), .B1(n_1797), .B2(n_1800), .C1(n_1801), .C2(n_1802), .Y(n_1794) );
AND2x4_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
INVx4_ASAP7_75t_L g594 ( .A(n_458), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_458), .B(n_459), .Y(n_789) );
INVx1_ASAP7_75t_SL g1024 ( .A(n_458), .Y(n_1024) );
INVx4_ASAP7_75t_L g1065 ( .A(n_458), .Y(n_1065) );
AND2x2_ASAP7_75t_SL g1331 ( .A(n_458), .B(n_461), .Y(n_1331) );
OAI21xp33_ASAP7_75t_L g1856 ( .A1(n_458), .A2(n_887), .B(n_1857), .Y(n_1856) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g604 ( .A(n_461), .B(n_531), .Y(n_604) );
OR2x2_ASAP7_75t_L g625 ( .A(n_461), .B(n_517), .Y(n_625) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_461), .Y(n_735) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g588 ( .A(n_464), .Y(n_588) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g1480 ( .A(n_467), .Y(n_1480) );
AOI22xp33_ASAP7_75t_SL g468 ( .A1(n_469), .A2(n_470), .B1(n_546), .B2(n_551), .Y(n_468) );
OAI31xp33_ASAP7_75t_SL g928 ( .A1(n_469), .A2(n_929), .A3(n_940), .B(n_944), .Y(n_928) );
AND3x4_ASAP7_75t_L g1003 ( .A(n_469), .B(n_484), .C(n_692), .Y(n_1003) );
INVx1_ASAP7_75t_L g1050 ( .A(n_469), .Y(n_1050) );
INVx2_ASAP7_75t_SL g1783 ( .A(n_469), .Y(n_1783) );
NAND3xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_497), .C(n_527), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_491), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_475), .A2(n_486), .B1(n_942), .B2(n_943), .Y(n_941) );
AOI221xp5_ASAP7_75t_L g1137 ( .A1(n_475), .A2(n_486), .B1(n_491), .B2(n_1138), .C(n_1139), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g1187 ( .A1(n_475), .A2(n_486), .B1(n_1188), .B2(n_1189), .Y(n_1187) );
INVx2_ASAP7_75t_L g1343 ( .A(n_475), .Y(n_1343) );
AOI22xp33_ASAP7_75t_L g1403 ( .A1(n_475), .A2(n_486), .B1(n_1404), .B2(n_1405), .Y(n_1403) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_480), .Y(n_475) );
INVx1_ASAP7_75t_L g620 ( .A(n_476), .Y(n_620) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x4_ASAP7_75t_L g507 ( .A(n_477), .B(n_489), .Y(n_507) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x4_ASAP7_75t_L g510 ( .A(n_478), .B(n_490), .Y(n_510) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g495 ( .A(n_479), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_479), .B(n_490), .Y(n_538) );
AND2x6_ASAP7_75t_L g486 ( .A(n_480), .B(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g496 ( .A(n_480), .Y(n_496) );
NAND2x1p5_ASAP7_75t_L g545 ( .A(n_480), .B(n_501), .Y(n_545) );
AND2x4_ASAP7_75t_L g480 ( .A(n_481), .B(n_483), .Y(n_480) );
NAND2x1p5_ASAP7_75t_L g521 ( .A(n_481), .B(n_522), .Y(n_521) );
OR2x4_ASAP7_75t_L g740 ( .A(n_481), .B(n_628), .Y(n_740) );
INVx1_ASAP7_75t_L g743 ( .A(n_481), .Y(n_743) );
AND2x4_ASAP7_75t_L g748 ( .A(n_481), .B(n_510), .Y(n_748) );
OR2x6_ASAP7_75t_L g764 ( .A(n_481), .B(n_636), .Y(n_764) );
NAND3x1_ASAP7_75t_L g808 ( .A(n_481), .B(n_522), .C(n_809), .Y(n_808) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NAND2xp33_ASAP7_75t_SL g517 ( .A(n_482), .B(n_484), .Y(n_517) );
BUFx3_ASAP7_75t_L g692 ( .A(n_482), .Y(n_692) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g691 ( .A(n_484), .B(n_692), .Y(n_691) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_484), .Y(n_733) );
INVx4_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g996 ( .A(n_487), .B(n_622), .Y(n_996) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_487), .B(n_622), .Y(n_1093) );
NAND2x1_ASAP7_75t_L g1259 ( .A(n_487), .B(n_622), .Y(n_1259) );
AND2x4_ASAP7_75t_SL g1834 ( .A(n_487), .B(n_622), .Y(n_1834) );
INVx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND2x1p5_ASAP7_75t_L g494 ( .A(n_489), .B(n_495), .Y(n_494) );
BUFx2_ASAP7_75t_L g753 ( .A(n_489), .Y(n_753) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g502 ( .A(n_490), .Y(n_502) );
OR2x2_ASAP7_75t_L g628 ( .A(n_490), .B(n_504), .Y(n_628) );
NOR3xp33_ASAP7_75t_L g1344 ( .A(n_491), .B(n_1345), .C(n_1349), .Y(n_1344) );
NOR3xp33_ASAP7_75t_L g1360 ( .A(n_491), .B(n_1361), .C(n_1366), .Y(n_1360) );
CKINVDCx5p33_ASAP7_75t_R g491 ( .A(n_492), .Y(n_491) );
OR2x6_ASAP7_75t_L g492 ( .A(n_493), .B(n_496), .Y(n_492) );
INVx1_ASAP7_75t_L g746 ( .A(n_493), .Y(n_746) );
OAI221xp5_ASAP7_75t_L g1367 ( .A1(n_493), .A2(n_520), .B1(n_627), .B2(n_1368), .C(n_1369), .Y(n_1367) );
INVx1_ASAP7_75t_L g1780 ( .A(n_493), .Y(n_1780) );
BUFx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_494), .Y(n_613) );
BUFx3_ASAP7_75t_L g621 ( .A(n_494), .Y(n_621) );
BUFx2_ASAP7_75t_L g757 ( .A(n_495), .Y(n_757) );
INVx1_ASAP7_75t_L g663 ( .A(n_496), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_508), .B1(n_518), .B2(n_523), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g618 ( .A1(n_499), .A2(n_569), .B(n_619), .C(n_622), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g1185 ( .A1(n_499), .A2(n_1129), .B1(n_1180), .B2(n_1186), .Y(n_1185) );
INVx8_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx3_ASAP7_75t_L g540 ( .A(n_500), .Y(n_540) );
INVx2_ASAP7_75t_L g602 ( .A(n_500), .Y(n_602) );
INVx2_ASAP7_75t_L g1147 ( .A(n_500), .Y(n_1147) );
INVx8_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g936 ( .A(n_501), .B(n_937), .Y(n_936) );
BUFx3_ASAP7_75t_L g1101 ( .A(n_501), .Y(n_1101) );
BUFx3_ASAP7_75t_L g1136 ( .A(n_501), .Y(n_1136) );
HB1xp67_ASAP7_75t_L g1280 ( .A(n_501), .Y(n_1280) );
AND2x4_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
AND2x4_ASAP7_75t_L g514 ( .A(n_502), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVxp67_ASAP7_75t_L g515 ( .A(n_505), .Y(n_515) );
BUFx2_ASAP7_75t_L g1106 ( .A(n_506), .Y(n_1106) );
BUFx12f_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
BUFx3_ASAP7_75t_L g652 ( .A(n_507), .Y(n_652) );
AND2x4_ASAP7_75t_L g933 ( .A(n_507), .B(n_530), .Y(n_933) );
INVx5_ASAP7_75t_L g1006 ( .A(n_507), .Y(n_1006) );
BUFx2_ASAP7_75t_L g1127 ( .A(n_507), .Y(n_1127) );
BUFx3_ASAP7_75t_L g1468 ( .A(n_507), .Y(n_1468) );
BUFx3_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
BUFx2_ASAP7_75t_L g541 ( .A(n_510), .Y(n_541) );
INVx2_ASAP7_75t_L g655 ( .A(n_510), .Y(n_655) );
AND2x2_ASAP7_75t_L g939 ( .A(n_510), .B(n_937), .Y(n_939) );
BUFx2_ASAP7_75t_L g1002 ( .A(n_510), .Y(n_1002) );
BUFx2_ASAP7_75t_L g1129 ( .A(n_510), .Y(n_1129) );
BUFx2_ASAP7_75t_L g1465 ( .A(n_510), .Y(n_1465) );
BUFx2_ASAP7_75t_L g1825 ( .A(n_510), .Y(n_1825) );
INVx8_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_512), .A2(n_633), .B1(n_634), .B2(n_637), .Y(n_632) );
INVx5_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_SL g659 ( .A(n_513), .Y(n_659) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_513), .Y(n_668) );
INVx2_ASAP7_75t_SL g1133 ( .A(n_513), .Y(n_1133) );
INVx3_ASAP7_75t_L g1144 ( .A(n_513), .Y(n_1144) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx8_ASAP7_75t_L g526 ( .A(n_514), .Y(n_526) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_514), .Y(n_534) );
INVx2_ASAP7_75t_L g609 ( .A(n_514), .Y(n_609) );
BUFx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OAI221xp5_ASAP7_75t_L g671 ( .A1(n_520), .A2(n_672), .B1(n_673), .B2(n_675), .C(n_676), .Y(n_671) );
OAI221xp5_ASAP7_75t_L g952 ( .A1(n_520), .A2(n_658), .B1(n_687), .B2(n_953), .C(n_954), .Y(n_952) );
OAI221xp5_ASAP7_75t_L g1197 ( .A1(n_520), .A2(n_851), .B1(n_1198), .B2(n_1200), .C(n_1201), .Y(n_1197) );
OAI221xp5_ASAP7_75t_L g1350 ( .A1(n_520), .A2(n_621), .B1(n_658), .B2(n_1314), .C(n_1324), .Y(n_1350) );
OAI221xp5_ASAP7_75t_L g1509 ( .A1(n_520), .A2(n_621), .B1(n_658), .B2(n_1510), .C(n_1511), .Y(n_1509) );
NAND2xp5_ASAP7_75t_L g1781 ( .A(n_520), .B(n_1782), .Y(n_1781) );
INVx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OAI221xp5_ASAP7_75t_L g945 ( .A1(n_525), .A2(n_631), .B1(n_691), .B2(n_946), .C(n_947), .Y(n_945) );
OAI22xp5_ASAP7_75t_L g955 ( .A1(n_525), .A2(n_956), .B1(n_957), .B2(n_958), .Y(n_955) );
OAI21xp33_ASAP7_75t_L g1499 ( .A1(n_525), .A2(n_691), .B(n_1500), .Y(n_1499) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x4_ASAP7_75t_L g1016 ( .A(n_526), .B(n_603), .Y(n_1016) );
INVx3_ASAP7_75t_L g1109 ( .A(n_526), .Y(n_1109) );
INVx2_ASAP7_75t_SL g1203 ( .A(n_526), .Y(n_1203) );
INVx1_ASAP7_75t_L g650 ( .A(n_528), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g1340 ( .A1(n_528), .A2(n_544), .B1(n_1335), .B2(n_1341), .C(n_1342), .Y(n_1340) );
AOI221xp5_ASAP7_75t_L g1373 ( .A1(n_528), .A2(n_544), .B1(n_1374), .B2(n_1375), .C(n_1379), .Y(n_1373) );
BUFx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g1142 ( .A(n_529), .Y(n_1142) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g931 ( .A(n_530), .Y(n_931) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g937 ( .A(n_531), .Y(n_937) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_534), .Y(n_689) );
AND2x4_ASAP7_75t_L g742 ( .A(n_534), .B(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g856 ( .A(n_534), .Y(n_856) );
INVx2_ASAP7_75t_L g1365 ( .A(n_534), .Y(n_1365) );
BUFx6f_ASAP7_75t_L g1417 ( .A(n_534), .Y(n_1417) );
INVx1_ASAP7_75t_L g1770 ( .A(n_534), .Y(n_1770) );
OAI22xp5_ASAP7_75t_L g1202 ( .A1(n_535), .A2(n_1203), .B1(n_1204), .B2(n_1205), .Y(n_1202) );
CKINVDCx8_ASAP7_75t_R g535 ( .A(n_536), .Y(n_535) );
INVx3_ASAP7_75t_L g804 ( .A(n_536), .Y(n_804) );
INVx3_ASAP7_75t_L g858 ( .A(n_536), .Y(n_858) );
INVx3_ASAP7_75t_L g951 ( .A(n_536), .Y(n_951) );
INVx1_ASAP7_75t_L g1503 ( .A(n_536), .Y(n_1503) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g617 ( .A(n_537), .Y(n_617) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx2_ASAP7_75t_L g636 ( .A(n_538), .Y(n_636) );
A2O1A1Ixp33_ASAP7_75t_L g660 ( .A1(n_540), .A2(n_661), .B(n_662), .C(n_663), .Y(n_660) );
AND2x4_ASAP7_75t_L g1017 ( .A(n_541), .B(n_622), .Y(n_1017) );
BUFx2_ASAP7_75t_L g1102 ( .A(n_541), .Y(n_1102) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_544), .A2(n_1141), .B1(n_1143), .B2(n_1149), .Y(n_1140) );
AOI211xp5_ASAP7_75t_L g1493 ( .A1(n_544), .A2(n_1494), .B(n_1495), .C(n_1496), .Y(n_1493) );
AOI211xp5_ASAP7_75t_SL g1763 ( .A1(n_544), .A2(n_1764), .B(n_1765), .C(n_1766), .Y(n_1763) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g990 ( .A(n_545), .B(n_991), .Y(n_990) );
OR2x6_ASAP7_75t_L g1088 ( .A(n_545), .B(n_991), .Y(n_1088) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_548), .B(n_963), .Y(n_962) );
HB1xp67_ASAP7_75t_L g1157 ( .A(n_548), .Y(n_1157) );
NAND2xp33_ASAP7_75t_SL g1353 ( .A(n_548), .B(n_1354), .Y(n_1353) );
INVx1_ASAP7_75t_L g1442 ( .A(n_548), .Y(n_1442) );
NAND2xp5_ASAP7_75t_L g1517 ( .A(n_548), .B(n_1518), .Y(n_1517) );
NAND2xp5_ASAP7_75t_L g1784 ( .A(n_548), .B(n_1785), .Y(n_1784) );
BUFx6f_ASAP7_75t_L g969 ( .A(n_550), .Y(n_969) );
INVx2_ASAP7_75t_L g1847 ( .A(n_550), .Y(n_1847) );
INVx1_ASAP7_75t_L g725 ( .A(n_553), .Y(n_725) );
XNOR2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_646), .Y(n_553) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_598), .Y(n_557) );
AOI21xp5_ASAP7_75t_SL g558 ( .A1(n_559), .A2(n_586), .B(n_597), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_572), .B(n_573), .Y(n_559) );
OAI22xp33_ASAP7_75t_L g1161 ( .A1(n_561), .A2(n_707), .B1(n_1162), .B2(n_1163), .Y(n_1161) );
INVx3_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx6f_ASAP7_75t_L g792 ( .A(n_562), .Y(n_792) );
INVx4_ASAP7_75t_L g1860 ( .A(n_562), .Y(n_1860) );
OAI22xp5_ASAP7_75t_L g1522 ( .A1(n_563), .A2(n_1500), .B1(n_1523), .B2(n_1524), .Y(n_1522) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g779 ( .A(n_564), .Y(n_779) );
INVx4_ASAP7_75t_L g1318 ( .A(n_564), .Y(n_1318) );
INVx4_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
BUFx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g706 ( .A(n_566), .Y(n_706) );
INVx2_ASAP7_75t_L g880 ( .A(n_566), .Y(n_880) );
BUFx3_ASAP7_75t_L g887 ( .A(n_566), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_569), .B1(n_570), .B2(n_571), .Y(n_567) );
INVx1_ASAP7_75t_SL g1431 ( .A(n_568), .Y(n_1431) );
A2O1A1Ixp33_ASAP7_75t_L g574 ( .A1(n_570), .A2(n_575), .B(n_577), .C(n_578), .Y(n_574) );
INVxp67_ASAP7_75t_L g1844 ( .A(n_572), .Y(n_1844) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_580), .Y(n_573) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g1297 ( .A(n_576), .Y(n_1297) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NOR2x1_ASAP7_75t_L g1041 ( .A(n_579), .B(n_1042), .Y(n_1041) );
AOI22xp33_ASAP7_75t_SL g580 ( .A1(n_581), .A2(n_583), .B1(n_584), .B2(n_585), .Y(n_580) );
AOI222xp33_ASAP7_75t_L g1290 ( .A1(n_581), .A2(n_1286), .B1(n_1287), .B2(n_1291), .C1(n_1292), .C2(n_1293), .Y(n_1290) );
INVx1_ASAP7_75t_L g1487 ( .A(n_581), .Y(n_1487) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_585), .A2(n_606), .B1(n_607), .B2(n_611), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_592), .B1(n_593), .B2(n_595), .Y(n_586) );
INVx3_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g1082 ( .A(n_591), .Y(n_1082) );
OAI221xp5_ASAP7_75t_L g1231 ( .A1(n_591), .A2(n_885), .B1(n_1232), .B2(n_1233), .C(n_1234), .Y(n_1231) );
INVx1_ASAP7_75t_L g1484 ( .A(n_591), .Y(n_1484) );
OAI221xp5_ASAP7_75t_L g1839 ( .A1(n_591), .A2(n_1391), .B1(n_1840), .B2(n_1841), .C(n_1842), .Y(n_1839) );
INVx1_ASAP7_75t_L g694 ( .A(n_597), .Y(n_694) );
BUFx2_ASAP7_75t_L g1150 ( .A(n_597), .Y(n_1150) );
NAND2xp5_ASAP7_75t_L g1221 ( .A(n_597), .B(n_933), .Y(n_1221) );
NAND3xp33_ASAP7_75t_SL g598 ( .A(n_599), .B(n_605), .C(n_614), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g1489 ( .A1(n_601), .A2(n_1016), .B1(n_1473), .B2(n_1474), .Y(n_1489) );
AND2x4_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
AND2x4_ASAP7_75t_L g1251 ( .A(n_602), .B(n_603), .Y(n_1251) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g610 ( .A(n_604), .Y(n_610) );
OR2x2_ASAP7_75t_L g612 ( .A(n_604), .B(n_613), .Y(n_612) );
OR2x2_ASAP7_75t_L g616 ( .A(n_604), .B(n_617), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g1250 ( .A1(n_607), .A2(n_1246), .B1(n_1247), .B2(n_1251), .Y(n_1250) );
AOI22xp33_ASAP7_75t_L g1302 ( .A1(n_607), .A2(n_1251), .B1(n_1299), .B2(n_1300), .Y(n_1302) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
INVx2_ASAP7_75t_L g639 ( .A(n_608), .Y(n_639) );
INVx2_ASAP7_75t_L g1376 ( .A(n_608), .Y(n_1376) );
INVx3_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
BUFx2_ASAP7_75t_L g860 ( .A(n_609), .Y(n_860) );
OR2x6_ASAP7_75t_SL g930 ( .A(n_609), .B(n_931), .Y(n_930) );
BUFx2_ASAP7_75t_L g1105 ( .A(n_609), .Y(n_1105) );
INVxp67_ASAP7_75t_L g1014 ( .A(n_610), .Y(n_1014) );
AOI222xp33_ASAP7_75t_L g1818 ( .A1(n_611), .A2(n_1251), .B1(n_1819), .B2(n_1820), .C1(n_1821), .C2(n_1822), .Y(n_1818) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_613), .Y(n_631) );
INVx4_ASAP7_75t_L g674 ( .A(n_613), .Y(n_674) );
INVx3_ASAP7_75t_L g813 ( .A(n_613), .Y(n_813) );
OAI221xp5_ASAP7_75t_L g1362 ( .A1(n_613), .A2(n_691), .B1(n_1363), .B2(n_1364), .C(n_1365), .Y(n_1362) );
NOR2xp33_ASAP7_75t_SL g614 ( .A(n_615), .B(n_623), .Y(n_614) );
INVx1_ASAP7_75t_L g1821 ( .A(n_616), .Y(n_1821) );
BUFx3_ASAP7_75t_L g862 ( .A(n_617), .Y(n_862) );
INVx1_ASAP7_75t_L g959 ( .A(n_617), .Y(n_959) );
INVx2_ASAP7_75t_L g999 ( .A(n_620), .Y(n_999) );
OAI22xp33_ASAP7_75t_L g642 ( .A1(n_621), .A2(n_627), .B1(n_643), .B2(n_644), .Y(n_642) );
BUFx6f_ASAP7_75t_L g869 ( .A(n_621), .Y(n_869) );
INVx2_ASAP7_75t_L g1199 ( .A(n_621), .Y(n_1199) );
OAI221xp5_ASAP7_75t_L g1348 ( .A1(n_621), .A2(n_639), .B1(n_691), .B2(n_1319), .C(n_1323), .Y(n_1348) );
AND2x4_ASAP7_75t_L g998 ( .A(n_622), .B(n_999), .Y(n_998) );
AND2x4_ASAP7_75t_SL g1261 ( .A(n_622), .B(n_999), .Y(n_1261) );
OAI33xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_626), .A3(n_632), .B1(n_638), .B2(n_642), .B3(n_645), .Y(n_623) );
BUFx3_ASAP7_75t_L g798 ( .A(n_624), .Y(n_798) );
BUFx4f_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
BUFx2_ASAP7_75t_L g848 ( .A(n_625), .Y(n_848) );
OAI22xp33_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_629), .B1(n_630), .B2(n_631), .Y(n_626) );
INVx1_ASAP7_75t_L g852 ( .A(n_627), .Y(n_852) );
BUFx4f_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
BUFx3_ASAP7_75t_L g658 ( .A(n_628), .Y(n_658) );
BUFx3_ASAP7_75t_L g675 ( .A(n_628), .Y(n_675) );
INVx2_ASAP7_75t_L g681 ( .A(n_628), .Y(n_681) );
OR2x4_ASAP7_75t_L g761 ( .A(n_628), .B(n_743), .Y(n_761) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_631), .Y(n_802) );
OAI22xp33_ASAP7_75t_L g849 ( .A1(n_631), .A2(n_850), .B1(n_851), .B2(n_853), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_634), .A2(n_639), .B1(n_640), .B2(n_641), .Y(n_638) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
BUFx2_ASAP7_75t_L g684 ( .A(n_635), .Y(n_684) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
BUFx3_ASAP7_75t_L g670 ( .A(n_636), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_639), .A2(n_670), .B1(n_780), .B2(n_796), .Y(n_805) );
NAND4xp75_ASAP7_75t_L g647 ( .A(n_648), .B(n_695), .C(n_719), .D(n_722), .Y(n_647) );
OAI21x1_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_664), .B(n_693), .Y(n_648) );
OAI21xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_651), .B(n_660), .Y(n_649) );
AOI221xp5_ASAP7_75t_SL g651 ( .A1(n_652), .A2(n_653), .B1(n_654), .B2(n_656), .C(n_657), .Y(n_651) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g1281 ( .A(n_655), .Y(n_1281) );
INVx1_ASAP7_75t_L g1829 ( .A(n_655), .Y(n_1829) );
INVx1_ASAP7_75t_L g801 ( .A(n_658), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_659), .A2(n_778), .B1(n_793), .B2(n_804), .Y(n_803) );
INVx2_ASAP7_75t_L g1130 ( .A(n_659), .Y(n_1130) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_671), .B1(n_677), .B2(n_685), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_667), .B1(n_669), .B2(n_670), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_666), .A2(n_678), .B1(n_699), .B2(n_701), .Y(n_698) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
OAI221xp5_ASAP7_75t_L g704 ( .A1(n_669), .A2(n_686), .B1(n_705), .B2(n_707), .C(n_712), .Y(n_704) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g687 ( .A(n_674), .Y(n_687) );
INVx2_ASAP7_75t_L g1772 ( .A(n_674), .Y(n_1772) );
OAI22xp5_ASAP7_75t_L g1501 ( .A1(n_675), .A2(n_1502), .B1(n_1503), .B2(n_1504), .Y(n_1501) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B1(n_682), .B2(n_683), .Y(n_677) );
BUFx4f_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g948 ( .A1(n_680), .A2(n_949), .B1(n_950), .B2(n_951), .Y(n_948) );
INVx3_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx2_ASAP7_75t_SL g811 ( .A(n_681), .Y(n_811) );
INVx3_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
OAI221xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_687), .B1(n_688), .B2(n_690), .C(n_691), .Y(n_685) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OAI221xp5_ASAP7_75t_L g1773 ( .A1(n_691), .A2(n_1006), .B1(n_1100), .B2(n_1774), .C(n_1775), .Y(n_1773) );
INVx3_ASAP7_75t_L g752 ( .A(n_692), .Y(n_752) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AOI211x1_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B(n_702), .C(n_715), .Y(n_695) );
INVx1_ASAP7_75t_L g875 ( .A(n_699), .Y(n_875) );
BUFx3_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
BUFx3_ASAP7_75t_L g1532 ( .A(n_700), .Y(n_1532) );
BUFx2_ASAP7_75t_L g816 ( .A(n_701), .Y(n_816) );
OAI22xp5_ASAP7_75t_L g1320 ( .A1(n_701), .A2(n_1321), .B1(n_1323), .B2(n_1324), .Y(n_1320) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx6_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx5_ASAP7_75t_L g776 ( .A(n_708), .Y(n_776) );
BUFx6f_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g795 ( .A(n_709), .Y(n_795) );
INVx4_ASAP7_75t_L g877 ( .A(n_709), .Y(n_877) );
INVx1_ASAP7_75t_L g1079 ( .A(n_709), .Y(n_1079) );
INVx2_ASAP7_75t_SL g1315 ( .A(n_709), .Y(n_1315) );
INVx2_ASAP7_75t_L g1527 ( .A(n_709), .Y(n_1527) );
INVx8_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
OR2x2_ASAP7_75t_L g835 ( .A(n_710), .B(n_823), .Y(n_835) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_SL g976 ( .A(n_714), .Y(n_976) );
INVx2_ASAP7_75t_L g1026 ( .A(n_714), .Y(n_1026) );
INVx1_ASAP7_75t_L g1429 ( .A(n_714), .Y(n_1429) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_728), .B1(n_844), .B2(n_919), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g842 ( .A(n_729), .Y(n_842) );
OAI211xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_736), .B(n_765), .C(n_814), .Y(n_729) );
CKINVDCx14_ASAP7_75t_R g730 ( .A(n_731), .Y(n_730) );
AND2x4_ASAP7_75t_L g731 ( .A(n_732), .B(n_734), .Y(n_731) );
AND2x2_ASAP7_75t_SL g918 ( .A(n_732), .B(n_734), .Y(n_918) );
INVx1_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NOR3xp33_ASAP7_75t_SL g736 ( .A(n_737), .B(n_744), .C(n_759), .Y(n_736) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g908 ( .A(n_742), .Y(n_908) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
CKINVDCx8_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_754), .B1(n_755), .B2(n_758), .Y(n_749) );
BUFx3_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
BUFx3_ASAP7_75t_L g911 ( .A(n_751), .Y(n_911) );
AND2x2_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
AND2x4_ASAP7_75t_L g756 ( .A(n_752), .B(n_757), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_754), .A2(n_821), .B1(n_824), .B2(n_825), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_755), .A2(n_895), .B1(n_911), .B2(n_912), .Y(n_910) );
BUFx6f_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
BUFx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx2_ASAP7_75t_SL g915 ( .A(n_761), .Y(n_915) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
BUFx3_ASAP7_75t_L g916 ( .A(n_764), .Y(n_916) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_797), .Y(n_765) );
OAI33xp33_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_769), .A3(n_777), .B1(n_782), .B2(n_787), .B3(n_790), .Y(n_766) );
INVx1_ASAP7_75t_L g1438 ( .A(n_767), .Y(n_1438) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
OAI22xp33_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_771), .B1(n_775), .B2(n_776), .Y(n_769) );
OAI22xp33_ASAP7_75t_L g799 ( .A1(n_770), .A2(n_783), .B1(n_800), .B2(n_802), .Y(n_799) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_775), .A2(n_786), .B1(n_811), .B2(n_812), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g1798 ( .A1(n_776), .A2(n_1313), .B1(n_1775), .B2(n_1799), .Y(n_1798) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_779), .B1(n_780), .B2(n_781), .Y(n_777) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_779), .A2(n_783), .B1(n_784), .B2(n_786), .Y(n_782) );
OAI221xp5_ASAP7_75t_L g1215 ( .A1(n_779), .A2(n_888), .B1(n_1191), .B2(n_1200), .C(n_1216), .Y(n_1215) );
OAI221xp5_ASAP7_75t_L g1390 ( .A1(n_781), .A2(n_1363), .B1(n_1368), .B2(n_1391), .C(n_1392), .Y(n_1390) );
INVx5_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
OAI33xp33_ASAP7_75t_L g871 ( .A1(n_787), .A2(n_872), .A3(n_873), .B1(n_878), .B2(n_884), .B3(n_889), .Y(n_871) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
OAI22xp5_ASAP7_75t_SL g1387 ( .A1(n_789), .A2(n_1310), .B1(n_1388), .B2(n_1390), .Y(n_1387) );
OAI22xp5_ASAP7_75t_L g790 ( .A1(n_791), .A2(n_793), .B1(n_794), .B2(n_796), .Y(n_790) );
INVx2_ASAP7_75t_SL g791 ( .A(n_792), .Y(n_791) );
INVx2_ASAP7_75t_L g1077 ( .A(n_792), .Y(n_1077) );
INVx2_ASAP7_75t_L g1237 ( .A(n_792), .Y(n_1237) );
INVx3_ASAP7_75t_L g1526 ( .A(n_792), .Y(n_1526) );
OAI22xp5_ASAP7_75t_L g1235 ( .A1(n_794), .A2(n_1236), .B1(n_1237), .B2(n_1238), .Y(n_1235) );
BUFx3_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
OAI33xp33_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_799), .A3(n_803), .B1(n_805), .B2(n_806), .B3(n_810), .Y(n_797) );
INVx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
AOI33xp33_ASAP7_75t_L g1095 ( .A1(n_807), .A2(n_1096), .A3(n_1097), .B1(n_1103), .B2(n_1107), .B3(n_1111), .Y(n_1095) );
INVx3_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx3_ASAP7_75t_L g866 ( .A(n_808), .Y(n_866) );
OR2x2_ASAP7_75t_L g1013 ( .A(n_811), .B(n_1014), .Y(n_1013) );
OR2x6_ASAP7_75t_L g1113 ( .A(n_811), .B(n_1014), .Y(n_1113) );
INVx2_ASAP7_75t_SL g1409 ( .A(n_811), .Y(n_1409) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx2_ASAP7_75t_L g1193 ( .A(n_813), .Y(n_1193) );
OAI31xp33_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_828), .A3(n_836), .B(n_839), .Y(n_814) );
INVx3_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
BUFx3_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_822), .A2(n_895), .B1(n_896), .B2(n_897), .Y(n_894) );
INVx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx2_ASAP7_75t_L g898 ( .A(n_827), .Y(n_898) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
HB1xp67_ASAP7_75t_L g900 ( .A(n_831), .Y(n_900) );
HB1xp67_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
BUFx2_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx2_ASAP7_75t_L g902 ( .A(n_835), .Y(n_902) );
CKINVDCx16_ASAP7_75t_R g837 ( .A(n_838), .Y(n_837) );
INVx3_ASAP7_75t_SL g905 ( .A(n_838), .Y(n_905) );
OAI31xp33_ASAP7_75t_L g892 ( .A1(n_839), .A2(n_893), .A3(n_899), .B(n_903), .Y(n_892) );
BUFx3_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g919 ( .A(n_844), .Y(n_919) );
NAND3xp33_ASAP7_75t_L g845 ( .A(n_846), .B(n_892), .C(n_906), .Y(n_845) );
NOR2xp33_ASAP7_75t_L g846 ( .A(n_847), .B(n_871), .Y(n_846) );
OAI33xp33_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_849), .A3(n_854), .B1(n_859), .B2(n_864), .B3(n_867), .Y(n_847) );
OAI22xp5_ASAP7_75t_SL g873 ( .A1(n_850), .A2(n_868), .B1(n_874), .B2(n_876), .Y(n_873) );
OAI22xp33_ASAP7_75t_L g867 ( .A1(n_851), .A2(n_868), .B1(n_869), .B2(n_870), .Y(n_867) );
INVx2_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_853), .A2(n_870), .B1(n_885), .B2(n_888), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_855), .A2(n_856), .B1(n_857), .B2(n_858), .Y(n_854) );
OAI22xp5_ASAP7_75t_L g878 ( .A1(n_855), .A2(n_861), .B1(n_879), .B2(n_881), .Y(n_878) );
INVx1_ASAP7_75t_L g1414 ( .A(n_856), .Y(n_1414) );
OAI22xp5_ASAP7_75t_L g889 ( .A1(n_857), .A2(n_863), .B1(n_874), .B2(n_890), .Y(n_889) );
OAI22xp5_ASAP7_75t_L g1370 ( .A1(n_858), .A2(n_1144), .B1(n_1371), .B2(n_1372), .Y(n_1370) );
OAI22xp5_ASAP7_75t_L g859 ( .A1(n_860), .A2(n_861), .B1(n_862), .B2(n_863), .Y(n_859) );
OAI221xp5_ASAP7_75t_L g1407 ( .A1(n_862), .A2(n_1408), .B1(n_1410), .B2(n_1411), .C(n_1412), .Y(n_1407) );
OAI221xp5_ASAP7_75t_L g1415 ( .A1(n_862), .A2(n_1416), .B1(n_1418), .B2(n_1419), .C(n_1420), .Y(n_1415) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
AOI33xp33_ASAP7_75t_L g1461 ( .A1(n_865), .A2(n_1096), .A3(n_1462), .B1(n_1466), .B2(n_1467), .B3(n_1469), .Y(n_1461) );
BUFx2_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
BUFx2_ASAP7_75t_L g1270 ( .A(n_866), .Y(n_1270) );
OAI33xp33_ASAP7_75t_L g1521 ( .A1(n_872), .A2(n_1330), .A3(n_1522), .B1(n_1525), .B2(n_1528), .B3(n_1531), .Y(n_1521) );
INVx2_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
HB1xp67_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx2_ASAP7_75t_L g891 ( .A(n_877), .Y(n_891) );
OAI22xp5_ASAP7_75t_L g1858 ( .A1(n_877), .A2(n_1859), .B1(n_1860), .B2(n_1861), .Y(n_1858) );
OAI221xp5_ASAP7_75t_L g1210 ( .A1(n_879), .A2(n_1204), .B1(n_1211), .B2(n_1212), .C(n_1213), .Y(n_1210) );
INVx2_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
BUFx2_ASAP7_75t_L g1322 ( .A(n_880), .Y(n_1322) );
INVx2_ASAP7_75t_L g1391 ( .A(n_880), .Y(n_1391) );
HB1xp67_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
OAI211xp5_ASAP7_75t_SL g1043 ( .A1(n_882), .A2(n_1044), .B(n_1045), .C(n_1046), .Y(n_1043) );
OAI22xp5_ASAP7_75t_L g1316 ( .A1(n_882), .A2(n_1317), .B1(n_1318), .B2(n_1319), .Y(n_1316) );
INVx2_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx2_ASAP7_75t_L g1167 ( .A(n_883), .Y(n_1167) );
INVx1_ASAP7_75t_L g1530 ( .A(n_883), .Y(n_1530) );
INVx2_ASAP7_75t_L g1840 ( .A(n_883), .Y(n_1840) );
OAI221xp5_ASAP7_75t_L g1165 ( .A1(n_885), .A2(n_1166), .B1(n_1167), .B2(n_1168), .C(n_1169), .Y(n_1165) );
INVx3_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx2_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
OAI221xp5_ASAP7_75t_L g1388 ( .A1(n_887), .A2(n_1212), .B1(n_1364), .B2(n_1371), .C(n_1389), .Y(n_1388) );
INVx2_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx2_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx2_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
OAI31xp33_ASAP7_75t_L g906 ( .A1(n_907), .A2(n_909), .A3(n_913), .B(n_917), .Y(n_906) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
BUFx2_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
XNOR2xp5_ASAP7_75t_L g921 ( .A(n_922), .B(n_1051), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
XNOR2xp5_ASAP7_75t_L g923 ( .A(n_924), .B(n_982), .Y(n_923) );
XOR2x2_ASAP7_75t_L g924 ( .A(n_925), .B(n_981), .Y(n_924) );
NOR2xp33_ASAP7_75t_L g925 ( .A(n_926), .B(n_960), .Y(n_925) );
INVx3_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
AOI22xp5_ASAP7_75t_L g934 ( .A1(n_935), .A2(n_936), .B1(n_938), .B2(n_939), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g1422 ( .A1(n_936), .A2(n_939), .B1(n_1423), .B2(n_1424), .Y(n_1422) );
INVx2_ASAP7_75t_L g1506 ( .A(n_936), .Y(n_1506) );
INVx1_ASAP7_75t_L g1507 ( .A(n_939), .Y(n_1507) );
OAI22xp5_ASAP7_75t_L g944 ( .A1(n_945), .A2(n_948), .B1(n_952), .B2(n_955), .Y(n_944) );
OAI22xp5_ASAP7_75t_L g1351 ( .A1(n_951), .A2(n_1109), .B1(n_1317), .B2(n_1329), .Y(n_1351) );
INVx1_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
NAND4xp25_ASAP7_75t_SL g960 ( .A(n_961), .B(n_962), .C(n_964), .D(n_967), .Y(n_960) );
BUFx3_ASAP7_75t_L g1796 ( .A(n_969), .Y(n_1796) );
HB1xp67_ASAP7_75t_L g1209 ( .A(n_972), .Y(n_1209) );
INVx2_ASAP7_75t_SL g972 ( .A(n_973), .Y(n_972) );
AND2x4_ASAP7_75t_L g977 ( .A(n_978), .B(n_979), .Y(n_977) );
NAND3xp33_ASAP7_75t_SL g983 ( .A(n_984), .B(n_992), .C(n_1018), .Y(n_983) );
AOI21xp33_ASAP7_75t_L g984 ( .A1(n_985), .A2(n_987), .B(n_988), .Y(n_984) );
AOI21xp5_ASAP7_75t_L g1084 ( .A1(n_985), .A2(n_1085), .B(n_1086), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1253 ( .A(n_985), .B(n_1254), .Y(n_1253) );
AOI221xp5_ASAP7_75t_L g1274 ( .A1(n_985), .A2(n_1264), .B1(n_1275), .B2(n_1276), .C(n_1277), .Y(n_1274) );
AOI221xp5_ASAP7_75t_L g1454 ( .A1(n_985), .A2(n_1264), .B1(n_1455), .B2(n_1456), .C(n_1457), .Y(n_1454) );
INVx8_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_990), .B(n_1179), .Y(n_1178) );
NOR3xp33_ASAP7_75t_L g992 ( .A(n_993), .B(n_1012), .C(n_1017), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_994), .B(n_1000), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_995), .A2(n_996), .B1(n_997), .B2(n_998), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g1285 ( .A1(n_996), .A2(n_998), .B1(n_1286), .B2(n_1287), .Y(n_1285) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_998), .A2(n_1092), .B1(n_1093), .B2(n_1094), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g1458 ( .A1(n_998), .A2(n_1258), .B1(n_1459), .B2(n_1460), .Y(n_1458) );
AOI33xp33_ASAP7_75t_L g1000 ( .A1(n_1001), .A2(n_1003), .A3(n_1004), .B1(n_1007), .B2(n_1009), .B3(n_1011), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_1002), .A2(n_1146), .B1(n_1147), .B2(n_1148), .Y(n_1145) );
HB1xp67_ASAP7_75t_L g1413 ( .A(n_1002), .Y(n_1413) );
BUFx3_ASAP7_75t_L g1096 ( .A(n_1003), .Y(n_1096) );
AOI33xp33_ASAP7_75t_L g1265 ( .A1(n_1003), .A2(n_1266), .A3(n_1267), .B1(n_1268), .B2(n_1269), .B3(n_1270), .Y(n_1265) );
AOI33xp33_ASAP7_75t_L g1278 ( .A1(n_1003), .A2(n_1009), .A3(n_1279), .B1(n_1282), .B2(n_1283), .B3(n_1284), .Y(n_1278) );
AOI33xp33_ASAP7_75t_L g1823 ( .A1(n_1003), .A2(n_1009), .A3(n_1824), .B1(n_1826), .B2(n_1827), .B3(n_1828), .Y(n_1823) );
INVx2_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
INVx2_ASAP7_75t_R g1008 ( .A(n_1006), .Y(n_1008) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1006), .Y(n_1110) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
INVx2_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g1830 ( .A(n_1016), .B(n_1831), .Y(n_1830) );
INVx3_ASAP7_75t_L g1115 ( .A(n_1017), .Y(n_1115) );
INVx3_ASAP7_75t_L g1271 ( .A(n_1017), .Y(n_1271) );
AOI221xp5_ASAP7_75t_L g1833 ( .A1(n_1017), .A2(n_1261), .B1(n_1834), .B2(n_1835), .C(n_1836), .Y(n_1833) );
OAI21xp5_ASAP7_75t_L g1018 ( .A1(n_1019), .A2(n_1034), .B(n_1047), .Y(n_1018) );
INVx2_ASAP7_75t_SL g1020 ( .A(n_1021), .Y(n_1020) );
INVx3_ASAP7_75t_L g1056 ( .A(n_1021), .Y(n_1056) );
AOI221xp5_ASAP7_75t_L g1294 ( .A1(n_1021), .A2(n_1028), .B1(n_1275), .B2(n_1295), .C(n_1296), .Y(n_1294) );
AOI221xp5_ASAP7_75t_L g1476 ( .A1(n_1021), .A2(n_1028), .B1(n_1455), .B2(n_1477), .C(n_1481), .Y(n_1476) );
AOI21xp5_ASAP7_75t_L g1022 ( .A1(n_1023), .A2(n_1025), .B(n_1028), .Y(n_1022) );
AOI21xp5_ASAP7_75t_L g1057 ( .A1(n_1028), .A2(n_1058), .B(n_1066), .Y(n_1057) );
AOI21xp5_ASAP7_75t_L g1240 ( .A1(n_1028), .A2(n_1241), .B(n_1244), .Y(n_1240) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_1030), .A2(n_1031), .B1(n_1032), .B2(n_1033), .Y(n_1029) );
HB1xp67_ASAP7_75t_L g1070 ( .A(n_1031), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1245 ( .A1(n_1031), .A2(n_1033), .B1(n_1246), .B2(n_1247), .Y(n_1245) );
AOI22xp33_ASAP7_75t_L g1298 ( .A1(n_1031), .A2(n_1033), .B1(n_1299), .B2(n_1300), .Y(n_1298) );
AOI22xp33_ASAP7_75t_L g1472 ( .A1(n_1031), .A2(n_1473), .B1(n_1474), .B2(n_1475), .Y(n_1472) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1033), .Y(n_1073) );
BUFx6f_ASAP7_75t_L g1475 ( .A(n_1033), .Y(n_1475) );
INVx1_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
INVx2_ASAP7_75t_L g1075 ( .A(n_1036), .Y(n_1075) );
INVx2_ASAP7_75t_L g1230 ( .A(n_1036), .Y(n_1230) );
INVx4_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
INVx2_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
BUFx3_ASAP7_75t_L g1291 ( .A(n_1038), .Y(n_1291) );
BUFx2_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
INVx2_ASAP7_75t_L g1040 ( .A(n_1041), .Y(n_1040) );
AOI21xp5_ASAP7_75t_L g1288 ( .A1(n_1047), .A2(n_1289), .B(n_1301), .Y(n_1288) );
INVx1_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
OAI21xp33_ASAP7_75t_L g1182 ( .A1(n_1048), .A2(n_1183), .B(n_1196), .Y(n_1182) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1049), .Y(n_1048) );
BUFx2_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
BUFx2_ASAP7_75t_L g1083 ( .A(n_1050), .Y(n_1083) );
HB1xp67_ASAP7_75t_L g1380 ( .A(n_1050), .Y(n_1380) );
OAI31xp33_ASAP7_75t_L g1837 ( .A1(n_1050), .A2(n_1838), .A3(n_1843), .B(n_1855), .Y(n_1837) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
NAND3xp33_ASAP7_75t_SL g1053 ( .A(n_1054), .B(n_1084), .C(n_1089), .Y(n_1053) );
OAI21xp33_ASAP7_75t_L g1054 ( .A1(n_1055), .A2(n_1074), .B(n_1083), .Y(n_1054) );
BUFx2_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
BUFx2_ASAP7_75t_L g1803 ( .A(n_1063), .Y(n_1803) );
AOI221xp5_ASAP7_75t_L g1845 ( .A1(n_1063), .A2(n_1831), .B1(n_1836), .B2(n_1846), .C(n_1848), .Y(n_1845) );
HB1xp67_ASAP7_75t_SL g1064 ( .A(n_1065), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_1069), .A2(n_1070), .B1(n_1071), .B2(n_1072), .Y(n_1068) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
OAI221xp5_ASAP7_75t_L g1076 ( .A1(n_1077), .A2(n_1078), .B1(n_1079), .B2(n_1080), .C(n_1081), .Y(n_1076) );
OAI22xp5_ASAP7_75t_SL g1435 ( .A1(n_1077), .A2(n_1410), .B1(n_1436), .B2(n_1437), .Y(n_1435) );
INVx3_ASAP7_75t_L g1264 ( .A(n_1088), .Y(n_1264) );
INVx5_ASAP7_75t_L g1864 ( .A(n_1088), .Y(n_1864) );
NOR3xp33_ASAP7_75t_L g1089 ( .A(n_1090), .B(n_1112), .C(n_1114), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_1091), .B(n_1095), .Y(n_1090) );
BUFx2_ASAP7_75t_SL g1098 ( .A(n_1099), .Y(n_1098) );
INVx2_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
INVx2_ASAP7_75t_SL g1100 ( .A(n_1101), .Y(n_1100) );
NAND2xp5_ASAP7_75t_L g1377 ( .A(n_1101), .B(n_1378), .Y(n_1377) );
BUFx3_ASAP7_75t_L g1421 ( .A(n_1101), .Y(n_1421) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1101), .Y(n_1464) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
INVx2_ASAP7_75t_SL g1114 ( .A(n_1115), .Y(n_1114) );
NAND3xp33_ASAP7_75t_SL g1457 ( .A(n_1115), .B(n_1458), .C(n_1461), .Y(n_1457) );
AOI22xp5_ASAP7_75t_L g1116 ( .A1(n_1117), .A2(n_1118), .B1(n_1394), .B2(n_1395), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1118), .Y(n_1117) );
HB1xp67_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
XNOR2x1_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1223), .Y(n_1119) );
XNOR2x2_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1173), .Y(n_1120) );
AOI21xp5_ASAP7_75t_L g1121 ( .A1(n_1122), .A2(n_1171), .B(n_1172), .Y(n_1121) );
AND3x1_ASAP7_75t_L g1122 ( .A(n_1123), .B(n_1152), .C(n_1158), .Y(n_1122) );
AOI31xp33_ASAP7_75t_L g1172 ( .A1(n_1123), .A2(n_1152), .A3(n_1158), .B(n_1171), .Y(n_1172) );
AOI21xp5_ASAP7_75t_L g1123 ( .A1(n_1124), .A2(n_1150), .B(n_1151), .Y(n_1123) );
NAND3xp33_ASAP7_75t_SL g1124 ( .A(n_1125), .B(n_1137), .C(n_1140), .Y(n_1124) );
AOI22xp5_ASAP7_75t_L g1125 ( .A1(n_1126), .A2(n_1128), .B1(n_1131), .B2(n_1134), .Y(n_1125) );
INVx2_ASAP7_75t_L g1132 ( .A(n_1133), .Y(n_1132) );
BUFx2_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1136), .Y(n_1347) );
INVxp67_ASAP7_75t_L g1184 ( .A(n_1141), .Y(n_1184) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1150), .Y(n_1248) );
INVx2_ASAP7_75t_L g1352 ( .A(n_1150), .Y(n_1352) );
OAI31xp33_ASAP7_75t_SL g1400 ( .A1(n_1150), .A2(n_1401), .A3(n_1402), .B(n_1406), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1153), .B(n_1155), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_1156), .B(n_1157), .Y(n_1155) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
NAND3xp33_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1182), .C(n_1206), .Y(n_1175) );
OAI211xp5_ASAP7_75t_L g1183 ( .A1(n_1184), .A2(n_1185), .B(n_1187), .C(n_1190), .Y(n_1183) );
OAI211xp5_ASAP7_75t_L g1190 ( .A1(n_1191), .A2(n_1192), .B(n_1194), .C(n_1195), .Y(n_1190) );
HB1xp67_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
NOR3xp33_ASAP7_75t_L g1206 ( .A(n_1207), .B(n_1214), .C(n_1218), .Y(n_1206) );
INVxp67_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
XNOR2xp5_ASAP7_75t_L g1223 ( .A(n_1224), .B(n_1303), .Y(n_1223) );
XNOR2xp5_ASAP7_75t_L g1224 ( .A(n_1225), .B(n_1272), .Y(n_1224) );
NOR2x1p5_ASAP7_75t_L g1226 ( .A(n_1227), .B(n_1252), .Y(n_1226) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
O2A1O1Ixp33_ASAP7_75t_SL g1228 ( .A1(n_1229), .A2(n_1239), .B(n_1248), .C(n_1249), .Y(n_1228) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
AOI21xp5_ASAP7_75t_SL g1470 ( .A1(n_1248), .A2(n_1471), .B(n_1488), .Y(n_1470) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_1253), .B(n_1255), .Y(n_1252) );
AND4x1_ASAP7_75t_L g1255 ( .A(n_1256), .B(n_1262), .C(n_1265), .D(n_1271), .Y(n_1255) );
AOI22xp5_ASAP7_75t_L g1256 ( .A1(n_1257), .A2(n_1258), .B1(n_1260), .B2(n_1261), .Y(n_1256) );
INVx2_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
NAND2xp5_ASAP7_75t_L g1262 ( .A(n_1263), .B(n_1264), .Y(n_1262) );
NAND3xp33_ASAP7_75t_L g1277 ( .A(n_1271), .B(n_1278), .C(n_1285), .Y(n_1277) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1274), .B(n_1288), .Y(n_1273) );
NAND3xp33_ASAP7_75t_L g1289 ( .A(n_1290), .B(n_1294), .C(n_1298), .Y(n_1289) );
AOI222xp33_ASAP7_75t_L g1482 ( .A1(n_1291), .A2(n_1459), .B1(n_1460), .B2(n_1483), .C1(n_1485), .C2(n_1486), .Y(n_1482) );
XNOR2x1_ASAP7_75t_L g1303 ( .A(n_1304), .B(n_1355), .Y(n_1303) );
XNOR2x1_ASAP7_75t_L g1304 ( .A(n_1305), .B(n_1306), .Y(n_1304) );
NOR2x1_ASAP7_75t_L g1306 ( .A(n_1307), .B(n_1339), .Y(n_1306) );
NAND3xp33_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1333), .C(n_1337), .Y(n_1307) );
NOR2xp33_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1332), .Y(n_1308) );
OAI33xp33_ASAP7_75t_L g1309 ( .A1(n_1310), .A2(n_1311), .A3(n_1316), .B1(n_1320), .B2(n_1325), .B3(n_1330), .Y(n_1309) );
OAI22xp5_ASAP7_75t_L g1311 ( .A1(n_1312), .A2(n_1313), .B1(n_1314), .B2(n_1315), .Y(n_1311) );
OAI22xp5_ASAP7_75t_L g1325 ( .A1(n_1315), .A2(n_1326), .B1(n_1328), .B2(n_1329), .Y(n_1325) );
HB1xp67_ASAP7_75t_L g1437 ( .A(n_1315), .Y(n_1437) );
OAI22xp5_ASAP7_75t_L g1531 ( .A1(n_1315), .A2(n_1504), .B1(n_1532), .B2(n_1533), .Y(n_1531) );
OAI22xp5_ASAP7_75t_L g1528 ( .A1(n_1321), .A2(n_1510), .B1(n_1529), .B2(n_1530), .Y(n_1528) );
INVx4_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1327), .Y(n_1326) );
INVx2_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
A2O1A1Ixp33_ASAP7_75t_L g1339 ( .A1(n_1340), .A2(n_1344), .B(n_1352), .C(n_1353), .Y(n_1339) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1347), .Y(n_1346) );
INVx1_ASAP7_75t_L g1512 ( .A(n_1352), .Y(n_1512) );
INVx2_ASAP7_75t_L g1355 ( .A(n_1356), .Y(n_1355) );
XNOR2x1_ASAP7_75t_L g1356 ( .A(n_1357), .B(n_1358), .Y(n_1356) );
OR2x2_ASAP7_75t_L g1358 ( .A(n_1359), .B(n_1382), .Y(n_1358) );
A2O1A1Ixp33_ASAP7_75t_L g1359 ( .A1(n_1360), .A2(n_1373), .B(n_1380), .C(n_1381), .Y(n_1359) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
OA22x2_ASAP7_75t_L g1395 ( .A1(n_1396), .A2(n_1450), .B1(n_1451), .B2(n_1534), .Y(n_1395) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1396), .Y(n_1534) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1398), .Y(n_1397) );
NOR2x1_ASAP7_75t_L g1398 ( .A(n_1399), .B(n_1425), .Y(n_1398) );
NAND3xp33_ASAP7_75t_L g1406 ( .A(n_1407), .B(n_1415), .C(n_1422), .Y(n_1406) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
NAND2xp5_ASAP7_75t_L g1425 ( .A(n_1426), .B(n_1439), .Y(n_1425) );
INVx1_ASAP7_75t_SL g1430 ( .A(n_1431), .Y(n_1430) );
AOI21xp5_ASAP7_75t_L g1439 ( .A1(n_1440), .A2(n_1441), .B(n_1443), .Y(n_1439) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1442), .Y(n_1441) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1451), .Y(n_1450) );
XNOR2xp5_ASAP7_75t_L g1451 ( .A(n_1452), .B(n_1490), .Y(n_1451) );
NAND2xp5_ASAP7_75t_L g1453 ( .A(n_1454), .B(n_1470), .Y(n_1453) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
NAND3xp33_ASAP7_75t_SL g1471 ( .A(n_1472), .B(n_1476), .C(n_1482), .Y(n_1471) );
INVx2_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1487), .Y(n_1486) );
AOI211x1_ASAP7_75t_L g1491 ( .A1(n_1492), .A2(n_1512), .B(n_1513), .C(n_1519), .Y(n_1491) );
NAND2xp5_ASAP7_75t_L g1492 ( .A(n_1493), .B(n_1497), .Y(n_1492) );
NOR3xp33_ASAP7_75t_L g1497 ( .A(n_1498), .B(n_1505), .C(n_1508), .Y(n_1497) );
OAI22xp5_ASAP7_75t_L g1525 ( .A1(n_1502), .A2(n_1511), .B1(n_1526), .B2(n_1527), .Y(n_1525) );
OAI22xp5_ASAP7_75t_L g1804 ( .A1(n_1527), .A2(n_1532), .B1(n_1774), .B2(n_1805), .Y(n_1804) );
OAI221xp5_ASAP7_75t_L g1535 ( .A1(n_1536), .A2(n_1755), .B1(n_1759), .B2(n_1806), .C(n_1810), .Y(n_1535) );
AOI211xp5_ASAP7_75t_L g1536 ( .A1(n_1537), .A2(n_1660), .B(n_1667), .C(n_1733), .Y(n_1536) );
NAND5xp2_ASAP7_75t_L g1537 ( .A(n_1538), .B(n_1611), .C(n_1638), .D(n_1641), .E(n_1646), .Y(n_1537) );
AOI211xp5_ASAP7_75t_L g1538 ( .A1(n_1539), .A2(n_1569), .B(n_1578), .C(n_1606), .Y(n_1538) );
INVx1_ASAP7_75t_L g1539 ( .A(n_1540), .Y(n_1539) );
OR2x2_ASAP7_75t_L g1540 ( .A(n_1541), .B(n_1556), .Y(n_1540) );
OAI321xp33_ASAP7_75t_L g1578 ( .A1(n_1541), .A2(n_1579), .A3(n_1586), .B1(n_1591), .B2(n_1592), .C(n_1597), .Y(n_1578) );
AND2x2_ASAP7_75t_L g1599 ( .A(n_1541), .B(n_1557), .Y(n_1599) );
AND3x1_ASAP7_75t_L g1632 ( .A(n_1541), .B(n_1566), .C(n_1590), .Y(n_1632) );
AND2x2_ASAP7_75t_L g1637 ( .A(n_1541), .B(n_1624), .Y(n_1637) );
NAND2xp5_ASAP7_75t_L g1657 ( .A(n_1541), .B(n_1566), .Y(n_1657) );
OR2x2_ASAP7_75t_L g1684 ( .A(n_1541), .B(n_1685), .Y(n_1684) );
AND2x2_ASAP7_75t_L g1687 ( .A(n_1541), .B(n_1587), .Y(n_1687) );
NAND2xp5_ASAP7_75t_L g1726 ( .A(n_1541), .B(n_1590), .Y(n_1726) );
INVx2_ASAP7_75t_L g1541 ( .A(n_1542), .Y(n_1541) );
AND2x2_ASAP7_75t_L g1596 ( .A(n_1542), .B(n_1587), .Y(n_1596) );
BUFx2_ASAP7_75t_L g1602 ( .A(n_1542), .Y(n_1602) );
OR2x2_ASAP7_75t_L g1693 ( .A(n_1542), .B(n_1679), .Y(n_1693) );
AND2x2_ASAP7_75t_L g1705 ( .A(n_1542), .B(n_1624), .Y(n_1705) );
AND2x2_ASAP7_75t_L g1542 ( .A(n_1543), .B(n_1551), .Y(n_1542) );
AND2x4_ASAP7_75t_L g1544 ( .A(n_1545), .B(n_1546), .Y(n_1544) );
AND2x6_ASAP7_75t_L g1549 ( .A(n_1545), .B(n_1550), .Y(n_1549) );
AND2x6_ASAP7_75t_L g1552 ( .A(n_1545), .B(n_1553), .Y(n_1552) );
AND2x2_ASAP7_75t_L g1554 ( .A(n_1545), .B(n_1555), .Y(n_1554) );
AND2x2_ASAP7_75t_L g1561 ( .A(n_1545), .B(n_1555), .Y(n_1561) );
AND2x2_ASAP7_75t_L g1573 ( .A(n_1545), .B(n_1555), .Y(n_1573) );
AND2x2_ASAP7_75t_L g1546 ( .A(n_1547), .B(n_1548), .Y(n_1546) );
INVx2_ASAP7_75t_L g1664 ( .A(n_1552), .Y(n_1664) );
OAI21xp5_ASAP7_75t_L g1868 ( .A1(n_1555), .A2(n_1869), .B(n_1870), .Y(n_1868) );
NAND2xp5_ASAP7_75t_L g1556 ( .A(n_1557), .B(n_1562), .Y(n_1556) );
AND2x2_ASAP7_75t_L g1580 ( .A(n_1557), .B(n_1581), .Y(n_1580) );
NOR2xp33_ASAP7_75t_L g1614 ( .A(n_1557), .B(n_1615), .Y(n_1614) );
INVx1_ASAP7_75t_L g1649 ( .A(n_1557), .Y(n_1649) );
NAND2xp5_ASAP7_75t_L g1675 ( .A(n_1557), .B(n_1619), .Y(n_1675) );
NOR2xp33_ASAP7_75t_L g1709 ( .A(n_1557), .B(n_1710), .Y(n_1709) );
NAND2xp5_ASAP7_75t_L g1744 ( .A(n_1557), .B(n_1587), .Y(n_1744) );
INVx2_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
INVx1_ASAP7_75t_L g1595 ( .A(n_1558), .Y(n_1595) );
AND2x2_ASAP7_75t_L g1601 ( .A(n_1558), .B(n_1602), .Y(n_1601) );
AND2x2_ASAP7_75t_L g1630 ( .A(n_1558), .B(n_1571), .Y(n_1630) );
NAND2xp5_ASAP7_75t_L g1679 ( .A(n_1558), .B(n_1562), .Y(n_1679) );
NOR2xp33_ASAP7_75t_L g1681 ( .A(n_1558), .B(n_1682), .Y(n_1681) );
AND2x2_ASAP7_75t_L g1725 ( .A(n_1558), .B(n_1582), .Y(n_1725) );
AND2x2_ASAP7_75t_L g1558 ( .A(n_1559), .B(n_1560), .Y(n_1558) );
INVxp67_ASAP7_75t_L g1666 ( .A(n_1561), .Y(n_1666) );
HB1xp67_ASAP7_75t_L g1758 ( .A(n_1561), .Y(n_1758) );
AND2x2_ASAP7_75t_L g1695 ( .A(n_1562), .B(n_1601), .Y(n_1695) );
AND2x2_ASAP7_75t_L g1562 ( .A(n_1563), .B(n_1566), .Y(n_1562) );
AND2x2_ASAP7_75t_L g1587 ( .A(n_1563), .B(n_1588), .Y(n_1587) );
INVx2_ASAP7_75t_L g1590 ( .A(n_1563), .Y(n_1590) );
NAND2xp5_ASAP7_75t_L g1615 ( .A(n_1563), .B(n_1602), .Y(n_1615) );
NAND3xp33_ASAP7_75t_L g1688 ( .A(n_1563), .B(n_1593), .C(n_1661), .Y(n_1688) );
OR2x2_ASAP7_75t_L g1563 ( .A(n_1564), .B(n_1565), .Y(n_1563) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1566), .Y(n_1588) );
AND2x2_ASAP7_75t_L g1589 ( .A(n_1566), .B(n_1590), .Y(n_1589) );
AND2x2_ASAP7_75t_L g1674 ( .A(n_1566), .B(n_1602), .Y(n_1674) );
OR2x2_ASAP7_75t_L g1710 ( .A(n_1566), .B(n_1602), .Y(n_1710) );
AND2x2_ASAP7_75t_L g1566 ( .A(n_1567), .B(n_1568), .Y(n_1566) );
A2O1A1Ixp33_ASAP7_75t_L g1677 ( .A1(n_1569), .A2(n_1661), .B(n_1678), .C(n_1680), .Y(n_1677) );
INVx1_ASAP7_75t_L g1569 ( .A(n_1570), .Y(n_1569) );
OR2x2_ASAP7_75t_L g1570 ( .A(n_1571), .B(n_1575), .Y(n_1570) );
CKINVDCx6p67_ASAP7_75t_R g1604 ( .A(n_1571), .Y(n_1604) );
OR2x2_ASAP7_75t_L g1608 ( .A(n_1571), .B(n_1609), .Y(n_1608) );
NAND2xp5_ASAP7_75t_L g1651 ( .A(n_1571), .B(n_1619), .Y(n_1651) );
AND2x2_ASAP7_75t_L g1659 ( .A(n_1571), .B(n_1575), .Y(n_1659) );
NAND2xp5_ASAP7_75t_L g1741 ( .A(n_1571), .B(n_1661), .Y(n_1741) );
NAND2xp5_ASAP7_75t_L g1748 ( .A(n_1571), .B(n_1749), .Y(n_1748) );
OR2x6_ASAP7_75t_L g1571 ( .A(n_1572), .B(n_1574), .Y(n_1571) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1575), .Y(n_1585) );
INVx3_ASAP7_75t_L g1591 ( .A(n_1575), .Y(n_1591) );
AND2x2_ASAP7_75t_L g1610 ( .A(n_1575), .B(n_1605), .Y(n_1610) );
OR2x2_ASAP7_75t_L g1613 ( .A(n_1575), .B(n_1582), .Y(n_1613) );
AND2x2_ASAP7_75t_L g1625 ( .A(n_1575), .B(n_1604), .Y(n_1625) );
AND2x2_ASAP7_75t_L g1628 ( .A(n_1575), .B(n_1582), .Y(n_1628) );
OR2x2_ASAP7_75t_L g1643 ( .A(n_1575), .B(n_1604), .Y(n_1643) );
OAI221xp5_ASAP7_75t_L g1702 ( .A1(n_1575), .A2(n_1703), .B1(n_1704), .B2(n_1706), .C(n_1707), .Y(n_1702) );
OAI32xp33_ASAP7_75t_L g1729 ( .A1(n_1575), .A2(n_1591), .A3(n_1593), .B1(n_1684), .B2(n_1730), .Y(n_1729) );
AND2x4_ASAP7_75t_L g1575 ( .A(n_1576), .B(n_1577), .Y(n_1575) );
OAI32xp33_ASAP7_75t_L g1746 ( .A1(n_1579), .A2(n_1593), .A3(n_1633), .B1(n_1747), .B2(n_1748), .Y(n_1746) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
INVx1_ASAP7_75t_L g1633 ( .A(n_1581), .Y(n_1633) );
AND2x2_ASAP7_75t_L g1690 ( .A(n_1581), .B(n_1604), .Y(n_1690) );
AND2x2_ASAP7_75t_L g1581 ( .A(n_1582), .B(n_1585), .Y(n_1581) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1582), .Y(n_1605) );
AND2x2_ASAP7_75t_L g1582 ( .A(n_1583), .B(n_1584), .Y(n_1582) );
OR2x2_ASAP7_75t_L g1586 ( .A(n_1587), .B(n_1589), .Y(n_1586) );
AND2x2_ASAP7_75t_L g1600 ( .A(n_1587), .B(n_1601), .Y(n_1600) );
AND2x2_ASAP7_75t_L g1624 ( .A(n_1588), .B(n_1590), .Y(n_1624) );
O2A1O1Ixp33_ASAP7_75t_L g1697 ( .A1(n_1588), .A2(n_1698), .B(n_1699), .C(n_1700), .Y(n_1697) );
AND2x2_ASAP7_75t_L g1598 ( .A(n_1589), .B(n_1599), .Y(n_1598) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1589), .Y(n_1607) );
AND2x2_ASAP7_75t_L g1645 ( .A(n_1589), .B(n_1602), .Y(n_1645) );
OAI322xp33_ASAP7_75t_L g1626 ( .A1(n_1590), .A2(n_1627), .A3(n_1629), .B1(n_1631), .B2(n_1633), .C1(n_1634), .C2(n_1636), .Y(n_1626) );
OR2x2_ASAP7_75t_L g1682 ( .A(n_1590), .B(n_1602), .Y(n_1682) );
AND2x2_ASAP7_75t_L g1731 ( .A(n_1590), .B(n_1602), .Y(n_1731) );
CKINVDCx14_ASAP7_75t_R g1722 ( .A(n_1591), .Y(n_1722) );
NAND2xp5_ASAP7_75t_L g1592 ( .A(n_1593), .B(n_1596), .Y(n_1592) );
NAND2xp5_ASAP7_75t_L g1719 ( .A(n_1593), .B(n_1687), .Y(n_1719) );
INVx1_ASAP7_75t_L g1593 ( .A(n_1594), .Y(n_1593) );
NAND2xp5_ASAP7_75t_L g1640 ( .A(n_1594), .B(n_1637), .Y(n_1640) );
NAND2xp5_ASAP7_75t_L g1698 ( .A(n_1594), .B(n_1635), .Y(n_1698) );
AND2x2_ASAP7_75t_L g1716 ( .A(n_1594), .B(n_1687), .Y(n_1716) );
INVx2_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
AND2x2_ASAP7_75t_L g1644 ( .A(n_1595), .B(n_1645), .Y(n_1644) );
NAND2xp5_ASAP7_75t_L g1685 ( .A(n_1595), .B(n_1624), .Y(n_1685) );
AND2x2_ASAP7_75t_L g1735 ( .A(n_1595), .B(n_1635), .Y(n_1735) );
AND2x2_ASAP7_75t_L g1752 ( .A(n_1596), .B(n_1619), .Y(n_1752) );
OAI21xp5_ASAP7_75t_L g1597 ( .A1(n_1598), .A2(n_1600), .B(n_1603), .Y(n_1597) );
INVx1_ASAP7_75t_L g1676 ( .A(n_1598), .Y(n_1676) );
AND2x2_ASAP7_75t_L g1654 ( .A(n_1599), .B(n_1624), .Y(n_1654) );
INVx1_ASAP7_75t_L g1739 ( .A(n_1600), .Y(n_1739) );
INVx1_ASAP7_75t_L g1622 ( .A(n_1601), .Y(n_1622) );
INVx1_ASAP7_75t_L g1692 ( .A(n_1603), .Y(n_1692) );
NAND2xp5_ASAP7_75t_L g1704 ( .A(n_1603), .B(n_1705), .Y(n_1704) );
AND2x2_ASAP7_75t_L g1603 ( .A(n_1604), .B(n_1605), .Y(n_1603) );
NOR2xp33_ASAP7_75t_L g1612 ( .A(n_1604), .B(n_1613), .Y(n_1612) );
NAND2xp5_ASAP7_75t_L g1634 ( .A(n_1604), .B(n_1635), .Y(n_1634) );
NOR2xp33_ASAP7_75t_SL g1696 ( .A(n_1604), .B(n_1633), .Y(n_1696) );
NAND2xp5_ASAP7_75t_L g1700 ( .A(n_1604), .B(n_1661), .Y(n_1700) );
AND2x2_ASAP7_75t_L g1714 ( .A(n_1604), .B(n_1619), .Y(n_1714) );
INVx2_ASAP7_75t_L g1619 ( .A(n_1605), .Y(n_1619) );
NOR2xp33_ASAP7_75t_L g1606 ( .A(n_1607), .B(n_1608), .Y(n_1606) );
INVx1_ASAP7_75t_L g1745 ( .A(n_1608), .Y(n_1745) );
OAI22xp5_ASAP7_75t_L g1712 ( .A1(n_1609), .A2(n_1684), .B1(n_1713), .B2(n_1715), .Y(n_1712) );
OAI211xp5_ASAP7_75t_L g1720 ( .A1(n_1609), .A2(n_1686), .B(n_1721), .C(n_1727), .Y(n_1720) );
CKINVDCx6p67_ASAP7_75t_R g1609 ( .A(n_1610), .Y(n_1609) );
NAND2xp5_ASAP7_75t_L g1648 ( .A(n_1610), .B(n_1649), .Y(n_1648) );
AOI221xp5_ASAP7_75t_L g1611 ( .A1(n_1612), .A2(n_1614), .B1(n_1616), .B2(n_1625), .C(n_1626), .Y(n_1611) );
INVx2_ASAP7_75t_L g1635 ( .A(n_1613), .Y(n_1635) );
AND2x2_ASAP7_75t_L g1616 ( .A(n_1617), .B(n_1620), .Y(n_1616) );
AND2x2_ASAP7_75t_L g1708 ( .A(n_1617), .B(n_1709), .Y(n_1708) );
A2O1A1Ixp33_ASAP7_75t_L g1736 ( .A1(n_1617), .A2(n_1685), .B(n_1686), .C(n_1737), .Y(n_1736) );
INVx2_ASAP7_75t_L g1617 ( .A(n_1618), .Y(n_1617) );
NAND2xp5_ASAP7_75t_L g1638 ( .A(n_1618), .B(n_1639), .Y(n_1638) );
NAND2xp5_ASAP7_75t_L g1658 ( .A(n_1618), .B(n_1659), .Y(n_1658) );
NOR2xp33_ASAP7_75t_L g1738 ( .A(n_1618), .B(n_1739), .Y(n_1738) );
NAND2xp5_ASAP7_75t_L g1754 ( .A(n_1618), .B(n_1716), .Y(n_1754) );
INVx2_ASAP7_75t_L g1618 ( .A(n_1619), .Y(n_1618) );
OR2x2_ASAP7_75t_L g1703 ( .A(n_1619), .B(n_1621), .Y(n_1703) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1621), .Y(n_1620) );
OR2x2_ASAP7_75t_L g1621 ( .A(n_1622), .B(n_1623), .Y(n_1621) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
INVx1_ASAP7_75t_L g1670 ( .A(n_1625), .Y(n_1670) );
AND2x2_ASAP7_75t_L g1680 ( .A(n_1625), .B(n_1681), .Y(n_1680) );
OAI22xp5_ASAP7_75t_L g1652 ( .A1(n_1627), .A2(n_1653), .B1(n_1655), .B2(n_1658), .Y(n_1652) );
NOR2xp33_ASAP7_75t_L g1728 ( .A(n_1627), .B(n_1631), .Y(n_1728) );
INVx2_ASAP7_75t_L g1627 ( .A(n_1628), .Y(n_1627) );
AOI22xp33_ASAP7_75t_L g1694 ( .A1(n_1628), .A2(n_1632), .B1(n_1695), .B2(n_1696), .Y(n_1694) );
CKINVDCx14_ASAP7_75t_R g1629 ( .A(n_1630), .Y(n_1629) );
INVx2_ASAP7_75t_L g1631 ( .A(n_1632), .Y(n_1631) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1637), .Y(n_1636) );
O2A1O1Ixp33_ASAP7_75t_L g1742 ( .A1(n_1639), .A2(n_1743), .B(n_1745), .C(n_1746), .Y(n_1742) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1640), .Y(n_1639) );
NAND2xp5_ASAP7_75t_L g1641 ( .A(n_1642), .B(n_1644), .Y(n_1641) );
INVx1_ASAP7_75t_L g1642 ( .A(n_1643), .Y(n_1642) );
O2A1O1Ixp33_ASAP7_75t_L g1646 ( .A1(n_1645), .A2(n_1647), .B(n_1650), .C(n_1652), .Y(n_1646) );
NOR2xp33_ASAP7_75t_L g1747 ( .A(n_1645), .B(n_1687), .Y(n_1747) );
INVx1_ASAP7_75t_L g1647 ( .A(n_1648), .Y(n_1647) );
NOR2xp33_ASAP7_75t_L g1656 ( .A(n_1649), .B(n_1657), .Y(n_1656) );
INVx1_ASAP7_75t_L g1650 ( .A(n_1651), .Y(n_1650) );
OAI221xp5_ASAP7_75t_L g1669 ( .A1(n_1651), .A2(n_1670), .B1(n_1671), .B2(n_1676), .C(n_1677), .Y(n_1669) );
INVx1_ASAP7_75t_L g1653 ( .A(n_1654), .Y(n_1653) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
OAI31xp33_ASAP7_75t_L g1750 ( .A1(n_1659), .A2(n_1751), .A3(n_1752), .B(n_1753), .Y(n_1750) );
INVx2_ASAP7_75t_SL g1660 ( .A(n_1661), .Y(n_1660) );
INVx2_ASAP7_75t_SL g1706 ( .A(n_1661), .Y(n_1706) );
OAI22xp5_ASAP7_75t_SL g1662 ( .A1(n_1663), .A2(n_1664), .B1(n_1665), .B2(n_1666), .Y(n_1662) );
NAND3xp33_ASAP7_75t_L g1667 ( .A(n_1668), .B(n_1701), .C(n_1717), .Y(n_1667) );
NOR4xp25_ASAP7_75t_L g1668 ( .A(n_1669), .B(n_1683), .C(n_1691), .D(n_1697), .Y(n_1668) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1672), .Y(n_1671) );
OAI21xp5_ASAP7_75t_L g1707 ( .A1(n_1672), .A2(n_1708), .B(n_1711), .Y(n_1707) );
NOR2xp33_ASAP7_75t_L g1672 ( .A(n_1673), .B(n_1675), .Y(n_1672) );
A2O1A1Ixp33_ASAP7_75t_L g1734 ( .A1(n_1673), .A2(n_1735), .B(n_1736), .C(n_1740), .Y(n_1734) );
INVx1_ASAP7_75t_L g1673 ( .A(n_1674), .Y(n_1673) );
INVx1_ASAP7_75t_L g1678 ( .A(n_1679), .Y(n_1678) );
AOI31xp33_ASAP7_75t_L g1683 ( .A1(n_1684), .A2(n_1686), .A3(n_1688), .B(n_1689), .Y(n_1683) );
INVx1_ASAP7_75t_L g1751 ( .A(n_1684), .Y(n_1751) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1687), .Y(n_1686) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1690), .Y(n_1689) );
OAI21xp33_ASAP7_75t_L g1691 ( .A1(n_1692), .A2(n_1693), .B(n_1694), .Y(n_1691) );
INVx1_ASAP7_75t_L g1699 ( .A(n_1695), .Y(n_1699) );
INVx1_ASAP7_75t_L g1711 ( .A(n_1700), .Y(n_1711) );
NOR2xp33_ASAP7_75t_L g1701 ( .A(n_1702), .B(n_1712), .Y(n_1701) );
INVx3_ASAP7_75t_L g1732 ( .A(n_1706), .Y(n_1732) );
INVx1_ASAP7_75t_L g1713 ( .A(n_1714), .Y(n_1713) );
INVx1_ASAP7_75t_L g1715 ( .A(n_1716), .Y(n_1715) );
OAI31xp33_ASAP7_75t_L g1717 ( .A1(n_1718), .A2(n_1720), .A3(n_1729), .B(n_1732), .Y(n_1717) );
INVx1_ASAP7_75t_L g1718 ( .A(n_1719), .Y(n_1718) );
NAND2xp5_ASAP7_75t_L g1721 ( .A(n_1722), .B(n_1723), .Y(n_1721) );
NOR2xp33_ASAP7_75t_L g1723 ( .A(n_1724), .B(n_1726), .Y(n_1723) );
CKINVDCx14_ASAP7_75t_R g1724 ( .A(n_1725), .Y(n_1724) );
INVx1_ASAP7_75t_L g1749 ( .A(n_1726), .Y(n_1749) );
INVx1_ASAP7_75t_L g1727 ( .A(n_1728), .Y(n_1727) );
CKINVDCx14_ASAP7_75t_R g1730 ( .A(n_1731), .Y(n_1730) );
NAND3xp33_ASAP7_75t_L g1733 ( .A(n_1734), .B(n_1742), .C(n_1750), .Y(n_1733) );
INVxp67_ASAP7_75t_L g1737 ( .A(n_1738), .Y(n_1737) );
INVx1_ASAP7_75t_L g1740 ( .A(n_1741), .Y(n_1740) );
INVx1_ASAP7_75t_L g1743 ( .A(n_1744), .Y(n_1743) );
INVx1_ASAP7_75t_L g1753 ( .A(n_1754), .Y(n_1753) );
CKINVDCx20_ASAP7_75t_R g1755 ( .A(n_1756), .Y(n_1755) );
CKINVDCx20_ASAP7_75t_R g1756 ( .A(n_1757), .Y(n_1756) );
INVx4_ASAP7_75t_L g1757 ( .A(n_1758), .Y(n_1757) );
HB1xp67_ASAP7_75t_L g1760 ( .A(n_1761), .Y(n_1760) );
NOR2x1_ASAP7_75t_L g1761 ( .A(n_1762), .B(n_1786), .Y(n_1761) );
A2O1A1Ixp33_ASAP7_75t_L g1762 ( .A1(n_1763), .A2(n_1767), .B(n_1783), .C(n_1784), .Y(n_1762) );
NOR3xp33_ASAP7_75t_SL g1767 ( .A(n_1768), .B(n_1776), .C(n_1777), .Y(n_1767) );
INVx1_ASAP7_75t_L g1769 ( .A(n_1770), .Y(n_1769) );
INVx1_ASAP7_75t_L g1771 ( .A(n_1772), .Y(n_1771) );
INVx1_ASAP7_75t_L g1778 ( .A(n_1779), .Y(n_1778) );
INVx1_ASAP7_75t_L g1779 ( .A(n_1780), .Y(n_1779) );
NAND2xp5_ASAP7_75t_L g1786 ( .A(n_1787), .B(n_1794), .Y(n_1786) );
INVx1_ASAP7_75t_L g1797 ( .A(n_1798), .Y(n_1797) );
CKINVDCx5p33_ASAP7_75t_R g1806 ( .A(n_1807), .Y(n_1806) );
HB1xp67_ASAP7_75t_L g1807 ( .A(n_1808), .Y(n_1807) );
BUFx3_ASAP7_75t_L g1808 ( .A(n_1809), .Y(n_1808) );
BUFx3_ASAP7_75t_L g1811 ( .A(n_1812), .Y(n_1811) );
INVx1_ASAP7_75t_L g1814 ( .A(n_1815), .Y(n_1814) );
XNOR2x1_ASAP7_75t_L g1815 ( .A(n_1816), .B(n_1865), .Y(n_1815) );
OR2x2_ASAP7_75t_L g1816 ( .A(n_1817), .B(n_1832), .Y(n_1816) );
NAND3xp33_ASAP7_75t_L g1817 ( .A(n_1818), .B(n_1823), .C(n_1830), .Y(n_1817) );
NAND3xp33_ASAP7_75t_SL g1832 ( .A(n_1833), .B(n_1837), .C(n_1862), .Y(n_1832) );
OAI21xp33_ASAP7_75t_L g1843 ( .A1(n_1844), .A2(n_1845), .B(n_1849), .Y(n_1843) );
INVx2_ASAP7_75t_L g1846 ( .A(n_1847), .Y(n_1846) );
INVx1_ASAP7_75t_L g1852 ( .A(n_1853), .Y(n_1852) );
NAND2xp5_ASAP7_75t_L g1862 ( .A(n_1863), .B(n_1864), .Y(n_1862) );
INVx1_ASAP7_75t_L g1866 ( .A(n_1867), .Y(n_1866) );
INVx1_ASAP7_75t_L g1867 ( .A(n_1868), .Y(n_1867) );
INVx1_ASAP7_75t_L g1870 ( .A(n_1871), .Y(n_1870) );
endmodule