module real_aes_7389_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_746;
wire n_153;
wire n_284;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_385;
wire n_358;
wire n_214;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g482 ( .A1(n_0), .A2(n_165), .B(n_483), .C(n_486), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_1), .B(n_477), .Y(n_488) );
INVx1_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
INVx1_ASAP7_75t_L g203 ( .A(n_3), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_4), .B(n_166), .Y(n_560) );
OAI22xp5_ASAP7_75t_SL g143 ( .A1(n_5), .A2(n_144), .B1(n_145), .B2(n_451), .Y(n_143) );
CKINVDCx16_ASAP7_75t_R g451 ( .A(n_5), .Y(n_451) );
OAI22xp5_ASAP7_75t_SL g749 ( .A1(n_5), .A2(n_98), .B1(n_451), .B2(n_750), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_6), .A2(n_106), .B1(n_117), .B2(n_757), .Y(n_105) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_7), .A2(n_462), .B(n_509), .Y(n_508) );
AO21x2_ASAP7_75t_L g539 ( .A1(n_8), .A2(n_172), .B(n_540), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_9), .A2(n_39), .B1(n_169), .B2(n_221), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_10), .B(n_172), .Y(n_189) );
AND2x6_ASAP7_75t_L g174 ( .A(n_11), .B(n_175), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_12), .A2(n_174), .B(n_465), .C(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g109 ( .A(n_13), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_13), .B(n_40), .Y(n_128) );
INVx1_ASAP7_75t_L g156 ( .A(n_14), .Y(n_156) );
INVx1_ASAP7_75t_L g195 ( .A(n_15), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_16), .B(n_162), .Y(n_215) );
OAI22xp5_ASAP7_75t_SL g753 ( .A1(n_17), .A2(n_42), .B1(n_537), .B2(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_17), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_18), .B(n_166), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_19), .B(n_152), .Y(n_151) );
AO32x2_ASAP7_75t_L g232 ( .A1(n_20), .A2(n_172), .A3(n_173), .B1(n_192), .B2(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_21), .B(n_169), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_22), .B(n_152), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_23), .A2(n_55), .B1(n_169), .B2(n_221), .Y(n_235) );
AOI22xp33_ASAP7_75t_SL g229 ( .A1(n_24), .A2(n_83), .B1(n_162), .B2(n_169), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_25), .B(n_169), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_26), .A2(n_173), .B(n_465), .C(n_467), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_27), .A2(n_173), .B(n_465), .C(n_543), .Y(n_542) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_28), .Y(n_160) );
OAI22xp5_ASAP7_75t_L g136 ( .A1(n_29), .A2(n_99), .B1(n_137), .B2(n_138), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_29), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_30), .B(n_211), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_31), .A2(n_462), .B(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_32), .B(n_211), .Y(n_248) );
INVx2_ASAP7_75t_L g164 ( .A(n_33), .Y(n_164) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_34), .A2(n_497), .B(n_498), .C(n_502), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_35), .B(n_169), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_36), .B(n_211), .Y(n_223) );
OAI22xp5_ASAP7_75t_SL g135 ( .A1(n_37), .A2(n_136), .B1(n_139), .B2(n_140), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_37), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_38), .B(n_217), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_40), .B(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_41), .B(n_461), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_42), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_43), .B(n_166), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_44), .B(n_462), .Y(n_541) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_45), .A2(n_497), .B(n_502), .C(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_46), .B(n_169), .Y(n_182) );
INVx1_ASAP7_75t_L g484 ( .A(n_47), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_48), .A2(n_752), .B1(n_753), .B2(n_755), .Y(n_751) );
INVx1_ASAP7_75t_L g755 ( .A(n_48), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_49), .A2(n_92), .B1(n_221), .B2(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g523 ( .A(n_50), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_51), .B(n_169), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_52), .B(n_169), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_53), .B(n_462), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_54), .B(n_187), .Y(n_186) );
AOI22xp33_ASAP7_75t_SL g168 ( .A1(n_56), .A2(n_61), .B1(n_162), .B2(n_169), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g132 ( .A1(n_57), .A2(n_133), .B1(n_134), .B2(n_135), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_57), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_58), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_59), .B(n_169), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_60), .B(n_169), .Y(n_268) );
INVx1_ASAP7_75t_L g175 ( .A(n_62), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_63), .B(n_462), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_64), .B(n_477), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_65), .A2(n_187), .B(n_198), .C(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_66), .B(n_169), .Y(n_204) );
INVx1_ASAP7_75t_L g155 ( .A(n_67), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_68), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_69), .B(n_166), .Y(n_500) );
AO32x2_ASAP7_75t_L g225 ( .A1(n_70), .A2(n_172), .A3(n_173), .B1(n_226), .B2(n_230), .Y(n_225) );
AOI222xp33_ASAP7_75t_SL g130 ( .A1(n_71), .A2(n_131), .B1(n_132), .B2(n_141), .C1(n_735), .C2(n_741), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_72), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_73), .B(n_167), .Y(n_534) );
INVx1_ASAP7_75t_L g267 ( .A(n_74), .Y(n_267) );
INVx1_ASAP7_75t_L g243 ( .A(n_75), .Y(n_243) );
CKINVDCx16_ASAP7_75t_R g480 ( .A(n_76), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_77), .B(n_469), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g557 ( .A1(n_78), .A2(n_465), .B(n_502), .C(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_79), .B(n_162), .Y(n_244) );
CKINVDCx16_ASAP7_75t_R g510 ( .A(n_80), .Y(n_510) );
INVx1_ASAP7_75t_L g116 ( .A(n_81), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_82), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_84), .B(n_221), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_85), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_86), .B(n_162), .Y(n_247) );
INVx2_ASAP7_75t_L g153 ( .A(n_87), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_88), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_89), .B(n_159), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_90), .B(n_162), .Y(n_183) );
INVx2_ASAP7_75t_L g113 ( .A(n_91), .Y(n_113) );
OR2x2_ASAP7_75t_L g125 ( .A(n_91), .B(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g452 ( .A(n_91), .B(n_127), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g161 ( .A1(n_93), .A2(n_104), .B1(n_162), .B2(n_163), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_94), .B(n_462), .Y(n_495) );
INVx1_ASAP7_75t_L g499 ( .A(n_95), .Y(n_499) );
INVxp67_ASAP7_75t_L g513 ( .A(n_96), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_97), .B(n_162), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_98), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_99), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_100), .B(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g530 ( .A(n_101), .Y(n_530) );
INVx1_ASAP7_75t_L g559 ( .A(n_102), .Y(n_559) );
AND2x2_ASAP7_75t_L g525 ( .A(n_103), .B(n_211), .Y(n_525) );
INVx2_ASAP7_75t_L g759 ( .A(n_106), .Y(n_759) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
CKINVDCx14_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_112), .B(n_113), .C(n_114), .Y(n_111) );
AND2x2_ASAP7_75t_L g127 ( .A(n_112), .B(n_128), .Y(n_127) );
OR2x2_ASAP7_75t_L g734 ( .A(n_113), .B(n_127), .Y(n_734) );
NOR2x2_ASAP7_75t_L g743 ( .A(n_113), .B(n_126), .Y(n_743) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
AOI22x1_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_130), .B1(n_744), .B2(n_745), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_122), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_SL g744 ( .A(n_120), .Y(n_744) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_122), .A2(n_746), .B(n_756), .Y(n_745) );
NOR2xp33_ASAP7_75t_SL g122 ( .A(n_123), .B(n_129), .Y(n_122) );
INVx1_ASAP7_75t_SL g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_SL g124 ( .A(n_125), .Y(n_124) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_125), .Y(n_756) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g139 ( .A(n_136), .Y(n_139) );
OAI22xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_452), .B1(n_453), .B2(n_734), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
OAI22xp5_ASAP7_75t_SL g735 ( .A1(n_143), .A2(n_736), .B1(n_738), .B2(n_739), .Y(n_735) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
XNOR2xp5_ASAP7_75t_L g748 ( .A(n_145), .B(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_SL g145 ( .A(n_146), .B(n_385), .Y(n_145) );
NOR5xp2_ASAP7_75t_L g146 ( .A(n_147), .B(n_298), .C(n_344), .D(n_357), .E(n_369), .Y(n_146) );
OAI211xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_206), .B(n_252), .C(n_279), .Y(n_147) );
INVx1_ASAP7_75t_SL g380 ( .A(n_148), .Y(n_380) );
OR2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_176), .Y(n_148) );
AND2x2_ASAP7_75t_L g304 ( .A(n_149), .B(n_177), .Y(n_304) );
AND2x2_ASAP7_75t_L g332 ( .A(n_149), .B(n_278), .Y(n_332) );
AND2x2_ASAP7_75t_L g340 ( .A(n_149), .B(n_283), .Y(n_340) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g270 ( .A(n_150), .B(n_178), .Y(n_270) );
INVx2_ASAP7_75t_L g282 ( .A(n_150), .Y(n_282) );
AND2x2_ASAP7_75t_L g407 ( .A(n_150), .B(n_349), .Y(n_407) );
OR2x2_ASAP7_75t_L g409 ( .A(n_150), .B(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g150 ( .A(n_151), .B(n_157), .Y(n_150) );
INVx1_ASAP7_75t_L g276 ( .A(n_151), .Y(n_276) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_152), .Y(n_172) );
INVx1_ASAP7_75t_L g192 ( .A(n_152), .Y(n_192) );
AND2x2_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
AND2x2_ASAP7_75t_SL g211 ( .A(n_153), .B(n_154), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
NAND3xp33_ASAP7_75t_L g157 ( .A(n_158), .B(n_171), .C(n_173), .Y(n_157) );
AO21x1_ASAP7_75t_L g275 ( .A1(n_158), .A2(n_171), .B(n_276), .Y(n_275) );
OAI22xp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_161), .B1(n_165), .B2(n_168), .Y(n_158) );
INVx2_ASAP7_75t_L g222 ( .A(n_159), .Y(n_222) );
OAI22xp5_ASAP7_75t_SL g226 ( .A1(n_159), .A2(n_167), .B1(n_227), .B2(n_229), .Y(n_226) );
OAI22xp5_ASAP7_75t_L g233 ( .A1(n_159), .A2(n_165), .B1(n_234), .B2(n_235), .Y(n_233) );
INVx4_ASAP7_75t_L g485 ( .A(n_159), .Y(n_485) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx3_ASAP7_75t_L g167 ( .A(n_160), .Y(n_167) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_160), .Y(n_200) );
INVx1_ASAP7_75t_L g217 ( .A(n_160), .Y(n_217) );
AND2x2_ASAP7_75t_L g463 ( .A(n_160), .B(n_188), .Y(n_463) );
INVx1_ASAP7_75t_L g466 ( .A(n_160), .Y(n_466) );
INVx2_ASAP7_75t_L g196 ( .A(n_162), .Y(n_196) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g170 ( .A(n_164), .Y(n_170) );
INVx1_ASAP7_75t_L g188 ( .A(n_164), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_165), .A2(n_185), .B(n_186), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_165), .A2(n_202), .B(n_203), .C(n_204), .Y(n_201) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_166), .A2(n_182), .B(n_183), .Y(n_181) );
O2A1O1Ixp5_ASAP7_75t_SL g241 ( .A1(n_166), .A2(n_242), .B(n_243), .C(n_244), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_166), .A2(n_264), .B(n_265), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_166), .B(n_513), .Y(n_512) );
INVx5_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx3_ASAP7_75t_L g242 ( .A(n_169), .Y(n_242) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_169), .Y(n_561) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g221 ( .A(n_170), .Y(n_221) );
BUFx3_ASAP7_75t_L g228 ( .A(n_170), .Y(n_228) );
AND2x6_ASAP7_75t_L g465 ( .A(n_170), .B(n_466), .Y(n_465) );
INVx3_ASAP7_75t_L g477 ( .A(n_171), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_171), .B(n_504), .Y(n_503) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_171), .A2(n_529), .B(n_536), .Y(n_528) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_171), .A2(n_556), .B(n_563), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_171), .B(n_564), .Y(n_563) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OA21x2_ASAP7_75t_L g179 ( .A1(n_172), .A2(n_180), .B(n_189), .Y(n_179) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_172), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_172), .A2(n_541), .B(n_542), .Y(n_540) );
OAI21xp5_ASAP7_75t_L g262 ( .A1(n_173), .A2(n_263), .B(n_266), .Y(n_262) );
BUFx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
OAI21xp5_ASAP7_75t_L g180 ( .A1(n_174), .A2(n_181), .B(n_184), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g193 ( .A1(n_174), .A2(n_194), .B(n_201), .Y(n_193) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_174), .A2(n_213), .B(n_218), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g240 ( .A1(n_174), .A2(n_241), .B(n_245), .Y(n_240) );
AND2x4_ASAP7_75t_L g462 ( .A(n_174), .B(n_463), .Y(n_462) );
INVx4_ASAP7_75t_SL g487 ( .A(n_174), .Y(n_487) );
NAND2x1p5_ASAP7_75t_L g531 ( .A(n_174), .B(n_463), .Y(n_531) );
INVx2_ASAP7_75t_SL g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g320 ( .A(n_177), .B(n_292), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_177), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g434 ( .A(n_177), .B(n_274), .Y(n_434) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_190), .Y(n_177) );
AND2x2_ASAP7_75t_L g277 ( .A(n_178), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g324 ( .A(n_178), .Y(n_324) );
AND2x2_ASAP7_75t_L g349 ( .A(n_178), .B(n_261), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_178), .B(n_382), .Y(n_419) );
INVx3_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g283 ( .A(n_179), .B(n_261), .Y(n_283) );
AND2x2_ASAP7_75t_L g297 ( .A(n_179), .B(n_260), .Y(n_297) );
AND2x2_ASAP7_75t_L g314 ( .A(n_179), .B(n_190), .Y(n_314) );
AND2x2_ASAP7_75t_L g371 ( .A(n_179), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_179), .B(n_278), .Y(n_384) );
AND2x2_ASAP7_75t_L g436 ( .A(n_179), .B(n_361), .Y(n_436) );
INVx2_ASAP7_75t_L g202 ( .A(n_187), .Y(n_202) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g259 ( .A(n_190), .B(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g278 ( .A(n_190), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_190), .B(n_261), .Y(n_355) );
OA21x2_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_193), .B(n_205), .Y(n_190) );
OA21x2_ASAP7_75t_L g261 ( .A1(n_191), .A2(n_262), .B(n_269), .Y(n_261) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_192), .B(n_537), .Y(n_536) );
O2A1O1Ixp33_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_197), .C(n_198), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_196), .A2(n_534), .B(n_535), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_196), .A2(n_544), .B(n_545), .Y(n_543) );
O2A1O1Ixp33_ASAP7_75t_L g558 ( .A1(n_198), .A2(n_559), .B(n_560), .C(n_561), .Y(n_558) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_199), .A2(n_246), .B(n_247), .Y(n_245) );
INVx4_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g469 ( .A(n_200), .Y(n_469) );
O2A1O1Ixp5_ASAP7_75t_L g266 ( .A1(n_202), .A2(n_222), .B(n_267), .C(n_268), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_202), .A2(n_468), .B(n_470), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_236), .B(n_249), .Y(n_206) );
INVx1_ASAP7_75t_SL g368 ( .A(n_207), .Y(n_368) );
AND2x4_ASAP7_75t_L g207 ( .A(n_208), .B(n_224), .Y(n_207) );
BUFx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_SL g256 ( .A(n_209), .B(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g251 ( .A(n_210), .Y(n_251) );
INVx1_ASAP7_75t_L g288 ( .A(n_210), .Y(n_288) );
AND2x2_ASAP7_75t_L g309 ( .A(n_210), .B(n_231), .Y(n_309) );
AND2x2_ASAP7_75t_L g343 ( .A(n_210), .B(n_232), .Y(n_343) );
OR2x2_ASAP7_75t_L g362 ( .A(n_210), .B(n_238), .Y(n_362) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_210), .Y(n_376) );
AND2x2_ASAP7_75t_L g389 ( .A(n_210), .B(n_390), .Y(n_389) );
OA21x2_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_223), .Y(n_210) );
INVx2_ASAP7_75t_L g230 ( .A(n_211), .Y(n_230) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_211), .A2(n_240), .B(n_248), .Y(n_239) );
INVx1_ASAP7_75t_L g475 ( .A(n_211), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_211), .A2(n_495), .B(n_496), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_211), .A2(n_520), .B(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_216), .Y(n_213) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_222), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g310 ( .A1(n_224), .A2(n_311), .B1(n_312), .B2(n_321), .Y(n_310) );
AND2x2_ASAP7_75t_L g394 ( .A(n_224), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_231), .Y(n_224) );
INVx1_ASAP7_75t_L g255 ( .A(n_225), .Y(n_255) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_225), .Y(n_292) );
INVx1_ASAP7_75t_L g303 ( .A(n_225), .Y(n_303) );
AND2x2_ASAP7_75t_L g318 ( .A(n_225), .B(n_232), .Y(n_318) );
INVx2_ASAP7_75t_L g486 ( .A(n_228), .Y(n_486) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_228), .Y(n_501) );
INVx1_ASAP7_75t_L g472 ( .A(n_230), .Y(n_472) );
OR2x2_ASAP7_75t_L g272 ( .A(n_231), .B(n_257), .Y(n_272) );
AND2x2_ASAP7_75t_L g302 ( .A(n_231), .B(n_303), .Y(n_302) );
NOR2xp67_ASAP7_75t_L g390 ( .A(n_231), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g250 ( .A(n_232), .B(n_251), .Y(n_250) );
BUFx2_ASAP7_75t_L g359 ( .A(n_232), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_236), .B(n_375), .Y(n_374) );
BUFx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g337 ( .A(n_237), .B(n_303), .Y(n_337) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g249 ( .A(n_238), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g308 ( .A(n_238), .Y(n_308) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g257 ( .A(n_239), .Y(n_257) );
OR2x2_ASAP7_75t_L g287 ( .A(n_239), .B(n_288), .Y(n_287) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_239), .Y(n_342) );
AOI32xp33_ASAP7_75t_L g379 ( .A1(n_249), .A2(n_309), .A3(n_380), .B1(n_381), .B2(n_383), .Y(n_379) );
AND2x2_ASAP7_75t_L g305 ( .A(n_250), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_250), .B(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_250), .B(n_337), .Y(n_423) );
INVx1_ASAP7_75t_L g428 ( .A(n_250), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_258), .B1(n_271), .B2(n_273), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
AND2x2_ASAP7_75t_L g358 ( .A(n_254), .B(n_359), .Y(n_358) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_255), .B(n_257), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_256), .A2(n_280), .B1(n_284), .B2(n_294), .Y(n_279) );
AND2x2_ASAP7_75t_L g301 ( .A(n_256), .B(n_302), .Y(n_301) );
A2O1A1Ixp33_ASAP7_75t_L g352 ( .A1(n_256), .A2(n_270), .B(n_318), .C(n_353), .Y(n_352) );
OAI332xp33_ASAP7_75t_L g357 ( .A1(n_256), .A2(n_358), .A3(n_360), .B1(n_362), .B2(n_363), .B3(n_365), .C1(n_366), .C2(n_368), .Y(n_357) );
INVx2_ASAP7_75t_L g398 ( .A(n_256), .Y(n_398) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_257), .Y(n_316) );
INVx1_ASAP7_75t_L g391 ( .A(n_257), .Y(n_391) );
AND2x2_ASAP7_75t_L g445 ( .A(n_257), .B(n_309), .Y(n_445) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_270), .Y(n_258) );
AND2x2_ASAP7_75t_L g325 ( .A(n_260), .B(n_275), .Y(n_325) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g274 ( .A(n_261), .B(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g373 ( .A(n_261), .B(n_275), .Y(n_373) );
INVx1_ASAP7_75t_L g382 ( .A(n_261), .Y(n_382) );
INVx1_ASAP7_75t_L g356 ( .A(n_270), .Y(n_356) );
INVxp67_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g440 ( .A(n_272), .B(n_292), .Y(n_440) );
INVx1_ASAP7_75t_SL g351 ( .A(n_273), .Y(n_351) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_277), .Y(n_273) );
AND2x2_ASAP7_75t_L g378 ( .A(n_274), .B(n_336), .Y(n_378) );
INVx1_ASAP7_75t_L g397 ( .A(n_274), .Y(n_397) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_274), .B(n_364), .Y(n_399) );
INVx1_ASAP7_75t_L g296 ( .A(n_275), .Y(n_296) );
AND2x2_ASAP7_75t_L g300 ( .A(n_277), .B(n_281), .Y(n_300) );
AND2x2_ASAP7_75t_L g367 ( .A(n_277), .B(n_325), .Y(n_367) );
INVx2_ASAP7_75t_L g410 ( .A(n_277), .Y(n_410) );
INVx2_ASAP7_75t_L g293 ( .A(n_278), .Y(n_293) );
AND2x2_ASAP7_75t_L g295 ( .A(n_278), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
INVx1_ASAP7_75t_L g311 ( .A(n_281), .Y(n_311) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_282), .B(n_355), .Y(n_361) );
OR2x2_ASAP7_75t_L g425 ( .A(n_282), .B(n_384), .Y(n_425) );
INVx1_ASAP7_75t_L g449 ( .A(n_282), .Y(n_449) );
INVx1_ASAP7_75t_L g405 ( .A(n_283), .Y(n_405) );
AND2x2_ASAP7_75t_L g450 ( .A(n_283), .B(n_293), .Y(n_450) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_289), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_287), .A2(n_313), .B1(n_315), .B2(n_319), .Y(n_312) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OAI322xp33_ASAP7_75t_SL g396 ( .A1(n_290), .A2(n_397), .A3(n_398), .B1(n_399), .B2(n_400), .C1(n_403), .C2(n_405), .Y(n_396) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
AND2x2_ASAP7_75t_L g393 ( .A(n_291), .B(n_309), .Y(n_393) );
OR2x2_ASAP7_75t_L g427 ( .A(n_291), .B(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g430 ( .A(n_291), .B(n_362), .Y(n_430) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g375 ( .A(n_292), .B(n_376), .Y(n_375) );
OR2x2_ASAP7_75t_L g431 ( .A(n_292), .B(n_362), .Y(n_431) );
INVx3_ASAP7_75t_L g364 ( .A(n_293), .Y(n_364) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
INVx1_ASAP7_75t_L g420 ( .A(n_295), .Y(n_420) );
AOI222xp33_ASAP7_75t_L g299 ( .A1(n_297), .A2(n_300), .B1(n_301), .B2(n_304), .C1(n_305), .C2(n_307), .Y(n_299) );
INVx1_ASAP7_75t_L g330 ( .A(n_297), .Y(n_330) );
NAND3xp33_ASAP7_75t_SL g298 ( .A(n_299), .B(n_310), .C(n_327), .Y(n_298) );
AND2x2_ASAP7_75t_L g415 ( .A(n_302), .B(n_316), .Y(n_415) );
BUFx2_ASAP7_75t_L g306 ( .A(n_303), .Y(n_306) );
INVx1_ASAP7_75t_L g347 ( .A(n_303), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_304), .A2(n_340), .B1(n_393), .B2(n_394), .C(n_396), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_306), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_309), .Y(n_333) );
AND2x2_ASAP7_75t_L g346 ( .A(n_309), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_314), .B(n_325), .Y(n_326) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
OAI21xp33_ASAP7_75t_L g321 ( .A1(n_316), .A2(n_322), .B(n_326), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_316), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g413 ( .A(n_318), .B(n_395), .Y(n_413) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g336 ( .A(n_324), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_325), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g442 ( .A(n_325), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_333), .B1(n_334), .B2(n_337), .C(n_338), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_329), .B(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g438 ( .A(n_337), .B(n_343), .Y(n_438) );
INVxp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
OAI31xp33_ASAP7_75t_SL g406 ( .A1(n_341), .A2(n_380), .A3(n_407), .B(n_408), .Y(n_406) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx1_ASAP7_75t_L g395 ( .A(n_342), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_343), .B(n_347), .Y(n_446) );
OAI221xp5_ASAP7_75t_SL g344 ( .A1(n_345), .A2(n_348), .B1(n_350), .B2(n_351), .C(n_352), .Y(n_344) );
INVx1_ASAP7_75t_L g350 ( .A(n_346), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_349), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g365 ( .A(n_358), .Y(n_365) );
INVx2_ASAP7_75t_L g401 ( .A(n_359), .Y(n_401) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g387 ( .A(n_364), .B(n_373), .Y(n_387) );
A2O1A1Ixp33_ASAP7_75t_L g437 ( .A1(n_364), .A2(n_381), .B(n_438), .C(n_439), .Y(n_437) );
OAI221xp5_ASAP7_75t_SL g369 ( .A1(n_365), .A2(n_370), .B1(n_374), .B2(n_377), .C(n_379), .Y(n_369) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
A2O1A1Ixp33_ASAP7_75t_L g432 ( .A1(n_368), .A2(n_433), .B(n_435), .C(n_437), .Y(n_432) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_371), .A2(n_422), .B1(n_424), .B2(n_426), .C(n_429), .Y(n_421) );
INVx1_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
NOR4xp25_ASAP7_75t_L g385 ( .A(n_386), .B(n_411), .C(n_432), .D(n_443), .Y(n_385) );
OAI211xp5_ASAP7_75t_SL g386 ( .A1(n_387), .A2(n_388), .B(n_392), .C(n_406), .Y(n_386) );
INVx1_ASAP7_75t_SL g441 ( .A(n_393), .Y(n_441) );
OR2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
INVx1_ASAP7_75t_SL g404 ( .A(n_402), .Y(n_404) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_409), .A2(n_418), .B1(n_430), .B2(n_431), .Y(n_429) );
A2O1A1Ixp33_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_414), .B(n_416), .C(n_421), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AOI31xp33_ASAP7_75t_L g443 ( .A1(n_414), .A2(n_444), .A3(n_446), .B(n_447), .Y(n_443) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OR2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
AOI21xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B(n_442), .Y(n_439) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_450), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g737 ( .A(n_452), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_453), .Y(n_738) );
AND2x2_ASAP7_75t_SL g453 ( .A(n_454), .B(n_670), .Y(n_453) );
NOR5xp2_ASAP7_75t_L g454 ( .A(n_455), .B(n_601), .C(n_630), .D(n_650), .E(n_657), .Y(n_454) );
OAI211xp5_ASAP7_75t_SL g455 ( .A1(n_456), .A2(n_489), .B(n_546), .C(n_588), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_457), .A2(n_673), .B1(n_675), .B2(n_676), .Y(n_672) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_476), .Y(n_457) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_458), .Y(n_549) );
AND2x4_ASAP7_75t_L g581 ( .A(n_458), .B(n_582), .Y(n_581) );
INVx5_ASAP7_75t_L g599 ( .A(n_458), .Y(n_599) );
AND2x2_ASAP7_75t_L g608 ( .A(n_458), .B(n_600), .Y(n_608) );
AND2x2_ASAP7_75t_L g620 ( .A(n_458), .B(n_493), .Y(n_620) );
AND2x2_ASAP7_75t_L g716 ( .A(n_458), .B(n_584), .Y(n_716) );
OR2x6_ASAP7_75t_L g458 ( .A(n_459), .B(n_473), .Y(n_458) );
AOI21xp5_ASAP7_75t_SL g459 ( .A1(n_460), .A2(n_464), .B(n_472), .Y(n_459) );
BUFx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx5_ASAP7_75t_L g481 ( .A(n_465), .Y(n_481) );
INVx2_ASAP7_75t_L g471 ( .A(n_469), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g498 ( .A1(n_471), .A2(n_499), .B(n_500), .C(n_501), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_471), .A2(n_501), .B(n_523), .C(n_524), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
INVx2_ASAP7_75t_L g582 ( .A(n_476), .Y(n_582) );
AND2x2_ASAP7_75t_L g600 ( .A(n_476), .B(n_555), .Y(n_600) );
AND2x2_ASAP7_75t_L g619 ( .A(n_476), .B(n_554), .Y(n_619) );
AND2x2_ASAP7_75t_L g659 ( .A(n_476), .B(n_599), .Y(n_659) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B(n_488), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_SL g479 ( .A1(n_480), .A2(n_481), .B(n_482), .C(n_487), .Y(n_479) );
INVx2_ASAP7_75t_L g497 ( .A(n_481), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_481), .A2(n_487), .B(n_510), .C(n_511), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
INVx1_ASAP7_75t_L g502 ( .A(n_487), .Y(n_502) );
INVxp67_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_491), .B(n_515), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AOI322xp5_ASAP7_75t_L g718 ( .A1(n_492), .A2(n_526), .A3(n_573), .B1(n_581), .B2(n_635), .C1(n_719), .C2(n_722), .Y(n_718) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_505), .Y(n_492) );
INVx5_ASAP7_75t_L g551 ( .A(n_493), .Y(n_551) );
AND2x2_ASAP7_75t_L g567 ( .A(n_493), .B(n_553), .Y(n_567) );
BUFx2_ASAP7_75t_L g645 ( .A(n_493), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_493), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g722 ( .A(n_493), .B(n_629), .Y(n_722) );
OR2x6_ASAP7_75t_L g493 ( .A(n_494), .B(n_503), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_505), .B(n_517), .Y(n_576) );
INVx1_ASAP7_75t_L g603 ( .A(n_505), .Y(n_603) );
AND2x2_ASAP7_75t_L g616 ( .A(n_505), .B(n_538), .Y(n_616) );
AND2x2_ASAP7_75t_L g717 ( .A(n_505), .B(n_635), .Y(n_717) );
INVx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g571 ( .A(n_506), .B(n_517), .Y(n_571) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_506), .Y(n_579) );
OR2x2_ASAP7_75t_L g586 ( .A(n_506), .B(n_538), .Y(n_586) );
AND2x2_ASAP7_75t_L g596 ( .A(n_506), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_506), .B(n_528), .Y(n_625) );
INVxp67_ASAP7_75t_L g649 ( .A(n_506), .Y(n_649) );
AND2x2_ASAP7_75t_L g656 ( .A(n_506), .B(n_526), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_506), .B(n_538), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_506), .B(n_527), .Y(n_682) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B(n_514), .Y(n_506) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_526), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_517), .B(n_539), .Y(n_626) );
OR2x2_ASAP7_75t_L g648 ( .A(n_517), .B(n_527), .Y(n_648) );
AND2x2_ASAP7_75t_L g661 ( .A(n_517), .B(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_517), .B(n_616), .Y(n_667) );
OAI211xp5_ASAP7_75t_SL g671 ( .A1(n_517), .A2(n_672), .B(n_677), .C(n_686), .Y(n_671) );
AND2x2_ASAP7_75t_L g732 ( .A(n_517), .B(n_538), .Y(n_732) );
INVx5_ASAP7_75t_SL g517 ( .A(n_518), .Y(n_517) );
OR2x2_ASAP7_75t_L g585 ( .A(n_518), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_518), .B(n_591), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_518), .B(n_580), .Y(n_592) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_518), .Y(n_594) );
OR2x2_ASAP7_75t_L g605 ( .A(n_518), .B(n_527), .Y(n_605) );
AND2x2_ASAP7_75t_SL g610 ( .A(n_518), .B(n_596), .Y(n_610) );
AND2x2_ASAP7_75t_L g635 ( .A(n_518), .B(n_527), .Y(n_635) );
AND2x2_ASAP7_75t_L g655 ( .A(n_518), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g693 ( .A(n_518), .B(n_526), .Y(n_693) );
OR2x2_ASAP7_75t_L g696 ( .A(n_518), .B(n_682), .Y(n_696) );
OR2x6_ASAP7_75t_L g518 ( .A(n_519), .B(n_525), .Y(n_518) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_538), .Y(n_526) );
A2O1A1Ixp33_ASAP7_75t_L g639 ( .A1(n_527), .A2(n_640), .B(n_643), .C(n_649), .Y(n_639) );
INVx5_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_528), .B(n_538), .Y(n_570) );
AND2x2_ASAP7_75t_L g574 ( .A(n_528), .B(n_539), .Y(n_574) );
OR2x2_ASAP7_75t_L g580 ( .A(n_528), .B(n_538), .Y(n_580) );
OAI21xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B(n_532), .Y(n_529) );
INVx1_ASAP7_75t_SL g597 ( .A(n_538), .Y(n_597) );
OR2x2_ASAP7_75t_L g725 ( .A(n_538), .B(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
O2A1O1Ixp33_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_565), .B(n_568), .C(n_577), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AOI31xp33_ASAP7_75t_L g650 ( .A1(n_548), .A2(n_651), .A3(n_653), .B(n_654), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_549), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_550), .B(n_581), .Y(n_587) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_551), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g607 ( .A(n_551), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g612 ( .A(n_551), .B(n_582), .Y(n_612) );
AND2x2_ASAP7_75t_L g622 ( .A(n_551), .B(n_581), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_551), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g642 ( .A(n_551), .B(n_599), .Y(n_642) );
AND2x2_ASAP7_75t_L g647 ( .A(n_551), .B(n_619), .Y(n_647) );
OR2x2_ASAP7_75t_L g666 ( .A(n_551), .B(n_553), .Y(n_666) );
OR2x2_ASAP7_75t_L g668 ( .A(n_551), .B(n_669), .Y(n_668) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_551), .Y(n_715) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g615 ( .A(n_553), .B(n_582), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_553), .B(n_599), .Y(n_638) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
BUFx2_ASAP7_75t_L g584 ( .A(n_555), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_562), .Y(n_556) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g675 ( .A(n_567), .B(n_599), .Y(n_675) );
AOI322xp5_ASAP7_75t_L g677 ( .A1(n_567), .A2(n_581), .A3(n_619), .B1(n_678), .B2(n_679), .C1(n_680), .C2(n_683), .Y(n_677) );
INVx1_ASAP7_75t_L g685 ( .A(n_567), .Y(n_685) );
NAND2xp33_ASAP7_75t_L g568 ( .A(n_569), .B(n_572), .Y(n_568) );
INVx1_ASAP7_75t_SL g679 ( .A(n_569), .Y(n_679) );
OR2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
OR2x2_ASAP7_75t_L g631 ( .A(n_570), .B(n_576), .Y(n_631) );
INVx1_ASAP7_75t_L g662 ( .A(n_570), .Y(n_662) );
INVx2_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OAI32xp33_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_581), .A3(n_583), .B1(n_585), .B2(n_587), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
AOI21xp33_ASAP7_75t_SL g617 ( .A1(n_580), .A2(n_595), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_SL g632 ( .A(n_581), .Y(n_632) );
AND2x4_ASAP7_75t_L g629 ( .A(n_582), .B(n_599), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_582), .B(n_665), .Y(n_664) );
AOI322xp5_ASAP7_75t_L g694 ( .A1(n_583), .A2(n_610), .A3(n_629), .B1(n_662), .B2(n_695), .C1(n_697), .C2(n_698), .Y(n_694) );
OAI221xp5_ASAP7_75t_L g723 ( .A1(n_583), .A2(n_660), .B1(n_724), .B2(n_725), .C(n_727), .Y(n_723) );
AND2x2_ASAP7_75t_L g611 ( .A(n_584), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_SL g591 ( .A(n_586), .Y(n_591) );
OR2x2_ASAP7_75t_L g663 ( .A(n_586), .B(n_648), .Y(n_663) );
OAI31xp33_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_592), .A3(n_593), .B(n_598), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_589), .A2(n_622), .B1(n_623), .B2(n_627), .Y(n_621) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g634 ( .A(n_591), .B(n_635), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_593), .A2(n_634), .B1(n_687), .B2(n_690), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g676 ( .A(n_596), .B(n_645), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_596), .B(n_635), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_597), .B(n_703), .Y(n_702) );
OR2x2_ASAP7_75t_L g710 ( .A(n_597), .B(n_648), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_598), .A2(n_693), .B1(n_706), .B2(n_709), .Y(n_705) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx2_ASAP7_75t_L g614 ( .A(n_599), .Y(n_614) );
AND2x2_ASAP7_75t_L g697 ( .A(n_599), .B(n_619), .Y(n_697) );
OR2x2_ASAP7_75t_L g699 ( .A(n_599), .B(n_666), .Y(n_699) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_599), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_600), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_600), .B(n_645), .Y(n_653) );
OAI211xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_606), .B(n_609), .C(n_621), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B1(n_613), .B2(n_616), .C(n_617), .Y(n_609) );
INVxp67_ASAP7_75t_L g721 ( .A(n_612), .Y(n_721) );
INVx1_ASAP7_75t_L g688 ( .A(n_613), .Y(n_688) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
AND2x2_ASAP7_75t_L g652 ( .A(n_614), .B(n_619), .Y(n_652) );
INVx1_ASAP7_75t_L g669 ( .A(n_615), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_615), .B(n_642), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
INVx1_ASAP7_75t_L g684 ( .A(n_619), .Y(n_684) );
AND2x2_ASAP7_75t_L g690 ( .A(n_619), .B(n_645), .Y(n_690) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
INVx1_ASAP7_75t_SL g678 ( .A(n_626), .Y(n_678) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_629), .B(n_665), .Y(n_689) );
OAI221xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .B1(n_633), .B2(n_636), .C(n_639), .Y(n_630) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g726 ( .A(n_635), .Y(n_726) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g644 ( .A(n_638), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_642), .B(n_701), .Y(n_700) );
AOI21xp33_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_646), .B(n_648), .Y(n_643) );
OAI211xp5_ASAP7_75t_SL g691 ( .A1(n_646), .A2(n_692), .B(n_694), .C(n_700), .Y(n_691) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g703 ( .A(n_648), .Y(n_703) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI222xp33_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_660), .B1(n_663), .B2(n_664), .C1(n_667), .C2(n_668), .Y(n_657) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g733 ( .A(n_664), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_665), .B(n_708), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_665), .A2(n_712), .B1(n_714), .B2(n_717), .Y(n_711) );
INVx2_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
NOR4xp25_ASAP7_75t_L g670 ( .A(n_671), .B(n_691), .C(n_704), .D(n_723), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_673), .B(n_703), .Y(n_713) );
INVx1_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g680 ( .A(n_678), .B(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_681), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_688), .B(n_689), .Y(n_687) );
INVx1_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NAND3xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_711), .C(n_718), .Y(n_704) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
INVx2_ASAP7_75t_L g720 ( .A(n_716), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
OAI21xp5_ASAP7_75t_SL g727 ( .A1(n_728), .A2(n_730), .B(n_733), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g740 ( .A(n_734), .Y(n_740) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
XOR2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_751), .Y(n_746) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
endmodule