module real_jpeg_3938_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_19;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

INVx8_ASAP7_75t_L g94 ( 
.A(n_0),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_1),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_2),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_2),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_2),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_2),
.B(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_2),
.B(n_30),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_3),
.Y(n_97)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_3),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_3),
.Y(n_138)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_3),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_4),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_4),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_4),
.B(n_138),
.Y(n_137)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_6),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_7),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_7),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_7),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_7),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_8),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_8),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_8),
.B(n_132),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_8),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_8),
.B(n_73),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_8),
.B(n_34),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_8),
.B(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_9),
.Y(n_134)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_11),
.B(n_91),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_11),
.B(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_11),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_11),
.B(n_34),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_12),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_13),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_14),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_14),
.B(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_14),
.B(n_41),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_14),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_14),
.B(n_177),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_14),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_14),
.B(n_218),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_15),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_15),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_15),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_15),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_15),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_15),
.B(n_91),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_15),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_168),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_166),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_143),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_21),
.B(n_143),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_100),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_64),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_36),
.B2(n_63),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_33),
.Y(n_28)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_32),
.Y(n_111)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_32),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_35),
.Y(n_109)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_46),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_37),
.A2(n_38),
.B(n_40),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_43),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_45),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_52),
.C(n_57),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_47),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_104)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_58),
.B(n_236),
.Y(n_235)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_62),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_62),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_82),
.C(n_83),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_65),
.B(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_74),
.C(n_76),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_66),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_71),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_67),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_237)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_75),
.B(n_77),
.Y(n_250)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_85),
.B(n_95),
.C(n_98),
.Y(n_142)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.Y(n_89)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_92),
.Y(n_219)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_95),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_97),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_121),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.C(n_112),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_102),
.A2(n_103),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_106),
.B(n_113),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_107),
.B(n_110),
.Y(n_162)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

MAJx2_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.C(n_118),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_118),
.Y(n_149)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_119),
.Y(n_236)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_135),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_142),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.C(n_163),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_144),
.B(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_147),
.B(n_163),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.C(n_162),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_148),
.B(n_253),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_150),
.A2(n_151),
.B1(n_162),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_151),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_156),
.C(n_160),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_152),
.A2(n_153),
.B1(n_160),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_156),
.B(n_243),
.Y(n_242)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_160),
.Y(n_244)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_162),
.Y(n_254)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI21x1_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_257),
.B(n_262),
.Y(n_168)
);

AOI21x1_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_246),
.B(n_256),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_228),
.B(n_245),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_209),
.B(n_227),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_192),
.B(n_208),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_188),
.B(n_191),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_183),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_183),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_182),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_182),
.Y(n_193)
);

INVx4_ASAP7_75t_SL g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_194),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_200),
.B2(n_201),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_203),
.C(n_206),
.Y(n_226)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_198),
.Y(n_215)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_206),
.B2(n_207),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_226),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_226),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_216),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_215),
.C(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_214),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_240),
.C(n_241),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_221),
.Y(n_240)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_231),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_238),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_239),
.C(n_242),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_235),
.C(n_237),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_242),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_255),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_255),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_252),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_251),
.C(n_261),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_260),
.Y(n_262)
);


endmodule