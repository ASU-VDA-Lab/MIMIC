module fake_jpeg_23914_n_327 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_5),
.B(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_39),
.B(n_27),
.Y(n_70)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_28),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_27),
.Y(n_56)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_48),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_51),
.Y(n_91)
);

AOI21xp33_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_35),
.B(n_24),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_61),
.Y(n_95)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_67),
.Y(n_98)
);

NAND2x1_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_25),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_60),
.A2(n_73),
.B(n_36),
.Y(n_113)
);

NAND2xp33_ASAP7_75t_SL g61 ( 
.A(n_46),
.B(n_25),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_28),
.B1(n_37),
.B2(n_41),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_64),
.A2(n_40),
.B1(n_29),
.B2(n_21),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_39),
.A2(n_23),
.B1(n_34),
.B2(n_24),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_66),
.A2(n_26),
.B1(n_20),
.B2(n_18),
.Y(n_105)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_70),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_38),
.A2(n_37),
.B1(n_28),
.B2(n_27),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_77),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_41),
.B(n_22),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_75),
.B(n_22),
.Y(n_99)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_0),
.Y(n_112)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_80),
.B(n_81),
.Y(n_126)
);

INVxp33_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_37),
.B1(n_31),
.B2(n_38),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_82),
.A2(n_83),
.B1(n_89),
.B2(n_93),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_41),
.B1(n_40),
.B2(n_38),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_85),
.B(n_94),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_56),
.B(n_31),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_116),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_72),
.A2(n_31),
.B1(n_33),
.B2(n_29),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_90),
.A2(n_102),
.B1(n_105),
.B2(n_114),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_45),
.C(n_44),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_55),
.C(n_71),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_72),
.A2(n_33),
.B1(n_30),
.B2(n_21),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_77),
.A2(n_30),
.B1(n_34),
.B2(n_23),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_96),
.A2(n_106),
.B1(n_109),
.B2(n_113),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_99),
.B(n_12),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_61),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_0),
.Y(n_118)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_103),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_54),
.A2(n_26),
.B1(n_20),
.B2(n_18),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_104),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_65),
.A2(n_67),
.B1(n_78),
.B2(n_59),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_108),
.Y(n_142)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_65),
.A2(n_26),
.B1(n_20),
.B2(n_18),
.Y(n_109)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_64),
.A2(n_36),
.B1(n_26),
.B2(n_20),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_71),
.B(n_45),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_117),
.B(n_108),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g173 ( 
.A1(n_118),
.A2(n_128),
.B(n_136),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_71),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_138),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_134),
.C(n_135),
.Y(n_156)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_127),
.Y(n_157)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_79),
.B(n_0),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_129),
.B(n_143),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_104),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_132),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_113),
.C(n_100),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_58),
.C(n_57),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_95),
.B(n_0),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_141),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_45),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_99),
.B(n_74),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_151),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_44),
.B1(n_42),
.B2(n_36),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_145),
.A2(n_117),
.B1(n_84),
.B2(n_91),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_105),
.A2(n_44),
.B1(n_42),
.B2(n_36),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_146),
.A2(n_101),
.B1(n_94),
.B2(n_80),
.Y(n_176)
);

AND2x4_ASAP7_75t_L g148 ( 
.A(n_83),
.B(n_88),
.Y(n_148)
);

AO21x1_ASAP7_75t_L g180 ( 
.A1(n_148),
.A2(n_87),
.B(n_3),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_90),
.B(n_1),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_152),
.C(n_1),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_150),
.Y(n_177)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_91),
.B(n_42),
.C(n_25),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_119),
.B(n_86),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_155),
.B(n_160),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_165),
.Y(n_201)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_86),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_161),
.B(n_5),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_162),
.A2(n_133),
.B1(n_135),
.B2(n_145),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_119),
.B(n_110),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_167),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_130),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_130),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_171),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_121),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_168),
.B(n_169),
.Y(n_197)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_110),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_172),
.Y(n_199)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_115),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_149),
.B(n_115),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_175),
.B(n_182),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_176),
.A2(n_148),
.B1(n_122),
.B2(n_132),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_103),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_178),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_120),
.A2(n_25),
.B1(n_87),
.B2(n_4),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_179),
.A2(n_148),
.B1(n_133),
.B2(n_144),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_180),
.A2(n_181),
.B(n_147),
.Y(n_193)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_124),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_183),
.A2(n_148),
.B(n_118),
.Y(n_202)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_184),
.B(n_185),
.Y(n_203)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_187),
.B(n_189),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_159),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_188),
.Y(n_227)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

OAI211xp5_ASAP7_75t_L g225 ( 
.A1(n_191),
.A2(n_193),
.B(n_202),
.C(n_173),
.Y(n_225)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_192),
.B(n_195),
.Y(n_234)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_194),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_177),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_196),
.A2(n_206),
.B1(n_132),
.B2(n_174),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_172),
.B(n_128),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_204),
.B(n_210),
.Y(n_223)
);

AND2x2_ASAP7_75t_SL g205 ( 
.A(n_153),
.B(n_167),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_169),
.B(n_154),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_153),
.B(n_118),
.Y(n_207)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_161),
.B(n_128),
.Y(n_208)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_208),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_170),
.B(n_123),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_177),
.B(n_140),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_214),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_183),
.C(n_156),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_157),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_213),
.A2(n_166),
.B(n_7),
.Y(n_237)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_180),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_127),
.Y(n_215)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_215),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_192),
.A2(n_184),
.B1(n_156),
.B2(n_179),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_217),
.A2(n_222),
.B1(n_200),
.B2(n_234),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_212),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_168),
.C(n_160),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_221),
.B(n_235),
.C(n_199),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_225),
.A2(n_237),
.B(n_214),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_158),
.Y(n_226)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_240),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_186),
.B(n_174),
.Y(n_230)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_231),
.A2(n_238),
.B1(n_241),
.B2(n_191),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_6),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_242),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_166),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_206),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_207),
.Y(n_239)
);

AND2x4_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_205),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_205),
.A2(n_203),
.B(n_193),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_196),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_250),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_194),
.Y(n_247)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_251),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_242),
.B(n_187),
.Y(n_249)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_227),
.B(n_213),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_235),
.B(n_240),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_202),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_261),
.C(n_263),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_254),
.A2(n_256),
.B(n_226),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_218),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_190),
.Y(n_257)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_217),
.A2(n_203),
.B1(n_200),
.B2(n_195),
.Y(n_258)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_228),
.Y(n_259)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_259),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_260),
.A2(n_223),
.B1(n_218),
.B2(n_220),
.Y(n_265)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_262),
.A2(n_194),
.B1(n_236),
.B2(n_228),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_221),
.B(n_215),
.Y(n_263)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_255),
.A2(n_254),
.B(n_253),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_224),
.B(n_230),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_251),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_244),
.A2(n_224),
.B1(n_209),
.B2(n_220),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_275),
.A2(n_278),
.B1(n_211),
.B2(n_198),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_222),
.C(n_229),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_263),
.C(n_252),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_254),
.A2(n_239),
.B1(n_233),
.B2(n_238),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_243),
.A2(n_241),
.B1(n_239),
.B2(n_237),
.Y(n_281)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_281),
.Y(n_285)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_282),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_279),
.Y(n_284)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_245),
.Y(n_286)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_286),
.Y(n_304)
);

AND2x2_ASAP7_75t_SL g287 ( 
.A(n_266),
.B(n_243),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_287),
.A2(n_289),
.B(n_273),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_288),
.A2(n_292),
.B(n_278),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_259),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_295),
.C(n_270),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_188),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_294),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_277),
.A2(n_197),
.B1(n_190),
.B2(n_210),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_268),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_248),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_301),
.B(n_286),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_298),
.A2(n_293),
.B(n_283),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_267),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_295),
.C(n_280),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_285),
.A2(n_272),
.B1(n_271),
.B2(n_275),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_303),
.A2(n_288),
.B1(n_281),
.B2(n_289),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_270),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_282),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_307),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_276),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_308),
.A2(n_304),
.B1(n_297),
.B2(n_299),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_298),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_311),
.C(n_312),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_296),
.A2(n_287),
.B(n_197),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_287),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_297),
.C(n_300),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_316),
.A2(n_318),
.B1(n_315),
.B2(n_204),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_317),
.A2(n_311),
.B(n_10),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_308),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_321),
.B(n_316),
.Y(n_322)
);

OAI21x1_ASAP7_75t_L g323 ( 
.A1(n_320),
.A2(n_9),
.B(n_10),
.Y(n_323)
);

OAI21x1_ASAP7_75t_SL g324 ( 
.A1(n_322),
.A2(n_323),
.B(n_11),
.Y(n_324)
);

AO21x1_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_13),
.B(n_16),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_13),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_16),
.Y(n_327)
);


endmodule