module fake_jpeg_13964_n_226 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_226);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_4),
.B(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx2_ASAP7_75t_SL g85 ( 
.A(n_42),
.Y(n_85)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_8),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_46),
.B(n_56),
.Y(n_84)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_53),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_21),
.B(n_14),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_L g58 ( 
.A1(n_23),
.A2(n_38),
.B(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_61),
.Y(n_71)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_16),
.Y(n_78)
);

BUFx12f_ASAP7_75t_SL g61 ( 
.A(n_21),
.Y(n_61)
);

INVxp67_ASAP7_75t_SL g62 ( 
.A(n_16),
.Y(n_62)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_22),
.B(n_13),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_64),
.B(n_10),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_18),
.C(n_25),
.Y(n_67)
);

A2O1A1O1Ixp25_ASAP7_75t_L g100 ( 
.A1(n_67),
.A2(n_52),
.B(n_59),
.C(n_57),
.D(n_60),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_40),
.A2(n_18),
.B1(n_25),
.B2(n_38),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_34),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_79),
.B(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_34),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_39),
.A2(n_36),
.B1(n_35),
.B2(n_23),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_47),
.B1(n_41),
.B2(n_4),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_22),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_82),
.B(n_88),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_49),
.A2(n_35),
.B1(n_26),
.B2(n_17),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_86),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_30),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_30),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_93),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_42),
.B(n_17),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_44),
.Y(n_110)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

AO22x1_ASAP7_75t_SL g99 ( 
.A1(n_71),
.A2(n_97),
.B1(n_68),
.B2(n_89),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_90),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_87),
.Y(n_134)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_103),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_67),
.A2(n_51),
.B1(n_48),
.B2(n_45),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_106),
.A2(n_87),
.B1(n_94),
.B2(n_75),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_26),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_110),
.Y(n_129)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_113),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_112),
.A2(n_116),
.B1(n_123),
.B2(n_66),
.Y(n_127)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_117),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_78),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_118),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_120),
.Y(n_145)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_11),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_122),
.B(n_125),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_78),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_70),
.B(n_13),
.Y(n_125)
);

NAND2x1_ASAP7_75t_SL g126 ( 
.A(n_76),
.B(n_95),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_126),
.A2(n_66),
.B(n_83),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_139),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_128),
.A2(n_132),
.B(n_134),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_130),
.A2(n_128),
.B1(n_145),
.B2(n_119),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_107),
.A2(n_115),
.B1(n_124),
.B2(n_99),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_107),
.A2(n_90),
.B1(n_94),
.B2(n_75),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_148),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_143),
.B(n_100),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_126),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_105),
.B(n_5),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_149),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_SL g143 ( 
.A(n_108),
.B(n_5),
.C(n_72),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_99),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_72),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_165),
.B(n_144),
.Y(n_183)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_106),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_163),
.Y(n_181)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_157),
.B(n_167),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_101),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_161),
.B(n_164),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_132),
.A2(n_112),
.B1(n_116),
.B2(n_120),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_162),
.A2(n_166),
.B1(n_153),
.B2(n_150),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_118),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_104),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_83),
.B(n_117),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_117),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_142),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_169),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_127),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_163),
.A2(n_135),
.B1(n_144),
.B2(n_143),
.Y(n_172)
);

AO221x1_ASAP7_75t_L g191 ( 
.A1(n_172),
.A2(n_183),
.B1(n_170),
.B2(n_180),
.C(n_174),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_134),
.C(n_133),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_174),
.C(n_176),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_130),
.C(n_138),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_156),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_175),
.B(n_155),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_138),
.C(n_147),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_165),
.A2(n_159),
.B(n_151),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_184),
.Y(n_195)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_188),
.B(n_189),
.Y(n_198)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_177),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_190),
.B(n_192),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_191),
.A2(n_193),
.B(n_196),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_185),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_178),
.B(n_160),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_197),
.Y(n_205)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_173),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_202),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_183),
.C(n_176),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_195),
.C(n_197),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_181),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_178),
.Y(n_206)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_211),
.Y(n_214)
);

OAI32xp33_ASAP7_75t_L g208 ( 
.A1(n_198),
.A2(n_182),
.A3(n_150),
.B1(n_189),
.B2(n_193),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_210),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_157),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_184),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_200),
.B(n_162),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_212),
.A2(n_203),
.B1(n_202),
.B2(n_201),
.Y(n_216)
);

BUFx24_ASAP7_75t_SL g215 ( 
.A(n_209),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_216),
.Y(n_220)
);

INVxp33_ASAP7_75t_L g218 ( 
.A(n_213),
.Y(n_218)
);

A2O1A1Ixp33_ASAP7_75t_SL g222 ( 
.A1(n_218),
.A2(n_166),
.B(n_196),
.C(n_152),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_214),
.B(n_209),
.Y(n_219)
);

MAJx2_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_221),
.C(n_154),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_212),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_222),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_220),
.C(n_218),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_223),
.Y(n_226)
);


endmodule