module fake_jpeg_15067_n_263 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_263);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_263;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_30),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_25),
.B1(n_18),
.B2(n_13),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_35),
.A2(n_25),
.B1(n_34),
.B2(n_30),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_25),
.B1(n_18),
.B2(n_21),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_42),
.B1(n_18),
.B2(n_25),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_44),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_18),
.B1(n_25),
.B2(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_13),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_13),
.Y(n_58)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_51),
.Y(n_69)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_61),
.B1(n_38),
.B2(n_30),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_46),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_64),
.B1(n_38),
.B2(n_36),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_58),
.B(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_13),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_14),
.Y(n_81)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_14),
.Y(n_62)
);

NAND3xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_19),
.C(n_15),
.Y(n_79)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_23),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_40),
.C(n_42),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_65),
.B(n_75),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

NAND2x1_ASAP7_75t_SL g71 ( 
.A(n_51),
.B(n_37),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_64),
.B(n_58),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_27),
.C(n_31),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_81),
.B1(n_82),
.B2(n_64),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_78),
.B(n_79),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_27),
.C(n_28),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_85),
.Y(n_103)
);

MAJx2_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_54),
.C(n_62),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_89),
.B(n_94),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_72),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_87),
.B(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_64),
.B(n_49),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_49),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_97),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_57),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_66),
.A2(n_48),
.B1(n_56),
.B2(n_57),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_98),
.A2(n_61),
.B1(n_38),
.B2(n_55),
.Y(n_111)
);

MAJx2_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_48),
.C(n_53),
.Y(n_99)
);

AOI322xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_81),
.A3(n_50),
.B1(n_63),
.B2(n_76),
.C1(n_72),
.C2(n_79),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_66),
.B1(n_77),
.B2(n_71),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_109),
.B1(n_111),
.B2(n_113),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_85),
.Y(n_102)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_61),
.B1(n_70),
.B2(n_53),
.Y(n_104)
);

OAI22x1_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_80),
.B1(n_63),
.B2(n_70),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_92),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_119),
.B(n_14),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_86),
.A2(n_98),
.B1(n_94),
.B2(n_88),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_74),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_115),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_99),
.A2(n_81),
.B1(n_78),
.B2(n_76),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_74),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_102),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_127),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_122),
.A2(n_139),
.B1(n_52),
.B2(n_125),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_110),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_126),
.B(n_137),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_108),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_88),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_132),
.C(n_133),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_99),
.B(n_81),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_129),
.Y(n_153)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_84),
.B1(n_89),
.B2(n_93),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_131),
.A2(n_134),
.B1(n_124),
.B2(n_121),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_84),
.C(n_93),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_29),
.C(n_28),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_111),
.A2(n_103),
.B1(n_109),
.B2(n_101),
.Y(n_134)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_63),
.B(n_55),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_141),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_119),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_108),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_23),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_114),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_113),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_156),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_103),
.B1(n_102),
.B2(n_106),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_145),
.A2(n_158),
.B1(n_45),
.B2(n_23),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_146),
.B(n_157),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_107),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_151),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_107),
.Y(n_149)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_150),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_116),
.Y(n_151)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_104),
.Y(n_155)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_52),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_39),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_178)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_164),
.A2(n_24),
.B1(n_15),
.B2(n_19),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_153),
.A2(n_124),
.B1(n_132),
.B2(n_139),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_165),
.A2(n_172),
.B1(n_176),
.B2(n_177),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_131),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_174),
.C(n_175),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_152),
.A2(n_135),
.B1(n_136),
.B2(n_47),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_39),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_29),
.C(n_28),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_47),
.B1(n_45),
.B2(n_39),
.Y(n_176)
);

OAI21x1_ASAP7_75t_L g177 ( 
.A1(n_147),
.A2(n_12),
.B(n_11),
.Y(n_177)
);

NOR2xp67_ASAP7_75t_SL g179 ( 
.A(n_151),
.B(n_47),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_179),
.A2(n_12),
.B(n_11),
.Y(n_190)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_33),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_29),
.C(n_31),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_171),
.A2(n_158),
.B1(n_157),
.B2(n_149),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_184),
.B(n_198),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_181),
.A2(n_144),
.B1(n_145),
.B2(n_143),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_199),
.Y(n_205)
);

OAI22x1_ASAP7_75t_L g186 ( 
.A1(n_180),
.A2(n_142),
.B1(n_150),
.B2(n_156),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_168),
.B(n_146),
.Y(n_189)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_166),
.A2(n_24),
.B(n_19),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_197),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_33),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_175),
.C(n_176),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_165),
.A2(n_11),
.B(n_9),
.Y(n_195)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_24),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_196),
.Y(n_212)
);

FAx1_ASAP7_75t_SL g197 ( 
.A(n_170),
.B(n_33),
.CI(n_31),
.CON(n_197),
.SN(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_178),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_200),
.B(n_0),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_172),
.Y(n_203)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_199),
.C(n_200),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_174),
.C(n_170),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_207),
.C(n_197),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_167),
.C(n_15),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_213),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_9),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_9),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_0),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_217),
.C(n_218),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_194),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_197),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_186),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_219),
.B(n_222),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_185),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_204),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_192),
.C(n_22),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_226),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_22),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_225),
.B(n_20),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_201),
.A2(n_22),
.B(n_20),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_17),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_214),
.A2(n_22),
.B(n_20),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_228),
.A2(n_20),
.B(n_17),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_212),
.Y(n_230)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_230),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_208),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_0),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_232),
.B(n_234),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_225),
.Y(n_239)
);

AOI21x1_ASAP7_75t_L g235 ( 
.A1(n_222),
.A2(n_205),
.B(n_8),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_235),
.A2(n_219),
.B(n_17),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_1),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_239),
.Y(n_248)
);

FAx1_ASAP7_75t_SL g240 ( 
.A(n_238),
.B(n_218),
.CI(n_216),
.CON(n_240),
.SN(n_240)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_245),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_SL g249 ( 
.A1(n_242),
.A2(n_236),
.B(n_4),
.C(n_5),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_238),
.A2(n_17),
.B(n_8),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_3),
.B(n_4),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_16),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_247),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_249),
.Y(n_254)
);

MAJx2_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_253),
.C(n_3),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_3),
.B(n_4),
.Y(n_253)
);

A2O1A1O1Ixp25_ASAP7_75t_L g255 ( 
.A1(n_251),
.A2(n_240),
.B(n_241),
.C(n_239),
.D(n_6),
.Y(n_255)
);

OAI321xp33_ASAP7_75t_L g259 ( 
.A1(n_255),
.A2(n_256),
.A3(n_257),
.B1(n_3),
.B2(n_5),
.C(n_6),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g256 ( 
.A(n_252),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_254),
.A2(n_248),
.B(n_4),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_258),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_260),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_259),
.Y(n_262)
);

OAI321xp33_ASAP7_75t_L g263 ( 
.A1(n_262),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_16),
.C(n_258),
.Y(n_263)
);


endmodule