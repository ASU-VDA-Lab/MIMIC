module fake_jpeg_30340_n_493 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_493);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_493;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_2),
.B(n_3),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_15),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_31),
.Y(n_51)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_51),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_53),
.B(n_70),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_57),
.Y(n_137)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_62),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_63),
.Y(n_148)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_65),
.Y(n_150)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_68),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_16),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_74),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_35),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_35),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_75),
.B(n_76),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_35),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_78),
.B(n_83),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_16),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_91),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_35),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_39),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_87),
.B(n_89),
.Y(n_154)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

OR2x2_ASAP7_75t_SL g89 ( 
.A(n_47),
.B(n_15),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_15),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_18),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_95),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_99),
.Y(n_143)
);

CKINVDCx9p33_ASAP7_75t_R g104 ( 
.A(n_56),
.Y(n_104)
);

INVx3_ASAP7_75t_SL g172 ( 
.A(n_104),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_95),
.A2(n_40),
.B1(n_41),
.B2(n_44),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_112),
.A2(n_119),
.B1(n_20),
.B2(n_38),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_89),
.B(n_29),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_115),
.B(n_132),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_52),
.A2(n_18),
.B1(n_44),
.B2(n_32),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_29),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_145),
.Y(n_158)
);

BUFx6f_ASAP7_75t_SL g127 ( 
.A(n_51),
.Y(n_127)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_127),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_79),
.B(n_19),
.Y(n_132)
);

BUFx24_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_133),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_50),
.A2(n_40),
.B1(n_43),
.B2(n_19),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_20),
.Y(n_169)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_55),
.Y(n_142)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_66),
.B(n_30),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_54),
.Y(n_149)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_96),
.B(n_30),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_28),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_111),
.B(n_92),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_159),
.B(n_163),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_160),
.B(n_169),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_162),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_38),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_165),
.B(n_176),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_101),
.Y(n_166)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_79),
.B(n_93),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_168),
.A2(n_143),
.B(n_103),
.Y(n_252)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

INVx13_ASAP7_75t_L g233 ( 
.A(n_170),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_107),
.Y(n_173)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_173),
.Y(n_219)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_175),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_129),
.B(n_80),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_109),
.B(n_28),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_177),
.B(n_187),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_141),
.A2(n_84),
.B1(n_32),
.B2(n_27),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_179),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_122),
.Y(n_180)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_180),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_141),
.A2(n_27),
.B1(n_24),
.B2(n_41),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_183),
.Y(n_222)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_184),
.Y(n_230)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_108),
.Y(n_186)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_186),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_43),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_117),
.Y(n_188)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_188),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_135),
.A2(n_65),
.B1(n_85),
.B2(n_81),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_189),
.A2(n_190),
.B1(n_197),
.B2(n_199),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_135),
.A2(n_63),
.B1(n_77),
.B2(n_73),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_105),
.B(n_34),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_191),
.B(n_194),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_112),
.A2(n_22),
.B1(n_24),
.B2(n_34),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_192),
.A2(n_193),
.B1(n_212),
.B2(n_153),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_120),
.A2(n_18),
.B1(n_62),
.B2(n_69),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_125),
.B(n_99),
.Y(n_194)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_108),
.Y(n_195)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_195),
.Y(n_254)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_110),
.Y(n_196)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_138),
.A2(n_68),
.B1(n_57),
.B2(n_18),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_123),
.B(n_18),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_198),
.B(n_204),
.Y(n_246)
);

AO22x1_ASAP7_75t_SL g199 ( 
.A1(n_100),
.A2(n_97),
.B1(n_25),
.B2(n_23),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_107),
.Y(n_200)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

NAND2xp33_ASAP7_75t_SL g202 ( 
.A(n_133),
.B(n_23),
.Y(n_202)
);

AND2x2_ASAP7_75t_SL g255 ( 
.A(n_202),
.B(n_124),
.Y(n_255)
);

OA22x2_ASAP7_75t_L g203 ( 
.A1(n_119),
.A2(n_25),
.B1(n_23),
.B2(n_3),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_203),
.A2(n_113),
.B1(n_25),
.B2(n_155),
.Y(n_224)
);

AOI21xp33_ASAP7_75t_L g204 ( 
.A1(n_133),
.A2(n_25),
.B(n_23),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_106),
.Y(n_205)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_136),
.Y(n_206)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_206),
.Y(n_245)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_114),
.Y(n_207)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_207),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_131),
.B(n_0),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_208),
.Y(n_218)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_128),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_209),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_126),
.B(n_1),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_211),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_102),
.A2(n_25),
.B1(n_23),
.B2(n_5),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_158),
.B(n_139),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_223),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_138),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_224),
.A2(n_172),
.B1(n_180),
.B2(n_162),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_176),
.B(n_137),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_231),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_176),
.B(n_137),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_169),
.B(n_147),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_242),
.B(n_244),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_168),
.A2(n_102),
.B1(n_136),
.B2(n_155),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_243),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_203),
.B(n_153),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_210),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_172),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_251),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_252),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_203),
.A2(n_150),
.B1(n_148),
.B2(n_147),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_173),
.B1(n_200),
.B2(n_195),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_255),
.Y(n_267)
);

AND2x6_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_152),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_259),
.B(n_268),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_214),
.A2(n_171),
.B(n_202),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_261),
.A2(n_216),
.B(n_227),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_213),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_262),
.B(n_265),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_263),
.A2(n_277),
.B1(n_286),
.B2(n_288),
.Y(n_302)
);

OAI22x1_ASAP7_75t_L g266 ( 
.A1(n_214),
.A2(n_203),
.B1(n_199),
.B2(n_186),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_266),
.A2(n_235),
.B1(n_245),
.B2(n_254),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_181),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_270),
.A2(n_296),
.B1(n_245),
.B2(n_228),
.Y(n_299)
);

AOI21xp33_ASAP7_75t_L g271 ( 
.A1(n_242),
.A2(n_174),
.B(n_161),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_271),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_244),
.A2(n_206),
.B1(n_118),
.B2(n_148),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_272),
.A2(n_274),
.B1(n_276),
.B2(n_239),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_248),
.A2(n_118),
.B1(n_150),
.B2(n_199),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_255),
.Y(n_275)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_275),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_248),
.A2(n_205),
.B1(n_209),
.B2(n_207),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_223),
.A2(n_184),
.B1(n_179),
.B2(n_143),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_218),
.B(n_201),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_278),
.B(n_285),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_215),
.B(n_188),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_279),
.B(n_287),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_185),
.C(n_167),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_295),
.Y(n_314)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_220),
.Y(n_281)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_281),
.Y(n_332)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_220),
.Y(n_282)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_282),
.Y(n_310)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_227),
.Y(n_283)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_283),
.Y(n_311)
);

INVx4_ASAP7_75t_SL g284 ( 
.A(n_229),
.Y(n_284)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_284),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_218),
.B(n_171),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_217),
.A2(n_238),
.B1(n_252),
.B2(n_257),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_213),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_217),
.A2(n_175),
.B1(n_170),
.B2(n_164),
.Y(n_288)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_229),
.Y(n_289)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_289),
.Y(n_323)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_230),
.Y(n_290)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_290),
.Y(n_325)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_230),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_291),
.A2(n_292),
.B1(n_219),
.B2(n_236),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_219),
.Y(n_292)
);

NAND3xp33_ASAP7_75t_L g294 ( 
.A(n_256),
.B(n_1),
.C(n_4),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_294),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_238),
.B(n_116),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_238),
.A2(n_234),
.B1(n_226),
.B2(n_231),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_221),
.B(n_164),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_298),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_237),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_299),
.B(n_306),
.Y(n_348)
);

INVx13_ASAP7_75t_L g346 ( 
.A(n_301),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_305),
.A2(n_330),
.B(n_262),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_293),
.A2(n_234),
.B1(n_222),
.B2(n_235),
.Y(n_306)
);

AO21x1_ASAP7_75t_L g345 ( 
.A1(n_308),
.A2(n_319),
.B(n_284),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_266),
.A2(n_236),
.B1(n_222),
.B2(n_254),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_309),
.A2(n_312),
.B1(n_321),
.B2(n_326),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_260),
.A2(n_258),
.B1(n_273),
.B2(n_296),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_273),
.A2(n_228),
.B1(n_250),
.B2(n_241),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_316),
.B(n_318),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_250),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_317),
.B(n_10),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_260),
.A2(n_241),
.B1(n_247),
.B2(n_216),
.Y(n_318)
);

NOR2x1_ASAP7_75t_SL g319 ( 
.A(n_258),
.B(n_233),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_279),
.B(n_239),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_320),
.B(n_335),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_267),
.A2(n_225),
.B1(n_249),
.B2(n_237),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_324),
.A2(n_328),
.B1(n_333),
.B2(n_334),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_269),
.A2(n_232),
.B1(n_225),
.B2(n_249),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_269),
.A2(n_232),
.B1(n_116),
.B2(n_233),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_267),
.A2(n_1),
.B(n_4),
.Y(n_330)
);

AND2x2_ASAP7_75t_SL g331 ( 
.A(n_264),
.B(n_1),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_331),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_270),
.A2(n_210),
.B1(n_6),
.B2(n_7),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_275),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_264),
.B(n_4),
.Y(n_335)
);

AOI32xp33_ASAP7_75t_L g336 ( 
.A1(n_329),
.A2(n_259),
.A3(n_261),
.B1(n_280),
.B2(n_263),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_336),
.A2(n_347),
.B(n_327),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_306),
.B(n_289),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_337),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_315),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_338),
.Y(n_374)
);

MAJx2_ASAP7_75t_L g340 ( 
.A(n_314),
.B(n_283),
.C(n_277),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_340),
.B(n_366),
.Y(n_389)
);

OAI21xp33_ASAP7_75t_L g342 ( 
.A1(n_313),
.A2(n_288),
.B(n_287),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_342),
.A2(n_325),
.B1(n_332),
.B2(n_13),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_315),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_343),
.Y(n_393)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_304),
.Y(n_344)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_344),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_345),
.A2(n_308),
.B(n_318),
.Y(n_370)
);

INVx13_ASAP7_75t_L g349 ( 
.A(n_319),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_356),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_302),
.A2(n_284),
.B1(n_292),
.B2(n_290),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_350),
.A2(n_352),
.B1(n_362),
.B2(n_323),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_307),
.B(n_291),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_351),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_302),
.A2(n_292),
.B1(n_282),
.B2(n_281),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_304),
.Y(n_354)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_354),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_314),
.B(n_210),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_355),
.B(n_317),
.C(n_300),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_303),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_311),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_357),
.B(n_358),
.Y(n_382)
);

NAND3xp33_ASAP7_75t_L g358 ( 
.A(n_322),
.B(n_7),
.C(n_8),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_311),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_359),
.B(n_363),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_312),
.A2(n_210),
.B1(n_10),
.B2(n_11),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_320),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_307),
.B(n_7),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_364),
.B(n_334),
.Y(n_378)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_303),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_365),
.B(n_367),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_335),
.B(n_11),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_370),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_347),
.A2(n_300),
.B(n_313),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_371),
.A2(n_372),
.B(n_392),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_344),
.A2(n_309),
.B1(n_299),
.B2(n_331),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_373),
.A2(n_387),
.B1(n_353),
.B2(n_350),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_375),
.B(n_379),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_356),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_376),
.B(n_385),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_316),
.C(n_331),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_377),
.B(n_352),
.C(n_362),
.Y(n_417)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_378),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_340),
.B(n_330),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_365),
.A2(n_326),
.B1(n_328),
.B2(n_333),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_383),
.A2(n_384),
.B1(n_394),
.B2(n_348),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_384),
.A2(n_394),
.B1(n_359),
.B2(n_360),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_357),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_348),
.A2(n_323),
.B1(n_331),
.B2(n_322),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_354),
.B(n_310),
.Y(n_388)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_388),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_361),
.B(n_310),
.Y(n_391)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_391),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_345),
.A2(n_325),
.B(n_332),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_375),
.B(n_345),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_399),
.B(n_400),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_375),
.B(n_366),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_373),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_401),
.B(n_407),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_389),
.B(n_361),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_404),
.B(n_377),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_376),
.B(n_363),
.Y(n_405)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_405),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_406),
.B(n_417),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_382),
.B(n_367),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_382),
.B(n_339),
.Y(n_408)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_408),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_410),
.A2(n_414),
.B1(n_415),
.B2(n_416),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_389),
.B(n_336),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_412),
.B(n_396),
.Y(n_437)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_368),
.Y(n_413)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_413),
.Y(n_436)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_368),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_383),
.A2(n_360),
.B1(n_339),
.B2(n_349),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_390),
.B(n_341),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_418),
.B(n_383),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_419),
.B(n_437),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_397),
.B(n_372),
.C(n_377),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_421),
.B(n_425),
.C(n_396),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_397),
.B(n_371),
.C(n_388),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_426),
.B(n_432),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_399),
.B(n_379),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_428),
.B(n_430),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_400),
.B(n_379),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_429),
.B(n_431),
.Y(n_441)
);

MAJx2_ASAP7_75t_L g430 ( 
.A(n_412),
.B(n_390),
.C(n_381),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_398),
.A2(n_341),
.B1(n_369),
.B2(n_380),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_410),
.A2(n_380),
.B1(n_381),
.B2(n_395),
.Y(n_432)
);

OAI21xp33_ASAP7_75t_L g434 ( 
.A1(n_405),
.A2(n_386),
.B(n_391),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_434),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_404),
.B(n_387),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_435),
.B(n_417),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_438),
.B(n_422),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_439),
.B(n_425),
.C(n_437),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_420),
.B(n_406),
.C(n_402),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_443),
.B(n_447),
.C(n_449),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_427),
.A2(n_409),
.B1(n_415),
.B2(n_385),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_448),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_433),
.B(n_418),
.Y(n_446)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_446),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_420),
.B(n_411),
.C(n_374),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_436),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_422),
.B(n_411),
.C(n_393),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_428),
.B(n_370),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_430),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_421),
.A2(n_403),
.B(n_392),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_451),
.A2(n_403),
.B(n_386),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_460),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_445),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_455),
.B(n_456),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_447),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_458),
.B(n_465),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_459),
.B(n_463),
.Y(n_469)
);

NOR2xp67_ASAP7_75t_SL g460 ( 
.A(n_452),
.B(n_439),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_442),
.B(n_424),
.C(n_426),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_462),
.B(n_449),
.C(n_443),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_450),
.B(n_434),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_442),
.B(n_423),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_464),
.B(n_452),
.C(n_441),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_466),
.B(n_470),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_457),
.A2(n_461),
.B1(n_440),
.B2(n_458),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_472),
.B(n_473),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_453),
.B(n_448),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_453),
.B(n_378),
.Y(n_474)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_474),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_346),
.C(n_12),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_475),
.B(n_11),
.Y(n_476)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_476),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_468),
.A2(n_463),
.B1(n_459),
.B2(n_346),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_478),
.B(n_475),
.Y(n_483)
);

CKINVDCx14_ASAP7_75t_R g479 ( 
.A(n_467),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_479),
.A2(n_480),
.B1(n_477),
.B2(n_469),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_481),
.A2(n_471),
.B(n_472),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_482),
.B(n_483),
.C(n_479),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_484),
.B(n_469),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_486),
.A2(n_487),
.B1(n_485),
.B2(n_13),
.Y(n_488)
);

OAI21xp33_ASAP7_75t_SL g489 ( 
.A1(n_488),
.A2(n_12),
.B(n_14),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_489),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_490),
.B(n_12),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_491),
.B(n_14),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_492),
.B(n_14),
.Y(n_493)
);


endmodule