module real_jpeg_5496_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_0),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_SL g45 ( 
.A(n_0),
.B(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_0),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_0),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_0),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_0),
.B(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_0),
.Y(n_183)
);

AND2x2_ASAP7_75t_SL g216 ( 
.A(n_0),
.B(n_217),
.Y(n_216)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_2),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_2),
.B(n_28),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_2),
.B(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_2),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_2),
.B(n_414),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_2),
.B(n_420),
.Y(n_419)
);

NAND2x1_ASAP7_75t_SL g53 ( 
.A(n_3),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_3),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_3),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_3),
.B(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_3),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_3),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_3),
.B(n_132),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_3),
.B(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_4),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_4),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_4),
.Y(n_399)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g20 ( 
.A(n_6),
.B(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_6),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_6),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_6),
.B(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_SL g242 ( 
.A(n_6),
.B(n_243),
.Y(n_242)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_7),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_7),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_7),
.Y(n_243)
);

BUFx5_ASAP7_75t_L g425 ( 
.A(n_7),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_8),
.Y(n_106)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_8),
.Y(n_148)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_10),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_10),
.B(n_179),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_10),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_10),
.B(n_252),
.Y(n_251)
);

AND2x2_ASAP7_75t_SL g301 ( 
.A(n_10),
.B(n_95),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_10),
.B(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_10),
.B(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_10),
.B(n_402),
.Y(n_401)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_11),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_11),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_12),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_12),
.B(n_56),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_12),
.B(n_126),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_12),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_12),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_12),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_12),
.B(n_313),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_12),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_13),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_13),
.B(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_13),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_13),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_13),
.B(n_386),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_13),
.B(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_13),
.B(n_425),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_14),
.B(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_14),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_14),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_14),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_14),
.B(n_410),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_15),
.Y(n_169)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_15),
.Y(n_187)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

O2A1O1Ixp33_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_109),
.B(n_327),
.C(n_505),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_36),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_19),
.B(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_26),
.C(n_31),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_20),
.A2(n_31),
.B1(n_73),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_20),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_20),
.A2(n_86),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_20),
.B(n_228),
.Y(n_227)
);

NOR3xp33_ASAP7_75t_L g505 ( 
.A(n_20),
.B(n_45),
.C(n_103),
.Y(n_505)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_24),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_24),
.Y(n_219)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g353 ( 
.A(n_25),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_26),
.A2(n_27),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_26),
.A2(n_27),
.B1(n_333),
.B2(n_339),
.Y(n_332)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_27),
.B(n_334),
.C(n_338),
.Y(n_487)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_31),
.A2(n_41),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_31),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_31),
.A2(n_73),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_31),
.B(n_153),
.C(n_158),
.Y(n_256)
);

OR2x2_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_35),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_33),
.Y(n_278)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_34),
.Y(n_180)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_34),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_34),
.Y(n_336)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_34),
.Y(n_383)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_42),
.Y(n_41)
);

OR2x2_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_35),
.B(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_97),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_81),
.C(n_82),
.Y(n_37)
);

FAx1_ASAP7_75t_SL g502 ( 
.A(n_38),
.B(n_81),
.CI(n_82),
.CON(n_502),
.SN(n_502)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_62),
.C(n_70),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_39),
.B(n_493),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_52),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_40),
.B(n_57),
.C(n_60),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.C(n_48),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_41),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_41),
.B(n_73),
.C(n_80),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_41),
.A2(n_74),
.B1(n_120),
.B2(n_124),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_41),
.B(n_120),
.C(n_125),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_41),
.A2(n_74),
.B1(n_482),
.B2(n_483),
.Y(n_481)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_43),
.Y(n_217)
);

INVx5_ASAP7_75t_L g378 ( 
.A(n_43),
.Y(n_378)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_44),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_44),
.Y(n_255)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_44),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_45),
.A2(n_100),
.B1(n_101),
.B2(n_107),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_45),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_45),
.A2(n_48),
.B1(n_49),
.B2(n_107),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_46),
.Y(n_328)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_47),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_48),
.A2(n_49),
.B1(n_135),
.B2(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_48),
.A2(n_49),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_49),
.B(n_131),
.C(n_135),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_49),
.B(n_194),
.C(n_327),
.Y(n_486)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_56),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_57),
.Y(n_61)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_59),
.B(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_62),
.B(n_70),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.C(n_69),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_63),
.A2(n_66),
.B1(n_67),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_63),
.Y(n_477)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_66),
.A2(n_67),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_67),
.B(n_140),
.C(n_242),
.Y(n_316)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_69),
.B(n_476),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_75),
.B2(n_80),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_75),
.A2(n_80),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_79),
.Y(n_206)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_79),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_80),
.B(n_194),
.C(n_297),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_87),
.B1(n_88),
.B2(n_96),
.Y(n_82)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_86),
.B(n_229),
.C(n_234),
.Y(n_292)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_91),
.C(n_96),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_108),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_102),
.A2(n_103),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_102),
.A2(n_103),
.B1(n_351),
.B2(n_354),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_102),
.B(n_347),
.C(n_354),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_103),
.B(n_312),
.C(n_316),
.Y(n_345)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_105),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_501),
.B(n_504),
.Y(n_109)
);

AOI21x1_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_469),
.B(n_498),
.Y(n_110)
);

AO21x1_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_319),
.B(n_355),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_286),
.B(n_318),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_257),
.B(n_285),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_114),
.B(n_467),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_221),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_115),
.B(n_221),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_173),
.C(n_207),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_116),
.B(n_284),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_149),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_117),
.B(n_150),
.C(n_160),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_130),
.C(n_138),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_118),
.B(n_281),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_125),
.Y(n_118)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_129),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_130),
.A2(n_138),
.B1(n_139),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_130),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_131),
.B(n_265),
.Y(n_264)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_134),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_135),
.Y(n_266)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_145),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_140),
.A2(n_241),
.B1(n_242),
.B2(n_244),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_140),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_140),
.A2(n_145),
.B1(n_146),
.B2(n_244),
.Y(n_279)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_143),
.Y(n_422)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_144),
.Y(n_214)
);

BUFx8_ASAP7_75t_L g366 ( 
.A(n_144),
.Y(n_366)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_160),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_157),
.B2(n_158),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_154),
.B(n_194),
.Y(n_372)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_156),
.Y(n_202)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_156),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx24_ASAP7_75t_SL g509 ( 
.A(n_160),
.Y(n_509)
);

FAx1_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.CI(n_170),
.CON(n_160),
.SN(n_160)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_162),
.B(n_163),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_161),
.B(n_165),
.C(n_170),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_171),
.B(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_173),
.B(n_207),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_189),
.C(n_191),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_174),
.A2(n_189),
.B1(n_190),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_174),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_178),
.C(n_182),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_176),
.B(n_429),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_176),
.B(n_415),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_181),
.B1(n_182),
.B2(n_188),
.Y(n_177)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_181),
.A2(n_182),
.B1(n_300),
.B2(n_303),
.Y(n_299)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_182),
.B(n_242),
.C(n_301),
.Y(n_348)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_186),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g371 ( 
.A(n_187),
.Y(n_371)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_191),
.B(n_261),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_198),
.C(n_203),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_192),
.A2(n_193),
.B1(n_456),
.B2(n_457),
.Y(n_455)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_194),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_194),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_194),
.A2(n_294),
.B1(n_327),
.B2(n_329),
.Y(n_326)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_198),
.A2(n_199),
.B1(n_203),
.B2(n_204),
.Y(n_457)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_201),
.Y(n_402)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_220),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_210),
.C(n_220),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_215),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_216),
.C(n_218),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_216),
.A2(n_334),
.B1(n_337),
.B2(n_338),
.Y(n_333)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_216),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_222),
.B(n_224),
.C(n_245),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_245),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_238),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_226),
.B(n_227),
.C(n_238),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_234),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_241),
.A2(n_242),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_241),
.A2(n_242),
.B1(n_363),
.B2(n_364),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_242),
.B(n_363),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_246),
.B(n_248),
.C(n_249),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_256),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_251),
.B(n_253),
.C(n_308),
.Y(n_307)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_256),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_283),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_258),
.B(n_283),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_263),
.C(n_280),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_259),
.A2(n_260),
.B1(n_461),
.B2(n_462),
.Y(n_460)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_263),
.B(n_280),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_267),
.C(n_279),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_264),
.B(n_451),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_267),
.B(n_279),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_271),
.C(n_274),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_268),
.A2(n_269),
.B1(n_274),
.B2(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_271),
.B(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_274),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_275),
.B(n_376),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_275),
.B(n_432),
.Y(n_431)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx8_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_287),
.B(n_319),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_288),
.B(n_289),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_289),
.B(n_320),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_289),
.B(n_320),
.Y(n_468)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_304),
.CI(n_317),
.CON(n_289),
.SN(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_299),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_292),
.B(n_293),
.C(n_299),
.Y(n_342)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_300),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_301),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_307),
.C(n_309),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_309),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_316),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_321),
.B(n_323),
.C(n_340),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_340),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_330),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_324),
.B(n_331),
.C(n_332),
.Y(n_478)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_327),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_333),
.Y(n_339)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_334),
.Y(n_337)
);

INVx6_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_342),
.B1(n_343),
.B2(n_344),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_341),
.B(n_345),
.C(n_346),
.Y(n_488)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

AO22x1_ASAP7_75t_SL g346 ( 
.A1(n_347),
.A2(n_348),
.B1(n_349),
.B2(n_350),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_351),
.Y(n_354)
);

INVx5_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

OAI31xp33_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_465),
.A3(n_466),
.B(n_468),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_459),
.B(n_464),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_358),
.A2(n_446),
.B(n_458),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_404),
.B(n_445),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_390),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_360),
.B(n_390),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_373),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_361),
.B(n_374),
.C(n_387),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_367),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_362),
.B(n_368),
.C(n_372),
.Y(n_454)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_372),
.Y(n_367)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx8_ASAP7_75t_L g386 ( 
.A(n_371),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_387),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_379),
.C(n_384),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_375),
.B(n_392),
.Y(n_391)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_379),
.A2(n_380),
.B1(n_384),
.B2(n_385),
.Y(n_392)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx6_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_393),
.C(n_403),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_391),
.B(n_442),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_393),
.A2(n_394),
.B1(n_403),
.B2(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_400),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_395),
.A2(n_396),
.B1(n_400),
.B2(n_401),
.Y(n_416)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_399),
.Y(n_430)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_403),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_439),
.B(n_444),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_426),
.B(n_438),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_407),
.B(n_417),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_407),
.B(n_417),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_416),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_413),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_409),
.B(n_413),
.C(n_416),
.Y(n_440)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_423),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_418),
.A2(n_419),
.B1(n_423),
.B2(n_424),
.Y(n_436)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_434),
.B(n_437),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_431),
.Y(n_427)
);

INVx5_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_436),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_435),
.B(n_436),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_441),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_440),
.B(n_441),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_447),
.B(n_448),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_449),
.A2(n_450),
.B1(n_452),
.B2(n_453),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_449),
.B(n_454),
.C(n_455),
.Y(n_463)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_455),
.Y(n_453)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_463),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_460),
.B(n_463),
.Y(n_464)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_461),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_494),
.Y(n_469)
);

OAI21xp33_ASAP7_75t_L g498 ( 
.A1(n_470),
.A2(n_499),
.B(n_500),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_489),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_471),
.B(n_489),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_479),
.C(n_488),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_472),
.B(n_479),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_473),
.B(n_478),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_475),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_474),
.B(n_475),
.C(n_478),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_480),
.A2(n_481),
.B1(n_484),
.B2(n_485),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_480),
.B(n_486),
.C(n_487),
.Y(n_491)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_487),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_488),
.B(n_497),
.Y(n_496)
);

BUFx24_ASAP7_75t_SL g507 ( 
.A(n_489),
.Y(n_507)
);

FAx1_ASAP7_75t_SL g489 ( 
.A(n_490),
.B(n_491),
.CI(n_492),
.CON(n_489),
.SN(n_489)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_490),
.B(n_491),
.C(n_492),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_496),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_495),
.B(n_496),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_503),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_502),
.B(n_503),
.Y(n_504)
);

BUFx24_ASAP7_75t_SL g508 ( 
.A(n_502),
.Y(n_508)
);


endmodule