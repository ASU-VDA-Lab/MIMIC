module fake_jpeg_5292_n_139 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_25),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_16),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_28),
.B(n_20),
.Y(n_44)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

NOR2x1_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_36),
.B1(n_43),
.B2(n_27),
.Y(n_45)
);

AO22x2_ASAP7_75t_SL g36 ( 
.A1(n_30),
.A2(n_14),
.B1(n_22),
.B2(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_44),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_11),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_16),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_49),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_25),
.C(n_24),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_52),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_18),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_21),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_34),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_L g58 ( 
.A1(n_54),
.A2(n_55),
.B(n_24),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_20),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_64),
.B(n_46),
.Y(n_78)
);

AO22x1_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_41),
.B1(n_43),
.B2(n_24),
.Y(n_59)
);

A2O1A1O1Ixp25_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_48),
.B(n_53),
.C(n_22),
.D(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_15),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_60),
.B(n_65),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_63),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_53),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g64 ( 
.A1(n_51),
.A2(n_32),
.B(n_13),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_29),
.B1(n_41),
.B2(n_31),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_38),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_35),
.B(n_17),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_46),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_73),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_65),
.B(n_51),
.Y(n_73)
);

NOR3xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_60),
.C(n_12),
.Y(n_94)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_76),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_78),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_15),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_68),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_83),
.B(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_62),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_91),
.B(n_13),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_67),
.C(n_66),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_70),
.C(n_57),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_78),
.C(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

NOR3xp33_ASAP7_75t_SL g96 ( 
.A(n_89),
.B(n_74),
.C(n_73),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_96),
.A2(n_83),
.B(n_92),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_86),
.A2(n_70),
.B1(n_80),
.B2(n_29),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_101),
.B1(n_84),
.B2(n_88),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_104),
.C(n_105),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

AO221x1_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_61),
.B1(n_56),
.B2(n_50),
.C(n_57),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_0),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_93),
.A2(n_31),
.B1(n_35),
.B2(n_40),
.Y(n_101)
);

OAI322xp33_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_12),
.A3(n_26),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_26),
.C(n_40),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_2),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_107),
.B(n_10),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_103),
.A2(n_56),
.B1(n_50),
.B2(n_31),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_109),
.A2(n_110),
.B1(n_101),
.B2(n_99),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_98),
.A2(n_40),
.B1(n_1),
.B2(n_0),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_112),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_1),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_100),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_106),
.A2(n_96),
.B(n_97),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_108),
.B(n_111),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_117),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_105),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_3),
.C(n_5),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_3),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_120),
.A2(n_114),
.B1(n_107),
.B2(n_113),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_124),
.C(n_127),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_115),
.A2(n_112),
.B1(n_114),
.B2(n_6),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_125),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_131)
);

OAI221xp5_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_121),
.B1(n_122),
.B2(n_125),
.C(n_127),
.Y(n_129)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

AO21x1_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_118),
.B(n_7),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_130),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_131),
.A2(n_132),
.B1(n_8),
.B2(n_9),
.Y(n_135)
);

NOR2xp67_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_8),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_10),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_128),
.C(n_131),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_137),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_134),
.Y(n_139)
);


endmodule