module real_aes_7972_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_841;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_852;
wire n_857;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_320;
wire n_884;
wire n_537;
wire n_551;
wire n_560;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_462;
wire n_289;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_356;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_892;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_656;
wire n_316;
wire n_532;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_617;
wire n_552;
wire n_602;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_898;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_365;
wire n_290;
wire n_526;
wire n_899;
wire n_637;
wire n_692;
wire n_789;
wire n_544;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_888;
wire n_836;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g509 ( .A1(n_0), .A2(n_253), .B1(n_510), .B2(n_511), .Y(n_509) );
AOI22xp33_ASAP7_75t_SL g512 ( .A1(n_1), .A2(n_126), .B1(n_513), .B2(n_516), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_2), .A2(n_104), .B1(n_405), .B2(n_525), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_3), .B(n_365), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_4), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_5), .A2(n_28), .B1(n_473), .B2(n_474), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_6), .A2(n_221), .B1(n_647), .B2(n_725), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g894 ( .A(n_7), .Y(n_894) );
AOI22xp33_ASAP7_75t_SL g590 ( .A1(n_8), .A2(n_114), .B1(n_384), .B2(n_436), .Y(n_590) );
OA22x2_ASAP7_75t_L g717 ( .A1(n_9), .A2(n_718), .B1(n_719), .B2(n_743), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_9), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_10), .A2(n_184), .B1(n_405), .B2(n_406), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_11), .A2(n_187), .B1(n_631), .B2(n_723), .Y(n_867) );
CKINVDCx20_ASAP7_75t_R g898 ( .A(n_12), .Y(n_898) );
AOI211xp5_ASAP7_75t_L g605 ( .A1(n_13), .A2(n_606), .B(n_607), .C(n_610), .Y(n_605) );
XOR2x2_ASAP7_75t_L g561 ( .A(n_14), .B(n_562), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_15), .A2(n_144), .B1(n_463), .B2(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g903 ( .A(n_16), .Y(n_903) );
CKINVDCx20_ASAP7_75t_R g667 ( .A(n_17), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_18), .A2(n_31), .B1(n_552), .B2(n_553), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_19), .A2(n_199), .B1(n_340), .B2(n_407), .Y(n_564) );
AOI22xp33_ASAP7_75t_SL g592 ( .A1(n_20), .A2(n_277), .B1(n_593), .B2(n_594), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_21), .Y(n_542) );
AOI22xp33_ASAP7_75t_SL g518 ( .A1(n_22), .A2(n_233), .B1(n_519), .B2(n_520), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_23), .Y(n_696) );
AOI22xp33_ASAP7_75t_SL g616 ( .A1(n_24), .A2(n_156), .B1(n_457), .B2(n_617), .Y(n_616) );
AOI22xp33_ASAP7_75t_SL g708 ( .A1(n_25), .A2(n_138), .B1(n_414), .B2(n_631), .Y(n_708) );
OA22x2_ASAP7_75t_L g533 ( .A1(n_26), .A2(n_534), .B1(n_535), .B2(n_559), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_26), .Y(n_534) );
AOI22xp33_ASAP7_75t_SL g705 ( .A1(n_27), .A2(n_206), .B1(n_457), .B2(n_680), .Y(n_705) );
AOI22xp33_ASAP7_75t_SL g722 ( .A1(n_29), .A2(n_249), .B1(n_603), .B2(n_723), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_30), .A2(n_245), .B1(n_520), .B2(n_556), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_32), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g891 ( .A(n_33), .Y(n_891) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_34), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_35), .A2(n_48), .B1(n_413), .B2(n_553), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_36), .A2(n_278), .B1(n_467), .B2(n_501), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_37), .A2(n_194), .B1(n_510), .B2(n_522), .Y(n_645) );
CKINVDCx20_ASAP7_75t_R g884 ( .A(n_38), .Y(n_884) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_39), .Y(n_776) );
AO22x2_ASAP7_75t_L g316 ( .A1(n_40), .A2(n_98), .B1(n_308), .B2(n_313), .Y(n_316) );
INVx1_ASAP7_75t_L g836 ( .A(n_40), .Y(n_836) );
AOI221xp5_ASAP7_75t_L g339 ( .A1(n_41), .A2(n_252), .B1(n_340), .B2(n_344), .C(n_349), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_42), .A2(n_46), .B1(n_390), .B2(n_594), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_43), .Y(n_811) );
AOI222xp33_ASAP7_75t_L g380 ( .A1(n_44), .A2(n_121), .B1(n_176), .B2(n_381), .C1(n_384), .C2(n_389), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_45), .A2(n_115), .B1(n_344), .B2(n_405), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g333 ( .A(n_47), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_49), .A2(n_50), .B1(n_650), .B2(n_742), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_51), .A2(n_397), .B1(n_443), .B2(n_444), .Y(n_396) );
INVx1_ASAP7_75t_L g443 ( .A(n_51), .Y(n_443) );
AOI222xp33_ASAP7_75t_L g475 ( .A1(n_52), .A2(n_146), .B1(n_212), .B2(n_476), .C1(n_477), .C2(n_479), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_53), .A2(n_279), .B1(n_465), .B2(n_627), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_54), .A2(n_70), .B1(n_477), .B2(n_479), .Y(n_799) );
AOI22xp33_ASAP7_75t_SL g729 ( .A1(n_55), .A2(n_139), .B1(n_513), .B2(n_730), .Y(n_729) );
AO22x2_ASAP7_75t_L g318 ( .A1(n_56), .A2(n_102), .B1(n_308), .B2(n_309), .Y(n_318) );
INVx1_ASAP7_75t_L g837 ( .A(n_56), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g881 ( .A1(n_57), .A2(n_142), .B1(n_391), .B2(n_468), .Y(n_881) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_58), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_59), .A2(n_78), .B1(n_467), .B2(n_653), .Y(n_652) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_60), .A2(n_287), .B(n_295), .C(n_838), .Y(n_286) );
AOI222xp33_ASAP7_75t_L g655 ( .A1(n_61), .A2(n_171), .B1(n_228), .B2(n_389), .C1(n_579), .C2(n_656), .Y(n_655) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_62), .Y(n_798) );
AOI22xp33_ASAP7_75t_SL g864 ( .A1(n_63), .A2(n_118), .B1(n_553), .B2(n_807), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_64), .A2(n_208), .B1(n_401), .B2(n_525), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_65), .B(n_435), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_66), .A2(n_285), .B1(n_335), .B2(n_526), .Y(n_618) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_67), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g367 ( .A(n_68), .Y(n_367) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_69), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_71), .A2(n_256), .B1(n_403), .B2(n_471), .Y(n_470) );
XNOR2xp5_ASAP7_75t_L g584 ( .A(n_72), .B(n_585), .Y(n_584) );
AOI22xp33_ASAP7_75t_SL g464 ( .A1(n_73), .A2(n_155), .B1(n_465), .B2(n_467), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_74), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_75), .A2(n_258), .B1(n_558), .B2(n_570), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_76), .Y(n_538) );
AOI22xp33_ASAP7_75t_SL g779 ( .A1(n_77), .A2(n_148), .B1(n_471), .B2(n_780), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_79), .A2(n_207), .B1(n_303), .B2(n_680), .Y(n_759) );
AOI221xp5_ASAP7_75t_L g300 ( .A1(n_80), .A2(n_159), .B1(n_301), .B2(n_319), .C(n_325), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_81), .B(n_463), .Y(n_754) );
INVx1_ASAP7_75t_L g580 ( .A(n_82), .Y(n_580) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_83), .A2(n_161), .B1(n_360), .B2(n_364), .C(n_366), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_84), .A2(n_179), .B1(n_335), .B2(n_410), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g781 ( .A1(n_85), .A2(n_131), .B1(n_414), .B2(n_567), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_86), .A2(n_236), .B1(n_410), .B2(n_558), .Y(n_557) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_87), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_88), .A2(n_172), .B1(n_346), .B2(n_617), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_89), .A2(n_273), .B1(n_385), .B2(n_391), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_90), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_91), .A2(n_299), .B1(n_393), .B2(n_394), .Y(n_298) );
INVx1_ASAP7_75t_L g393 ( .A(n_91), .Y(n_393) );
AOI22xp5_ASAP7_75t_SL g839 ( .A1(n_92), .A2(n_840), .B1(n_841), .B2(n_868), .Y(n_839) );
CKINVDCx20_ASAP7_75t_R g868 ( .A(n_92), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_93), .A2(n_224), .B1(n_468), .B2(n_576), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_94), .A2(n_175), .B1(n_413), .B2(n_417), .Y(n_412) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_95), .A2(n_145), .B1(n_335), .B2(n_572), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_96), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_97), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g887 ( .A(n_99), .Y(n_887) );
CKINVDCx20_ASAP7_75t_R g633 ( .A(n_100), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_101), .A2(n_149), .B1(n_401), .B2(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_SL g862 ( .A1(n_103), .A2(n_198), .B1(n_301), .B2(n_863), .Y(n_862) );
AOI22xp33_ASAP7_75t_SL g601 ( .A1(n_105), .A2(n_271), .B1(n_602), .B2(n_603), .Y(n_601) );
INVx1_ASAP7_75t_L g294 ( .A(n_106), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g674 ( .A(n_107), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_108), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_109), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_110), .A2(n_205), .B1(n_346), .B2(n_617), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_111), .A2(n_231), .B1(n_432), .B2(n_545), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_112), .A2(n_130), .B1(n_452), .B2(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g290 ( .A(n_113), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_116), .A2(n_158), .B1(n_390), .B2(n_478), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g851 ( .A(n_117), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_119), .B(n_516), .Y(n_609) );
CKINVDCx20_ASAP7_75t_R g373 ( .A(n_120), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_122), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g854 ( .A(n_123), .Y(n_854) );
INVx1_ASAP7_75t_L g883 ( .A(n_124), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_125), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_127), .A2(n_160), .B1(n_473), .B2(n_553), .Y(n_643) );
OA22x2_ASAP7_75t_L g764 ( .A1(n_128), .A2(n_765), .B1(n_766), .B2(n_767), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_128), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_129), .A2(n_151), .B1(n_385), .B2(n_465), .Y(n_702) );
AOI22xp33_ASAP7_75t_SL g740 ( .A1(n_132), .A2(n_162), .B1(n_593), .B2(n_594), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_133), .A2(n_229), .B1(n_452), .B2(n_780), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_134), .A2(n_247), .B1(n_600), .B2(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_135), .A2(n_143), .B1(n_344), .B2(n_453), .Y(n_642) );
AOI22xp33_ASAP7_75t_SL g595 ( .A1(n_136), .A2(n_238), .B1(n_463), .B2(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_137), .A2(n_178), .B1(n_455), .B2(n_457), .Y(n_454) );
INVx1_ASAP7_75t_L g874 ( .A(n_140), .Y(n_874) );
AOI22xp33_ASAP7_75t_SL g747 ( .A1(n_141), .A2(n_234), .B1(n_342), .B2(n_515), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_147), .B(n_500), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_150), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_152), .A2(n_230), .B1(n_522), .B2(n_525), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_153), .Y(n_505) );
XNOR2x2_ASAP7_75t_L g639 ( .A(n_154), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g293 ( .A(n_157), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g710 ( .A(n_163), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_164), .B(n_579), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_165), .B(n_365), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_166), .B(n_361), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_167), .A2(n_280), .B1(n_474), .B2(n_807), .Y(n_806) );
AND2x6_ASAP7_75t_L g289 ( .A(n_168), .B(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_168), .Y(n_830) );
AO22x2_ASAP7_75t_L g307 ( .A1(n_169), .A2(n_241), .B1(n_308), .B2(n_309), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_170), .A2(n_222), .B1(n_340), .B2(n_457), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g847 ( .A(n_173), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g671 ( .A(n_174), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_177), .A2(n_269), .B1(n_467), .B2(n_501), .Y(n_622) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_180), .Y(n_886) );
CKINVDCx20_ASAP7_75t_R g895 ( .A(n_181), .Y(n_895) );
CKINVDCx20_ASAP7_75t_R g350 ( .A(n_182), .Y(n_350) );
AOI22xp33_ASAP7_75t_SL g783 ( .A1(n_183), .A2(n_257), .B1(n_321), .B2(n_335), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_185), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_186), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_188), .A2(n_227), .B1(n_386), .B2(n_465), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_189), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_190), .B(n_700), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_191), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g326 ( .A(n_192), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_193), .A2(n_284), .B1(n_361), .B2(n_364), .Y(n_574) );
AO22x2_ASAP7_75t_L g312 ( .A1(n_195), .A2(n_259), .B1(n_308), .B2(n_313), .Y(n_312) );
AOI22xp33_ASAP7_75t_SL g784 ( .A1(n_196), .A2(n_202), .B1(n_570), .B2(n_599), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_197), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_200), .A2(n_282), .B1(n_303), .B2(n_473), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_201), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_203), .A2(n_237), .B1(n_303), .B2(n_519), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_204), .A2(n_270), .B1(n_566), .B2(n_567), .Y(n_565) );
INVx1_ASAP7_75t_L g880 ( .A(n_209), .Y(n_880) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_210), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_211), .A2(n_232), .B1(n_328), .B2(n_647), .Y(n_646) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_213), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g859 ( .A(n_214), .Y(n_859) );
CKINVDCx20_ASAP7_75t_R g608 ( .A(n_215), .Y(n_608) );
AOI22xp33_ASAP7_75t_SL g598 ( .A1(n_216), .A2(n_254), .B1(n_599), .B2(n_600), .Y(n_598) );
INVx1_ASAP7_75t_L g901 ( .A(n_217), .Y(n_901) );
AOI22xp33_ASAP7_75t_SL g629 ( .A1(n_218), .A2(n_281), .B1(n_630), .B2(n_631), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_219), .A2(n_255), .B1(n_401), .B2(n_403), .Y(n_400) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_220), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_223), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_225), .B(n_365), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g892 ( .A(n_226), .B(n_617), .Y(n_892) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_235), .Y(n_818) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_239), .Y(n_794) );
AOI22x1_ASAP7_75t_L g662 ( .A1(n_240), .A2(n_663), .B1(n_687), .B2(n_688), .Y(n_662) );
INVx1_ASAP7_75t_L g687 ( .A(n_240), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_241), .B(n_835), .Y(n_834) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_242), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g844 ( .A(n_243), .Y(n_844) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_244), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g621 ( .A(n_246), .Y(n_621) );
CKINVDCx20_ASAP7_75t_R g611 ( .A(n_248), .Y(n_611) );
AOI22xp33_ASAP7_75t_SL g758 ( .A1(n_250), .A2(n_283), .B1(n_330), .B2(n_524), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g899 ( .A(n_251), .Y(n_899) );
INVx1_ASAP7_75t_L g833 ( .A(n_259), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_260), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g857 ( .A(n_261), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_262), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_263), .B(n_478), .Y(n_855) );
OA22x2_ASAP7_75t_L g786 ( .A1(n_264), .A2(n_787), .B1(n_788), .B2(n_789), .Y(n_786) );
CKINVDCx16_ASAP7_75t_R g787 ( .A(n_264), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_265), .B(n_462), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_266), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g666 ( .A(n_267), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_268), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_272), .Y(n_430) );
INVx1_ASAP7_75t_L g308 ( .A(n_274), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_274), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_275), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_276), .Y(n_502) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_290), .Y(n_829) );
OAI21xp5_ASAP7_75t_L g872 ( .A1(n_291), .A2(n_828), .B(n_873), .Y(n_872) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_292), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_529), .B1(n_823), .B2(n_824), .C(n_825), .Y(n_295) );
INVx1_ASAP7_75t_L g823 ( .A(n_296), .Y(n_823) );
AOI22xp5_ASAP7_75t_SL g296 ( .A1(n_297), .A2(n_485), .B1(n_527), .B2(n_528), .Y(n_296) );
INVx1_ASAP7_75t_L g527 ( .A(n_297), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_395), .B1(n_483), .B2(n_484), .Y(n_297) );
INVx1_ASAP7_75t_L g483 ( .A(n_298), .Y(n_483) );
INVx1_ASAP7_75t_L g394 ( .A(n_299), .Y(n_394) );
AND4x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_339), .C(n_359), .D(n_380), .Y(n_299) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
BUFx3_ASAP7_75t_L g405 ( .A(n_303), .Y(n_405) );
BUFx3_ASAP7_75t_L g510 ( .A(n_303), .Y(n_510) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g456 ( .A(n_304), .Y(n_456) );
BUFx2_ASAP7_75t_SL g558 ( .A(n_304), .Y(n_558) );
BUFx2_ASAP7_75t_SL g606 ( .A(n_304), .Y(n_606) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_314), .Y(n_304) );
AND2x6_ASAP7_75t_L g330 ( .A(n_305), .B(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g342 ( .A(n_305), .B(n_343), .Y(n_342) );
AND2x6_ASAP7_75t_L g383 ( .A(n_305), .B(n_377), .Y(n_383) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_311), .Y(n_305) );
AND2x2_ASAP7_75t_L g348 ( .A(n_306), .B(n_312), .Y(n_348) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g323 ( .A(n_307), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_307), .B(n_312), .Y(n_338) );
AND2x2_ASAP7_75t_L g371 ( .A(n_307), .B(n_316), .Y(n_371) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g313 ( .A(n_310), .Y(n_313) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g324 ( .A(n_312), .Y(n_324) );
INVx1_ASAP7_75t_L g388 ( .A(n_312), .Y(n_388) );
AND2x2_ASAP7_75t_L g322 ( .A(n_314), .B(n_323), .Y(n_322) );
AND2x4_ASAP7_75t_L g336 ( .A(n_314), .B(n_337), .Y(n_336) );
AND2x4_ASAP7_75t_L g347 ( .A(n_314), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_314), .B(n_323), .Y(n_814) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
OR2x2_ASAP7_75t_L g332 ( .A(n_315), .B(n_318), .Y(n_332) );
AND2x2_ASAP7_75t_L g343 ( .A(n_315), .B(n_318), .Y(n_343) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g377 ( .A(n_316), .B(n_318), .Y(n_377) );
INVx1_ASAP7_75t_L g372 ( .A(n_317), .Y(n_372) );
AND2x2_ASAP7_75t_L g387 ( .A(n_317), .B(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g358 ( .A(n_318), .Y(n_358) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx2_ASAP7_75t_L g600 ( .A(n_321), .Y(n_600) );
BUFx3_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx3_ASAP7_75t_L g407 ( .A(n_322), .Y(n_407) );
BUFx3_ASAP7_75t_L g457 ( .A(n_322), .Y(n_457) );
BUFx3_ASAP7_75t_L g524 ( .A(n_322), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g352 ( .A(n_323), .B(n_343), .Y(n_352) );
AND2x2_ASAP7_75t_L g416 ( .A(n_323), .B(n_343), .Y(n_416) );
INVx1_ASAP7_75t_L g379 ( .A(n_324), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_327), .B1(n_333), .B2(n_334), .Y(n_325) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVx4_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g452 ( .A(n_329), .Y(n_452) );
INVx5_ASAP7_75t_SL g519 ( .A(n_329), .Y(n_519) );
INVx2_ASAP7_75t_SL g630 ( .A(n_329), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g902 ( .A(n_329), .B(n_903), .Y(n_902) );
INVx11_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx11_ASAP7_75t_L g402 ( .A(n_330), .Y(n_402) );
AND2x4_ASAP7_75t_L g363 ( .A(n_331), .B(n_348), .Y(n_363) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g422 ( .A(n_332), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx3_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx3_ASAP7_75t_L g453 ( .A(n_336), .Y(n_453) );
BUFx2_ASAP7_75t_SL g520 ( .A(n_336), .Y(n_520) );
INVx1_ASAP7_75t_L g604 ( .A(n_336), .Y(n_604) );
BUFx3_ASAP7_75t_L g680 ( .A(n_336), .Y(n_680) );
BUFx2_ASAP7_75t_SL g863 ( .A(n_336), .Y(n_863) );
AND2x2_ASAP7_75t_L g617 ( .A(n_337), .B(n_372), .Y(n_617) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OR2x6_ASAP7_75t_L g357 ( .A(n_338), .B(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g810 ( .A(n_340), .Y(n_810) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx3_ASAP7_75t_L g403 ( .A(n_341), .Y(n_403) );
INVx2_ASAP7_75t_L g647 ( .A(n_341), .Y(n_647) );
OAI22xp5_ASAP7_75t_SL g893 ( .A1(n_341), .A2(n_456), .B1(n_894), .B2(n_895), .Y(n_893) );
INVx6_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx3_ASAP7_75t_L g511 ( .A(n_342), .Y(n_511) );
BUFx3_ASAP7_75t_L g599 ( .A(n_342), .Y(n_599) );
BUFx3_ASAP7_75t_L g631 ( .A(n_342), .Y(n_631) );
AND2x6_ASAP7_75t_L g365 ( .A(n_343), .B(n_348), .Y(n_365) );
NAND2x1p5_ASAP7_75t_L g427 ( .A(n_343), .B(n_348), .Y(n_427) );
INVx4_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx4_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g411 ( .A(n_347), .Y(n_411) );
BUFx3_ASAP7_75t_L g471 ( .A(n_347), .Y(n_471) );
BUFx3_ASAP7_75t_L g526 ( .A(n_347), .Y(n_526) );
BUFx3_ASAP7_75t_L g572 ( .A(n_347), .Y(n_572) );
INVx1_ASAP7_75t_L g423 ( .A(n_348), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_351), .B1(n_353), .B2(n_354), .Y(n_349) );
OAI21xp33_ASAP7_75t_L g607 ( .A1(n_351), .A2(n_608), .B(n_609), .Y(n_607) );
BUFx2_ASAP7_75t_R g351 ( .A(n_352), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g897 ( .A1(n_352), .A2(n_604), .B1(n_898), .B2(n_899), .Y(n_897) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx4f_ASAP7_75t_SL g417 ( .A(n_356), .Y(n_417) );
BUFx2_ASAP7_75t_L g474 ( .A(n_356), .Y(n_474) );
BUFx2_ASAP7_75t_L g567 ( .A(n_356), .Y(n_567) );
INVx6_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g516 ( .A(n_357), .Y(n_516) );
INVx1_ASAP7_75t_L g553 ( .A(n_357), .Y(n_553) );
INVx1_ASAP7_75t_SL g730 ( .A(n_357), .Y(n_730) );
INVx1_ASAP7_75t_L g466 ( .A(n_358), .Y(n_466) );
BUFx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx5_ASAP7_75t_L g463 ( .A(n_362), .Y(n_463) );
INVx2_ASAP7_75t_L g700 ( .A(n_362), .Y(n_700) );
INVx2_ASAP7_75t_L g742 ( .A(n_362), .Y(n_742) );
INVx4_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx4f_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx2_ASAP7_75t_L g596 ( .A(n_365), .Y(n_596) );
INVx1_ASAP7_75t_SL g651 ( .A(n_365), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B1(n_373), .B2(n_374), .Y(n_366) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx3_ASAP7_75t_SL g439 ( .A(n_369), .Y(n_439) );
INVx4_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx3_ASAP7_75t_L g504 ( .A(n_370), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_370), .A2(n_538), .B1(n_539), .B2(n_540), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_370), .A2(n_375), .B1(n_776), .B2(n_777), .Y(n_775) );
OAI22xp33_ASAP7_75t_SL g800 ( .A1(n_370), .A2(n_441), .B1(n_801), .B2(n_802), .Y(n_800) );
HB1xp67_ASAP7_75t_L g858 ( .A(n_370), .Y(n_858) );
OAI22xp5_ASAP7_75t_L g882 ( .A1(n_370), .A2(n_492), .B1(n_883), .B2(n_884), .Y(n_882) );
NAND2x1p5_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
AND2x4_ASAP7_75t_L g386 ( .A(n_371), .B(n_387), .Y(n_386) );
AND2x4_ASAP7_75t_L g391 ( .A(n_371), .B(n_392), .Y(n_391) );
AND2x4_ASAP7_75t_L g465 ( .A(n_371), .B(n_466), .Y(n_465) );
BUFx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
CKINVDCx16_ASAP7_75t_R g442 ( .A(n_375), .Y(n_442) );
OR2x6_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g468 ( .A(n_377), .B(n_379), .Y(n_468) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx4_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx2_ASAP7_75t_L g429 ( .A(n_382), .Y(n_429) );
OAI21xp5_ASAP7_75t_L g620 ( .A1(n_382), .A2(n_621), .B(n_622), .Y(n_620) );
OAI21xp5_ASAP7_75t_L g750 ( .A1(n_382), .A2(n_751), .B(n_752), .Y(n_750) );
INVx4_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_383), .Y(n_476) );
INVx2_ASAP7_75t_SL g497 ( .A(n_383), .Y(n_497) );
INVx2_ASAP7_75t_L g543 ( .A(n_383), .Y(n_543) );
BUFx3_ASAP7_75t_L g579 ( .A(n_383), .Y(n_579) );
INVx2_ASAP7_75t_SL g495 ( .A(n_384), .Y(n_495) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_386), .Y(n_432) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_386), .Y(n_478) );
BUFx4f_ASAP7_75t_SL g627 ( .A(n_386), .Y(n_627) );
BUFx2_ASAP7_75t_L g656 ( .A(n_386), .Y(n_656) );
INVx1_ASAP7_75t_L g392 ( .A(n_388), .Y(n_392) );
BUFx4f_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g480 ( .A(n_390), .Y(n_480) );
BUFx12f_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_391), .Y(n_436) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_391), .Y(n_501) );
INVx1_ASAP7_75t_L g737 ( .A(n_391), .Y(n_737) );
INVx1_ASAP7_75t_L g484 ( .A(n_395), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_445), .B1(n_446), .B2(n_482), .Y(n_395) );
INVx1_ASAP7_75t_L g482 ( .A(n_396), .Y(n_482) );
INVx1_ASAP7_75t_SL g444 ( .A(n_397), .Y(n_444) );
AND2x2_ASAP7_75t_SL g397 ( .A(n_398), .B(n_418), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_399), .B(n_408), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_404), .Y(n_399) );
INVx2_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVx4_ASAP7_75t_L g556 ( .A(n_402), .Y(n_556) );
INVx4_ASAP7_75t_L g570 ( .A(n_402), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_402), .B(n_611), .Y(n_610) );
BUFx3_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_412), .Y(n_408) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OAI21xp5_ASAP7_75t_SL g890 ( .A1(n_411), .A2(n_891), .B(n_892), .Y(n_890) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx2_ASAP7_75t_L g552 ( .A(n_414), .Y(n_552) );
INVx5_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx3_ASAP7_75t_L g473 ( .A(n_415), .Y(n_473) );
INVx4_ASAP7_75t_L g515 ( .A(n_415), .Y(n_515) );
INVx2_ASAP7_75t_L g566 ( .A(n_415), .Y(n_566) );
INVx8_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NOR3xp33_ASAP7_75t_L g418 ( .A(n_419), .B(n_428), .C(n_437), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B1(n_424), .B2(n_425), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_421), .A2(n_425), .B1(n_670), .B2(n_671), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_421), .A2(n_492), .B1(n_770), .B2(n_771), .Y(n_769) );
BUFx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_422), .Y(n_490) );
INVx2_ASAP7_75t_L g846 ( .A(n_422), .Y(n_846) );
OAI21xp5_ASAP7_75t_L g879 ( .A1(n_422), .A2(n_880), .B(n_881), .Y(n_879) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g460 ( .A(n_426), .Y(n_460) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx3_ASAP7_75t_L g492 ( .A(n_427), .Y(n_492) );
OAI221xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_430), .B1(n_431), .B2(n_433), .C(n_434), .Y(n_428) );
OAI221xp5_ASAP7_75t_L g665 ( .A1(n_431), .A2(n_543), .B1(n_666), .B2(n_667), .C(n_668), .Y(n_665) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_432), .Y(n_431) );
BUFx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g546 ( .A(n_436), .Y(n_546) );
BUFx3_ASAP7_75t_L g853 ( .A(n_436), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_439), .B1(n_440), .B2(n_441), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_439), .A2(n_540), .B1(n_673), .B2(n_674), .Y(n_672) );
OAI22xp5_ASAP7_75t_SL g503 ( .A1(n_441), .A2(n_504), .B1(n_505), .B2(n_506), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_441), .A2(n_857), .B1(n_858), .B2(n_859), .Y(n_856) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g540 ( .A(n_442), .Y(n_540) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
XOR2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_481), .Y(n_448) );
NAND4xp75_ASAP7_75t_L g449 ( .A(n_450), .B(n_458), .C(n_469), .D(n_475), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_454), .Y(n_450) );
INVx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx3_ASAP7_75t_L g780 ( .A(n_456), .Y(n_780) );
OA211x2_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_460), .B(n_461), .C(n_464), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_460), .A2(n_490), .B1(n_548), .B2(n_549), .Y(n_547) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx3_ASAP7_75t_L g576 ( .A(n_465), .Y(n_576) );
BUFx2_ASAP7_75t_L g593 ( .A(n_465), .Y(n_593) );
INVx1_ASAP7_75t_L g654 ( .A(n_465), .Y(n_654) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx3_ASAP7_75t_L g594 ( .A(n_468), .Y(n_594) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_472), .Y(n_469) );
INVx1_ASAP7_75t_L g817 ( .A(n_471), .Y(n_817) );
INVx2_ASAP7_75t_L g588 ( .A(n_476), .Y(n_588) );
INVx2_ASAP7_75t_SL g733 ( .A(n_476), .Y(n_733) );
BUFx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx4_ASAP7_75t_L g888 ( .A(n_478), .Y(n_888) );
INVx3_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g528 ( .A(n_485), .Y(n_528) );
XNOR2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_507), .Y(n_487) );
NOR3xp33_ASAP7_75t_L g488 ( .A(n_489), .B(n_494), .C(n_503), .Y(n_488) );
OAI22xp5_ASAP7_75t_SL g489 ( .A1(n_490), .A2(n_491), .B1(n_492), .B2(n_493), .Y(n_489) );
INVx1_ASAP7_75t_L g793 ( .A(n_490), .Y(n_793) );
BUFx3_ASAP7_75t_L g795 ( .A(n_492), .Y(n_795) );
INVx2_ASAP7_75t_L g849 ( .A(n_492), .Y(n_849) );
OAI222xp33_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B1(n_497), .B2(n_498), .C1(n_499), .C2(n_502), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g885 ( .A1(n_497), .A2(n_886), .B1(n_887), .B2(n_888), .Y(n_885) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx4f_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_508), .B(n_517), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_512), .Y(n_508) );
INVx1_ASAP7_75t_L g686 ( .A(n_511), .Y(n_686) );
INVx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx6f_ASAP7_75t_L g807 ( .A(n_515), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_521), .Y(n_517) );
INVx1_ASAP7_75t_L g726 ( .A(n_519), .Y(n_726) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx4f_ASAP7_75t_SL g723 ( .A(n_524), .Y(n_723) );
BUFx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g824 ( .A(n_529), .Y(n_824) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B1(n_638), .B2(n_822), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B1(n_560), .B2(n_637), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g559 ( .A(n_535), .Y(n_559) );
NAND2x1_ASAP7_75t_L g535 ( .A(n_536), .B(n_550), .Y(n_535) );
NOR3xp33_ASAP7_75t_SL g536 ( .A(n_537), .B(n_541), .C(n_547), .Y(n_536) );
OAI21xp33_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_543), .B(n_544), .Y(n_541) );
OAI21xp5_ASAP7_75t_L g695 ( .A1(n_543), .A2(n_696), .B(n_697), .Y(n_695) );
OAI221xp5_ASAP7_75t_L g850 ( .A1(n_543), .A2(n_851), .B1(n_852), .B2(n_854), .C(n_855), .Y(n_850) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND4x1_ASAP7_75t_L g550 ( .A(n_551), .B(n_554), .C(n_555), .D(n_557), .Y(n_550) );
INVx1_ASAP7_75t_L g637 ( .A(n_560), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_582), .B1(n_583), .B2(n_636), .Y(n_560) );
INVx1_ASAP7_75t_SL g636 ( .A(n_561), .Y(n_636) );
NOR4xp75_ASAP7_75t_L g562 ( .A(n_563), .B(n_568), .C(n_573), .D(n_577), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_569), .B(n_571), .Y(n_568) );
BUFx2_ASAP7_75t_L g602 ( .A(n_572), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_574), .B(n_575), .Y(n_573) );
OAI21xp5_ASAP7_75t_SL g577 ( .A1(n_578), .A2(n_580), .B(n_581), .Y(n_577) );
OAI21xp33_ASAP7_75t_SL g797 ( .A1(n_578), .A2(n_798), .B(n_799), .Y(n_797) );
INVx3_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
OAI22x1_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_612), .B1(n_634), .B2(n_635), .Y(n_583) );
INVx1_ASAP7_75t_L g634 ( .A(n_584), .Y(n_634) );
NAND3x1_ASAP7_75t_L g585 ( .A(n_586), .B(n_597), .C(n_605), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_591), .Y(n_586) );
OAI21xp5_ASAP7_75t_SL g587 ( .A1(n_588), .A2(n_589), .B(n_590), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_595), .Y(n_591) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_601), .Y(n_597) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_604), .A2(n_816), .B1(n_817), .B2(n_818), .Y(n_815) );
INVx1_ASAP7_75t_L g635 ( .A(n_612), .Y(n_635) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
XOR2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_633), .Y(n_613) );
NAND3x1_ASAP7_75t_L g614 ( .A(n_615), .B(n_619), .C(n_628), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
NOR2x1_ASAP7_75t_L g619 ( .A(n_620), .B(n_623), .Y(n_619) );
NAND3xp33_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .C(n_626), .Y(n_623) );
INVx1_ASAP7_75t_L g735 ( .A(n_627), .Y(n_735) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_632), .Y(n_628) );
INVx1_ASAP7_75t_L g822 ( .A(n_638), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_657), .B1(n_820), .B2(n_821), .Y(n_638) );
INVx2_ASAP7_75t_L g820 ( .A(n_639), .Y(n_820) );
NAND4xp75_ASAP7_75t_L g640 ( .A(n_641), .B(n_644), .C(n_648), .D(n_655), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
AND2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
AND2x2_ASAP7_75t_SL g648 ( .A(n_649), .B(n_652), .Y(n_648) );
INVx1_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g821 ( .A(n_657), .Y(n_821) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_659), .B1(n_712), .B2(n_713), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_689), .B1(n_690), .B2(n_711), .Y(n_661) );
INVx1_ASAP7_75t_L g711 ( .A(n_662), .Y(n_711) );
INVx2_ASAP7_75t_SL g688 ( .A(n_663), .Y(n_688) );
AND2x4_ASAP7_75t_L g663 ( .A(n_664), .B(n_675), .Y(n_663) );
NOR3xp33_ASAP7_75t_SL g664 ( .A(n_665), .B(n_669), .C(n_672), .Y(n_664) );
NOR2x1_ASAP7_75t_L g675 ( .A(n_676), .B(n_682), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_681), .Y(n_676) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx3_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
XOR2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_710), .Y(n_692) );
NAND2x1p5_ASAP7_75t_L g693 ( .A(n_694), .B(n_703), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_698), .Y(n_694) );
NAND3xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_701), .C(n_702), .Y(n_698) );
NOR2x1_ASAP7_75t_L g703 ( .A(n_704), .B(n_707), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
OAI22xp5_ASAP7_75t_SL g713 ( .A1(n_714), .A2(n_715), .B1(n_762), .B2(n_819), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_717), .B1(n_744), .B2(n_761), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g743 ( .A(n_719), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_731), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_727), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_724), .Y(n_721) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_732), .B(n_739), .Y(n_731) );
OAI222xp33_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_734), .B1(n_735), .B2(n_736), .C1(n_737), .C2(n_738), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
INVx3_ASAP7_75t_L g761 ( .A(n_744), .Y(n_761) );
XOR2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_760), .Y(n_744) );
NAND3x1_ASAP7_75t_SL g745 ( .A(n_746), .B(n_749), .C(n_757), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
NOR2x1_ASAP7_75t_L g749 ( .A(n_750), .B(n_753), .Y(n_749) );
NAND3xp33_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .C(n_756), .Y(n_753) );
AND2x2_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
INVx1_ASAP7_75t_L g819 ( .A(n_762), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_764), .B1(n_785), .B2(n_786), .Y(n_762) );
INVx2_ASAP7_75t_SL g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
AND3x1_ASAP7_75t_L g767 ( .A(n_768), .B(n_778), .C(n_782), .Y(n_767) );
NOR3xp33_ASAP7_75t_L g768 ( .A(n_769), .B(n_772), .C(n_775), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
AND2x2_ASAP7_75t_L g778 ( .A(n_779), .B(n_781), .Y(n_778) );
AND2x2_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
AND2x2_ASAP7_75t_L g789 ( .A(n_790), .B(n_803), .Y(n_789) );
NOR3xp33_ASAP7_75t_L g790 ( .A(n_791), .B(n_797), .C(n_800), .Y(n_790) );
OAI22xp5_ASAP7_75t_SL g791 ( .A1(n_792), .A2(n_794), .B1(n_795), .B2(n_796), .Y(n_791) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
NOR3xp33_ASAP7_75t_L g803 ( .A(n_804), .B(n_808), .C(n_815), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_805), .B(n_806), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_810), .B1(n_811), .B2(n_812), .Y(n_808) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
NOR2xp33_ASAP7_75t_L g900 ( .A(n_814), .B(n_901), .Y(n_900) );
INVx1_ASAP7_75t_SL g825 ( .A(n_826), .Y(n_825) );
NOR2x1_ASAP7_75t_L g826 ( .A(n_827), .B(n_831), .Y(n_826) );
OR2x2_ASAP7_75t_SL g906 ( .A(n_827), .B(n_832), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_828), .B(n_830), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
OAI322xp33_ASAP7_75t_L g838 ( .A1(n_829), .A2(n_839), .A3(n_869), .B1(n_871), .B2(n_874), .C1(n_875), .C2(n_904), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_829), .B(n_870), .Y(n_873) );
CKINVDCx16_ASAP7_75t_R g870 ( .A(n_830), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_832), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_833), .B(n_834), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_836), .B(n_837), .Y(n_835) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_842), .B(n_860), .Y(n_841) );
NOR3xp33_ASAP7_75t_L g842 ( .A(n_843), .B(n_850), .C(n_856), .Y(n_842) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_845), .B1(n_847), .B2(n_848), .Y(n_843) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx2_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx2_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
NOR2xp33_ASAP7_75t_L g860 ( .A(n_861), .B(n_865), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_862), .B(n_864), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
CKINVDCx16_ASAP7_75t_R g871 ( .A(n_872), .Y(n_871) );
XNOR2x1_ASAP7_75t_L g876 ( .A(n_874), .B(n_877), .Y(n_876) );
BUFx2_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
AND3x2_ASAP7_75t_L g877 ( .A(n_878), .B(n_889), .C(n_896), .Y(n_877) );
NOR3xp33_ASAP7_75t_L g878 ( .A(n_879), .B(n_882), .C(n_885), .Y(n_878) );
NOR2xp33_ASAP7_75t_L g889 ( .A(n_890), .B(n_893), .Y(n_889) );
NOR3xp33_ASAP7_75t_L g896 ( .A(n_897), .B(n_900), .C(n_902), .Y(n_896) );
CKINVDCx20_ASAP7_75t_R g904 ( .A(n_905), .Y(n_904) );
CKINVDCx20_ASAP7_75t_R g905 ( .A(n_906), .Y(n_905) );
endmodule