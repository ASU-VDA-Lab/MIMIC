module fake_jpeg_17184_n_378 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_378);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_378;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx8_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx2_ASAP7_75t_SL g16 ( 
.A(n_8),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_5),
.B(n_2),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_39),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_13),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_40),
.B(n_46),
.Y(n_84)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx2_ASAP7_75t_SL g90 ( 
.A(n_42),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_49),
.Y(n_74)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_56),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_35),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_19),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_58),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx5_ASAP7_75t_SL g81 ( 
.A(n_59),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_18),
.B(n_12),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_64),
.Y(n_120)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_25),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_68),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_26),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_25),
.B(n_0),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_73),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_26),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_46),
.B(n_20),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_75),
.B(n_114),
.Y(n_140)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_23),
.B1(n_16),
.B2(n_29),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_77),
.A2(n_116),
.B1(n_70),
.B2(n_72),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_41),
.A2(n_16),
.B1(n_27),
.B2(n_37),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_80),
.A2(n_97),
.B1(n_101),
.B2(n_122),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_52),
.A2(n_33),
.B1(n_28),
.B2(n_29),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_82),
.A2(n_85),
.B1(n_86),
.B2(n_105),
.Y(n_158)
);

AO22x1_ASAP7_75t_SL g85 ( 
.A1(n_59),
.A2(n_37),
.B1(n_27),
.B2(n_15),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_44),
.A2(n_20),
.B1(n_27),
.B2(n_37),
.Y(n_86)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_47),
.A2(n_37),
.B1(n_27),
.B2(n_28),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_99),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_42),
.A2(n_33),
.B1(n_15),
.B2(n_14),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_39),
.A2(n_14),
.B1(n_30),
.B2(n_21),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_65),
.A2(n_14),
.B1(n_15),
.B2(n_31),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_106),
.A2(n_59),
.B1(n_53),
.B2(n_50),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_56),
.B(n_32),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_119),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_66),
.B(n_30),
.C(n_21),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_108),
.B(n_4),
.C(n_5),
.Y(n_160)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_57),
.B(n_30),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_62),
.A2(n_15),
.B1(n_32),
.B2(n_21),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_30),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_118),
.B(n_4),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_32),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_49),
.A2(n_15),
.B1(n_1),
.B2(n_2),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_51),
.A2(n_30),
.B1(n_21),
.B2(n_3),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_123),
.A2(n_53),
.B1(n_61),
.B2(n_60),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_SL g187 ( 
.A1(n_124),
.A2(n_85),
.B(n_81),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_127),
.A2(n_144),
.B1(n_172),
.B2(n_78),
.Y(n_176)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_129),
.A2(n_143),
.B1(n_154),
.B2(n_166),
.Y(n_198)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_130),
.Y(n_188)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_132),
.Y(n_196)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_136),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_58),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_134),
.B(n_141),
.Y(n_180)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_135),
.Y(n_197)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_137),
.Y(n_202)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_148),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_54),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_76),
.A2(n_55),
.B1(n_64),
.B2(n_70),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_74),
.A2(n_43),
.B1(n_66),
.B2(n_3),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g145 ( 
.A(n_92),
.B(n_66),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_145),
.B(n_160),
.C(n_144),
.Y(n_211)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_146),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_82),
.B(n_0),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_165),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_80),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_95),
.B(n_0),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_149),
.B(n_150),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_96),
.B(n_1),
.Y(n_150)
);

NAND2x1_ASAP7_75t_SL g151 ( 
.A(n_85),
.B(n_3),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_151),
.A2(n_109),
.B(n_117),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_102),
.Y(n_152)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

INVxp33_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_155),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_L g154 ( 
.A1(n_88),
.A2(n_111),
.B1(n_94),
.B2(n_104),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_99),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_97),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_162),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g157 ( 
.A(n_79),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_159),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_163),
.Y(n_208)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_89),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_113),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_169),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_84),
.B(n_4),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_122),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_108),
.B(n_6),
.Y(n_168)
);

AOI21xp33_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_9),
.B(n_101),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_121),
.B(n_10),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_113),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_170),
.B(n_152),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_79),
.Y(n_171)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_171),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_98),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_78),
.A2(n_10),
.B1(n_7),
.B2(n_9),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_173),
.A2(n_98),
.B1(n_81),
.B2(n_88),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_176),
.A2(n_189),
.B1(n_200),
.B2(n_214),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_181),
.A2(n_125),
.B1(n_142),
.B2(n_138),
.Y(n_229)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_183),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_187),
.A2(n_164),
.B1(n_130),
.B2(n_157),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_156),
.A2(n_104),
.B1(n_115),
.B2(n_120),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_191),
.Y(n_232)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_136),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_203),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_128),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_206),
.Y(n_222)
);

OAI21xp33_ASAP7_75t_L g242 ( 
.A1(n_195),
.A2(n_161),
.B(n_152),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_L g200 ( 
.A1(n_167),
.A2(n_115),
.B1(n_100),
.B2(n_110),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_123),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_211),
.Y(n_225)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_139),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_137),
.Y(n_204)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_204),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_132),
.Y(n_206)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_133),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_190),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_208),
.B(n_194),
.Y(n_235)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_212),
.Y(n_245)
);

NOR2x1_ASAP7_75t_L g213 ( 
.A(n_151),
.B(n_147),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_213),
.B(n_126),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_148),
.A2(n_127),
.B1(n_168),
.B2(n_158),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_131),
.B(n_140),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_157),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_145),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_218),
.B(n_230),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_213),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_220),
.A2(n_179),
.B1(n_174),
.B2(n_183),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_214),
.A2(n_158),
.B1(n_125),
.B2(n_142),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_221),
.A2(n_251),
.B1(n_252),
.B2(n_205),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_176),
.A2(n_211),
.B1(n_185),
.B2(n_210),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_223),
.A2(n_234),
.B1(n_188),
.B2(n_175),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_182),
.B(n_151),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_227),
.A2(n_231),
.B(n_235),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_177),
.A2(n_145),
.B(n_155),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_228),
.A2(n_236),
.B(n_243),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_182),
.B(n_140),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_166),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_208),
.B(n_165),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_239),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_198),
.A2(n_138),
.B1(n_159),
.B2(n_135),
.Y(n_234)
);

AO22x1_ASAP7_75t_SL g237 ( 
.A1(n_198),
.A2(n_154),
.B1(n_126),
.B2(n_170),
.Y(n_237)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_238),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_199),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_240),
.B(n_248),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_242),
.A2(n_247),
.B(n_228),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_180),
.B(n_157),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_253),
.Y(n_276)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_193),
.A2(n_206),
.B(n_184),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_197),
.B(n_171),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_186),
.Y(n_249)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_249),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_178),
.B(n_204),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_250),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_200),
.A2(n_196),
.B1(n_216),
.B2(n_197),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_196),
.A2(n_216),
.B1(n_188),
.B2(n_202),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_205),
.B(n_202),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_254),
.B(n_265),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_191),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_257),
.B(n_266),
.C(n_269),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_258),
.A2(n_263),
.B1(n_270),
.B2(n_256),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_237),
.A2(n_179),
.B1(n_209),
.B2(n_174),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_264),
.A2(n_277),
.B1(n_237),
.B2(n_251),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_222),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_225),
.B(n_178),
.C(n_207),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_218),
.B(n_239),
.C(n_235),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_221),
.A2(n_192),
.B1(n_203),
.B2(n_207),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_223),
.B(n_233),
.C(n_220),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_273),
.C(n_248),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_230),
.B(n_247),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_274),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_236),
.B(n_244),
.C(n_217),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_222),
.B(n_227),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_227),
.B(n_240),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_282),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_237),
.A2(n_217),
.B1(n_243),
.B2(n_234),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_279),
.B(n_278),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_246),
.Y(n_280)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_280),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_231),
.B(n_245),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_249),
.Y(n_284)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_263),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_285),
.B(n_290),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_287),
.A2(n_300),
.B1(n_307),
.B2(n_264),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_268),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_283),
.A2(n_245),
.B(n_231),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_291),
.A2(n_274),
.B1(n_283),
.B2(n_265),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_267),
.A2(n_241),
.B1(n_219),
.B2(n_232),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_292),
.A2(n_296),
.B1(n_258),
.B2(n_270),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_260),
.B(n_241),
.Y(n_293)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_293),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_254),
.Y(n_294)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_294),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_256),
.A2(n_219),
.B1(n_232),
.B2(n_252),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_306),
.C(n_308),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_262),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_268),
.Y(n_301)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_301),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_281),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_302),
.Y(n_311)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_280),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_303),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_260),
.B(n_224),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_304),
.B(n_286),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_271),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_257),
.B(n_226),
.C(n_266),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_257),
.B(n_226),
.C(n_269),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_281),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_309),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_313),
.C(n_315),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_273),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_278),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_316),
.A2(n_285),
.B1(n_292),
.B2(n_287),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_319),
.B(n_255),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_320),
.A2(n_282),
.B1(n_289),
.B2(n_275),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_295),
.B(n_259),
.C(n_261),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_323),
.C(n_324),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_259),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_261),
.C(n_276),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_298),
.B(n_279),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_326),
.B(n_329),
.C(n_272),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_328),
.B(n_300),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_291),
.B(n_276),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_327),
.A2(n_294),
.B(n_297),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_330),
.A2(n_341),
.B(n_322),
.Y(n_349)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_331),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_318),
.A2(n_288),
.B1(n_303),
.B2(n_289),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_336),
.Y(n_354)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_333),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_320),
.A2(n_288),
.B1(n_277),
.B2(n_309),
.Y(n_334)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_334),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_338),
.B(n_342),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_328),
.A2(n_296),
.B1(n_299),
.B2(n_301),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_339),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_314),
.B(n_255),
.C(n_299),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_340),
.B(n_343),
.C(n_344),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_310),
.A2(n_262),
.B1(n_284),
.B2(n_329),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_314),
.B(n_313),
.C(n_315),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_324),
.Y(n_344)
);

AOI21x1_ASAP7_75t_L g345 ( 
.A1(n_321),
.A2(n_317),
.B(n_326),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_345),
.A2(n_325),
.B(n_332),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_349),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_330),
.A2(n_312),
.B(n_323),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_351),
.A2(n_337),
.B(n_349),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_335),
.B(n_311),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_355),
.B(n_357),
.C(n_343),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_356),
.B(n_342),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_335),
.B(n_338),
.Y(n_357)
);

NOR2xp67_ASAP7_75t_SL g359 ( 
.A(n_356),
.B(n_340),
.Y(n_359)
);

AOI31xp67_ASAP7_75t_SL g369 ( 
.A1(n_359),
.A2(n_350),
.A3(n_351),
.B(n_346),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_362),
.Y(n_368)
);

BUFx24_ASAP7_75t_SL g361 ( 
.A(n_352),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_361),
.B(n_363),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_348),
.A2(n_331),
.B1(n_339),
.B2(n_334),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_364),
.B(n_355),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_366),
.B(n_367),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_358),
.Y(n_367)
);

AOI221xp5_ASAP7_75t_L g370 ( 
.A1(n_369),
.A2(n_354),
.B1(n_350),
.B2(n_362),
.C(n_353),
.Y(n_370)
);

NAND3xp33_ASAP7_75t_L g374 ( 
.A(n_370),
.B(n_371),
.C(n_368),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_367),
.A2(n_346),
.B(n_357),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_372),
.B(n_365),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_373),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_375),
.B(n_374),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_376),
.B(n_337),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_377),
.B(n_347),
.Y(n_378)
);


endmodule