module real_aes_6677_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_746;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_733;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g112 ( .A(n_0), .Y(n_112) );
INVx1_ASAP7_75t_L g510 ( .A(n_1), .Y(n_510) );
INVx1_ASAP7_75t_L g267 ( .A(n_2), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_3), .A2(n_38), .B1(n_186), .B2(n_538), .Y(n_537) );
AOI21xp33_ASAP7_75t_L g174 ( .A1(n_4), .A2(n_175), .B(n_176), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_5), .B(n_173), .Y(n_487) );
AND2x6_ASAP7_75t_L g148 ( .A(n_6), .B(n_149), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_7), .A2(n_243), .B(n_244), .Y(n_242) );
INVx1_ASAP7_75t_L g110 ( .A(n_8), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_8), .B(n_39), .Y(n_451) );
INVx1_ASAP7_75t_L g183 ( .A(n_9), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_10), .B(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g145 ( .A(n_11), .Y(n_145) );
INVx1_ASAP7_75t_L g506 ( .A(n_12), .Y(n_506) );
INVx1_ASAP7_75t_L g249 ( .A(n_13), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_14), .B(n_151), .Y(n_544) );
AOI222xp33_ASAP7_75t_SL g455 ( .A1(n_15), .A2(n_456), .B1(n_457), .B2(n_466), .C1(n_754), .C2(n_755), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_16), .B(n_141), .Y(n_515) );
XNOR2xp5_ASAP7_75t_L g123 ( .A(n_17), .B(n_124), .Y(n_123) );
AO32x2_ASAP7_75t_L g535 ( .A1(n_17), .A2(n_140), .A3(n_173), .B1(n_498), .B2(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_18), .B(n_186), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_19), .B(n_194), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_20), .B(n_141), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_21), .A2(n_51), .B1(n_186), .B2(n_538), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_22), .B(n_175), .Y(n_203) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_23), .A2(n_78), .B1(n_151), .B2(n_186), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_24), .B(n_186), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_25), .B(n_171), .Y(n_197) );
OAI22xp5_ASAP7_75t_SL g457 ( .A1(n_26), .A2(n_458), .B1(n_459), .B2(n_465), .Y(n_457) );
INVx1_ASAP7_75t_L g465 ( .A(n_26), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_27), .A2(n_247), .B(n_248), .C(n_250), .Y(n_246) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_28), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_29), .B(n_188), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_30), .B(n_181), .Y(n_268) );
INVx1_ASAP7_75t_L g159 ( .A(n_31), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_32), .B(n_188), .Y(n_532) );
INVx2_ASAP7_75t_L g153 ( .A(n_33), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_34), .B(n_186), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_35), .B(n_188), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g128 ( .A1(n_36), .A2(n_42), .B1(n_129), .B2(n_130), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_36), .Y(n_130) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_37), .A2(n_148), .B(n_160), .C(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_39), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g157 ( .A(n_40), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_41), .B(n_181), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_42), .Y(n_129) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_43), .A2(n_105), .B1(n_116), .B2(n_759), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_44), .B(n_186), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_45), .A2(n_88), .B1(n_211), .B2(n_538), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_46), .B(n_186), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_47), .B(n_186), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g163 ( .A(n_48), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_49), .B(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_50), .B(n_175), .Y(n_237) );
AOI22xp33_ASAP7_75t_SL g519 ( .A1(n_52), .A2(n_61), .B1(n_151), .B2(n_186), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g150 ( .A1(n_53), .A2(n_151), .B1(n_154), .B2(n_160), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g214 ( .A(n_54), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_55), .B(n_186), .Y(n_497) );
CKINVDCx16_ASAP7_75t_R g264 ( .A(n_56), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_57), .B(n_186), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_58), .A2(n_180), .B(n_182), .C(n_185), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_59), .Y(n_224) );
INVx1_ASAP7_75t_L g177 ( .A(n_60), .Y(n_177) );
INVx1_ASAP7_75t_L g149 ( .A(n_62), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_63), .B(n_186), .Y(n_511) );
INVx1_ASAP7_75t_L g144 ( .A(n_64), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_65), .Y(n_121) );
AO32x2_ASAP7_75t_L g555 ( .A1(n_66), .A2(n_173), .A3(n_229), .B1(n_498), .B2(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g495 ( .A(n_67), .Y(n_495) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_68), .A2(n_127), .B1(n_128), .B2(n_131), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_68), .Y(n_131) );
INVx1_ASAP7_75t_L g527 ( .A(n_69), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_SL g193 ( .A1(n_70), .A2(n_185), .B(n_194), .C(n_195), .Y(n_193) );
INVxp67_ASAP7_75t_L g196 ( .A(n_71), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_72), .B(n_151), .Y(n_528) );
INVx1_ASAP7_75t_L g115 ( .A(n_73), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_74), .Y(n_168) );
INVx1_ASAP7_75t_L g217 ( .A(n_75), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_76), .A2(n_102), .B1(n_463), .B2(n_464), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_76), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_77), .B(n_453), .Y(n_452) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_79), .A2(n_148), .B(n_160), .C(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_80), .B(n_538), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_81), .B(n_151), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_82), .B(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g142 ( .A(n_83), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_84), .B(n_194), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_85), .B(n_151), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_86), .A2(n_148), .B(n_160), .C(n_266), .Y(n_265) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_87), .B(n_112), .C(n_113), .Y(n_111) );
OR2x2_ASAP7_75t_L g448 ( .A(n_87), .B(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g469 ( .A(n_87), .B(n_450), .Y(n_469) );
INVx2_ASAP7_75t_L g753 ( .A(n_87), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_89), .A2(n_103), .B1(n_151), .B2(n_152), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_90), .B(n_188), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g271 ( .A(n_91), .Y(n_271) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_92), .A2(n_148), .B(n_160), .C(n_232), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_93), .Y(n_239) );
INVx1_ASAP7_75t_L g192 ( .A(n_94), .Y(n_192) );
CKINVDCx16_ASAP7_75t_R g245 ( .A(n_95), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_96), .B(n_207), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_97), .A2(n_460), .B1(n_461), .B2(n_462), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_97), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_98), .B(n_151), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_99), .B(n_173), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_100), .B(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_101), .A2(n_175), .B(n_191), .Y(n_190) );
CKINVDCx16_ASAP7_75t_R g464 ( .A(n_102), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx5_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
CKINVDCx9p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_108), .Y(n_760) );
OR2x4_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
AND2x2_ASAP7_75t_L g450 ( .A(n_112), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
OA21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_122), .B(n_454), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g758 ( .A(n_121), .Y(n_758) );
OAI21x1_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_445), .B(n_452), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_126), .B1(n_132), .B2(n_133), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_126), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_128), .Y(n_127) );
OAI22xp5_ASAP7_75t_SL g466 ( .A1(n_132), .A2(n_467), .B1(n_470), .B2(n_750), .Y(n_466) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OAI22xp5_ASAP7_75t_SL g755 ( .A1(n_133), .A2(n_467), .B1(n_756), .B2(n_757), .Y(n_755) );
AND3x1_ASAP7_75t_L g133 ( .A(n_134), .B(n_370), .C(n_419), .Y(n_133) );
NOR3xp33_ASAP7_75t_SL g134 ( .A(n_135), .B(n_277), .C(n_315), .Y(n_134) );
OAI222xp33_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_198), .B1(n_252), .B2(n_258), .C1(n_272), .C2(n_275), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_169), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_137), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_137), .B(n_320), .Y(n_411) );
BUFx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OR2x2_ASAP7_75t_L g288 ( .A(n_138), .B(n_189), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_138), .B(n_170), .Y(n_296) );
AND2x2_ASAP7_75t_L g331 ( .A(n_138), .B(n_308), .Y(n_331) );
OR2x2_ASAP7_75t_L g355 ( .A(n_138), .B(n_170), .Y(n_355) );
OR2x2_ASAP7_75t_L g363 ( .A(n_138), .B(n_262), .Y(n_363) );
AND2x2_ASAP7_75t_L g366 ( .A(n_138), .B(n_189), .Y(n_366) );
INVx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OR2x2_ASAP7_75t_L g260 ( .A(n_139), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g274 ( .A(n_139), .B(n_189), .Y(n_274) );
AND2x2_ASAP7_75t_L g324 ( .A(n_139), .B(n_262), .Y(n_324) );
AND2x2_ASAP7_75t_L g337 ( .A(n_139), .B(n_170), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_139), .B(n_423), .Y(n_444) );
AO21x2_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_146), .B(n_167), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_140), .B(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g212 ( .A(n_140), .Y(n_212) );
AO21x2_ASAP7_75t_L g262 ( .A1(n_140), .A2(n_263), .B(n_270), .Y(n_262) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_141), .Y(n_173) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AND2x2_ASAP7_75t_SL g188 ( .A(n_142), .B(n_143), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
OAI22xp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_150), .B1(n_163), .B2(n_164), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_L g176 ( .A1(n_147), .A2(n_177), .B(n_178), .C(n_179), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_L g191 ( .A1(n_147), .A2(n_178), .B(n_192), .C(n_193), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_147), .A2(n_178), .B(n_245), .C(n_246), .Y(n_244) );
INVx4_ASAP7_75t_SL g147 ( .A(n_148), .Y(n_147) );
NAND2x1p5_ASAP7_75t_L g164 ( .A(n_148), .B(n_165), .Y(n_164) );
AND2x4_ASAP7_75t_L g175 ( .A(n_148), .B(n_165), .Y(n_175) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_148), .A2(n_479), .B(n_482), .Y(n_478) );
BUFx3_ASAP7_75t_L g498 ( .A(n_148), .Y(n_498) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_148), .A2(n_505), .B(n_509), .Y(n_504) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_148), .A2(n_526), .B(n_529), .Y(n_525) );
OAI21xp5_ASAP7_75t_L g541 ( .A1(n_148), .A2(n_542), .B(n_546), .Y(n_541) );
INVx2_ASAP7_75t_L g269 ( .A(n_151), .Y(n_269) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g161 ( .A(n_153), .Y(n_161) );
INVx1_ASAP7_75t_L g166 ( .A(n_153), .Y(n_166) );
OAI22xp5_ASAP7_75t_SL g154 ( .A1(n_155), .A2(n_157), .B1(n_158), .B2(n_159), .Y(n_154) );
INVx2_ASAP7_75t_L g158 ( .A(n_155), .Y(n_158) );
INVx4_ASAP7_75t_L g247 ( .A(n_155), .Y(n_247) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g162 ( .A(n_156), .Y(n_162) );
AND2x2_ASAP7_75t_L g165 ( .A(n_156), .B(n_166), .Y(n_165) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_156), .Y(n_181) );
INVx3_ASAP7_75t_L g184 ( .A(n_156), .Y(n_184) );
INVx1_ASAP7_75t_L g194 ( .A(n_156), .Y(n_194) );
INVx5_ASAP7_75t_L g178 ( .A(n_160), .Y(n_178) );
AND2x6_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_161), .Y(n_186) );
BUFx3_ASAP7_75t_L g211 ( .A(n_161), .Y(n_211) );
INVx1_ASAP7_75t_L g538 ( .A(n_161), .Y(n_538) );
OAI21xp5_ASAP7_75t_L g216 ( .A1(n_164), .A2(n_217), .B(n_218), .Y(n_216) );
OAI21xp5_ASAP7_75t_L g263 ( .A1(n_164), .A2(n_264), .B(n_265), .Y(n_263) );
INVx1_ASAP7_75t_L g485 ( .A(n_166), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_L g362 ( .A1(n_169), .A2(n_363), .B(n_364), .C(n_367), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_169), .B(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_169), .B(n_307), .Y(n_429) );
AND2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_189), .Y(n_169) );
AND2x2_ASAP7_75t_SL g273 ( .A(n_170), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g287 ( .A(n_170), .Y(n_287) );
AND2x2_ASAP7_75t_L g314 ( .A(n_170), .B(n_308), .Y(n_314) );
INVx1_ASAP7_75t_SL g322 ( .A(n_170), .Y(n_322) );
AND2x2_ASAP7_75t_L g345 ( .A(n_170), .B(n_346), .Y(n_345) );
BUFx2_ASAP7_75t_L g423 ( .A(n_170), .Y(n_423) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_174), .B(n_187), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_SL g213 ( .A(n_172), .B(n_214), .Y(n_213) );
NAND3xp33_ASAP7_75t_L g516 ( .A(n_172), .B(n_498), .C(n_517), .Y(n_516) );
AO21x1_ASAP7_75t_L g561 ( .A1(n_172), .A2(n_517), .B(n_562), .Y(n_561) );
INVx4_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
OA21x2_ASAP7_75t_L g189 ( .A1(n_173), .A2(n_190), .B(n_197), .Y(n_189) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_173), .A2(n_478), .B(n_487), .Y(n_477) );
BUFx2_ASAP7_75t_L g243 ( .A(n_175), .Y(n_243) );
O2A1O1Ixp5_ASAP7_75t_L g494 ( .A1(n_180), .A2(n_495), .B(n_496), .C(n_497), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_180), .A2(n_547), .B(n_548), .Y(n_546) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx4_ASAP7_75t_L g235 ( .A(n_181), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_181), .A2(n_486), .B1(n_518), .B2(n_519), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_181), .A2(n_486), .B1(n_537), .B2(n_539), .Y(n_536) );
OAI22xp5_ASAP7_75t_SL g556 ( .A1(n_181), .A2(n_184), .B1(n_557), .B2(n_558), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_183), .B(n_184), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_184), .B(n_196), .Y(n_195) );
INVx5_ASAP7_75t_L g207 ( .A(n_184), .Y(n_207) );
O2A1O1Ixp5_ASAP7_75t_SL g526 ( .A1(n_185), .A2(n_207), .B(n_527), .C(n_528), .Y(n_526) );
INVx3_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_186), .Y(n_236) );
INVx1_ASAP7_75t_L g225 ( .A(n_188), .Y(n_225) );
INVx2_ASAP7_75t_L g229 ( .A(n_188), .Y(n_229) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_188), .A2(n_242), .B(n_251), .Y(n_241) );
OA21x2_ASAP7_75t_L g524 ( .A1(n_188), .A2(n_525), .B(n_532), .Y(n_524) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_188), .A2(n_541), .B(n_549), .Y(n_540) );
BUFx2_ASAP7_75t_L g259 ( .A(n_189), .Y(n_259) );
INVx1_ASAP7_75t_L g321 ( .A(n_189), .Y(n_321) );
INVx3_ASAP7_75t_L g346 ( .A(n_189), .Y(n_346) );
INVx1_ASAP7_75t_L g545 ( .A(n_194), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_198), .B(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_226), .Y(n_198) );
INVx1_ASAP7_75t_L g342 ( .A(n_199), .Y(n_342) );
OAI32xp33_ASAP7_75t_L g348 ( .A1(n_199), .A2(n_287), .A3(n_349), .B1(n_350), .B2(n_351), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_199), .A2(n_353), .B1(n_356), .B2(n_361), .Y(n_352) );
INVx4_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g290 ( .A(n_200), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g368 ( .A(n_200), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g438 ( .A(n_200), .B(n_384), .Y(n_438) );
AND2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_215), .Y(n_200) );
AND2x2_ASAP7_75t_L g253 ( .A(n_201), .B(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g283 ( .A(n_201), .Y(n_283) );
INVx1_ASAP7_75t_L g302 ( .A(n_201), .Y(n_302) );
OR2x2_ASAP7_75t_L g310 ( .A(n_201), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g317 ( .A(n_201), .B(n_291), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_201), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g338 ( .A(n_201), .B(n_256), .Y(n_338) );
INVx3_ASAP7_75t_L g360 ( .A(n_201), .Y(n_360) );
AND2x2_ASAP7_75t_L g385 ( .A(n_201), .B(n_257), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_201), .B(n_350), .Y(n_433) );
OR2x6_ASAP7_75t_L g201 ( .A(n_202), .B(n_213), .Y(n_201) );
AOI21xp5_ASAP7_75t_SL g202 ( .A1(n_203), .A2(n_204), .B(n_212), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_208), .B(n_209), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g266 ( .A1(n_207), .A2(n_267), .B(n_268), .C(n_269), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_207), .A2(n_480), .B(n_481), .Y(n_479) );
INVx2_ASAP7_75t_L g486 ( .A(n_207), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_207), .A2(n_492), .B(n_493), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_209), .A2(n_220), .B(n_221), .Y(n_219) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g250 ( .A(n_211), .Y(n_250) );
INVx1_ASAP7_75t_L g222 ( .A(n_212), .Y(n_222) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_212), .A2(n_490), .B(n_499), .Y(n_489) );
OA21x2_ASAP7_75t_L g503 ( .A1(n_212), .A2(n_504), .B(n_512), .Y(n_503) );
INVx2_ASAP7_75t_L g257 ( .A(n_215), .Y(n_257) );
AND2x2_ASAP7_75t_L g389 ( .A(n_215), .B(n_227), .Y(n_389) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_222), .B(n_223), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_225), .B(n_239), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_225), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g431 ( .A(n_226), .Y(n_431) );
OR2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_240), .Y(n_226) );
INVx1_ASAP7_75t_L g276 ( .A(n_227), .Y(n_276) );
AND2x2_ASAP7_75t_L g303 ( .A(n_227), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_227), .B(n_257), .Y(n_311) );
AND2x2_ASAP7_75t_L g369 ( .A(n_227), .B(n_292), .Y(n_369) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g255 ( .A(n_228), .Y(n_255) );
AND2x2_ASAP7_75t_L g282 ( .A(n_228), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g291 ( .A(n_228), .B(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_228), .B(n_257), .Y(n_357) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_238), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_237), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_236), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_240), .B(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g304 ( .A(n_240), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_240), .B(n_257), .Y(n_350) );
AND2x2_ASAP7_75t_L g359 ( .A(n_240), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g384 ( .A(n_240), .Y(n_384) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g256 ( .A(n_241), .B(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g292 ( .A(n_241), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_247), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g508 ( .A(n_247), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_247), .A2(n_530), .B(n_531), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_252), .A2(n_262), .B1(n_421), .B2(n_424), .Y(n_420) );
INVx1_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
OAI21xp5_ASAP7_75t_SL g443 ( .A1(n_254), .A2(n_365), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_255), .B(n_360), .Y(n_377) );
INVx1_ASAP7_75t_L g402 ( .A(n_255), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_256), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g329 ( .A(n_256), .B(n_282), .Y(n_329) );
INVx2_ASAP7_75t_L g285 ( .A(n_257), .Y(n_285) );
INVx1_ASAP7_75t_L g335 ( .A(n_257), .Y(n_335) );
OAI221xp5_ASAP7_75t_L g426 ( .A1(n_258), .A2(n_410), .B1(n_427), .B2(n_430), .C(n_432), .Y(n_426) );
OR2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
INVx1_ASAP7_75t_L g297 ( .A(n_259), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_259), .B(n_308), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_260), .B(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g351 ( .A(n_260), .B(n_297), .Y(n_351) );
INVx3_ASAP7_75t_SL g392 ( .A(n_260), .Y(n_392) );
AND2x2_ASAP7_75t_L g336 ( .A(n_261), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g365 ( .A(n_261), .B(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_261), .B(n_274), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_261), .B(n_320), .Y(n_406) );
INVx3_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx3_ASAP7_75t_L g308 ( .A(n_262), .Y(n_308) );
OAI322xp33_ASAP7_75t_L g403 ( .A1(n_262), .A2(n_334), .A3(n_356), .B1(n_404), .B2(n_406), .C1(n_407), .C2(n_408), .Y(n_403) );
O2A1O1Ixp33_ASAP7_75t_L g505 ( .A1(n_269), .A2(n_506), .B(n_507), .C(n_508), .Y(n_505) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AOI21xp33_ASAP7_75t_L g427 ( .A1(n_273), .A2(n_276), .B(n_428), .Y(n_427) );
NOR2xp33_ASAP7_75t_SL g353 ( .A(n_274), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g375 ( .A(n_274), .B(n_287), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_274), .B(n_314), .Y(n_390) );
INVxp67_ASAP7_75t_L g341 ( .A(n_276), .Y(n_341) );
AOI211xp5_ASAP7_75t_L g347 ( .A1(n_276), .A2(n_348), .B(n_352), .C(n_362), .Y(n_347) );
OAI221xp5_ASAP7_75t_SL g277 ( .A1(n_278), .A2(n_286), .B1(n_289), .B2(n_293), .C(n_298), .Y(n_277) );
INVxp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_284), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g301 ( .A(n_285), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g418 ( .A(n_285), .Y(n_418) );
OAI221xp5_ASAP7_75t_L g434 ( .A1(n_286), .A2(n_435), .B1(n_440), .B2(n_441), .C(n_443), .Y(n_434) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_287), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_SL g334 ( .A(n_287), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_287), .B(n_365), .Y(n_372) );
AND2x2_ASAP7_75t_L g414 ( .A(n_287), .B(n_392), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_288), .B(n_313), .Y(n_312) );
OAI22xp33_ASAP7_75t_L g409 ( .A1(n_288), .A2(n_300), .B1(n_410), .B2(n_411), .Y(n_409) );
OR2x2_ASAP7_75t_L g440 ( .A(n_288), .B(n_308), .Y(n_440) );
CKINVDCx16_ASAP7_75t_R g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g417 ( .A(n_291), .Y(n_417) );
AND2x2_ASAP7_75t_L g442 ( .A(n_291), .B(n_385), .Y(n_442) );
INVxp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NOR2xp33_ASAP7_75t_SL g294 ( .A(n_295), .B(n_297), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g306 ( .A(n_296), .B(n_307), .Y(n_306) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_305), .B1(n_309), .B2(n_312), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVx1_ASAP7_75t_L g373 ( .A(n_301), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_301), .B(n_341), .Y(n_408) );
AOI322xp5_ASAP7_75t_L g332 ( .A1(n_303), .A2(n_333), .A3(n_335), .B1(n_336), .B2(n_338), .C1(n_339), .C2(n_343), .Y(n_332) );
INVxp67_ASAP7_75t_L g326 ( .A(n_304), .Y(n_326) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_306), .A2(n_311), .B1(n_328), .B2(n_330), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_307), .B(n_320), .Y(n_407) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_308), .B(n_346), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_308), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g404 ( .A(n_310), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
NAND3xp33_ASAP7_75t_SL g315 ( .A(n_316), .B(n_332), .C(n_347), .Y(n_315) );
AOI221xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_318), .B1(n_323), .B2(n_325), .C(n_327), .Y(n_316) );
AND2x2_ASAP7_75t_L g323 ( .A(n_319), .B(n_324), .Y(n_323) );
INVx3_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
AND2x4_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
AND2x2_ASAP7_75t_L g333 ( .A(n_324), .B(n_334), .Y(n_333) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_326), .Y(n_405) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_331), .B(n_345), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_334), .B(n_392), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_335), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g410 ( .A(n_338), .Y(n_410) );
AND2x2_ASAP7_75t_L g425 ( .A(n_338), .B(n_402), .Y(n_425) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AOI211xp5_ASAP7_75t_L g419 ( .A1(n_349), .A2(n_420), .B(n_426), .C(n_434), .Y(n_419) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g388 ( .A(n_359), .B(n_389), .Y(n_388) );
NAND2x1_ASAP7_75t_SL g430 ( .A(n_360), .B(n_431), .Y(n_430) );
CKINVDCx16_ASAP7_75t_R g400 ( .A(n_363), .Y(n_400) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g395 ( .A(n_369), .Y(n_395) );
AND2x2_ASAP7_75t_L g399 ( .A(n_369), .B(n_385), .Y(n_399) );
NOR5xp2_ASAP7_75t_L g370 ( .A(n_371), .B(n_386), .C(n_403), .D(n_409), .E(n_412), .Y(n_370) );
OAI221xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_373), .B1(n_374), .B2(n_376), .C(n_378), .Y(n_371) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_375), .B(n_433), .Y(n_432) );
INVxp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g401 ( .A(n_385), .B(n_402), .Y(n_401) );
OAI221xp5_ASAP7_75t_SL g386 ( .A1(n_387), .A2(n_390), .B1(n_391), .B2(n_393), .C(n_396), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_399), .B1(n_400), .B2(n_401), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g439 ( .A(n_399), .Y(n_439) );
AOI211xp5_ASAP7_75t_SL g412 ( .A1(n_413), .A2(n_415), .B(n_417), .C(n_418), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_439), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
CKINVDCx14_ASAP7_75t_R g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g453 ( .A(n_448), .Y(n_453) );
NOR2x2_ASAP7_75t_L g754 ( .A(n_449), .B(n_753), .Y(n_754) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g752 ( .A(n_450), .B(n_753), .Y(n_752) );
NAND3xp33_ASAP7_75t_L g454 ( .A(n_452), .B(n_455), .C(n_758), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
CKINVDCx14_ASAP7_75t_R g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g756 ( .A(n_470), .Y(n_756) );
NAND2x1p5_ASAP7_75t_L g470 ( .A(n_471), .B(n_674), .Y(n_470) );
AND2x2_ASAP7_75t_SL g471 ( .A(n_472), .B(n_632), .Y(n_471) );
NOR4xp25_ASAP7_75t_L g472 ( .A(n_473), .B(n_572), .C(n_608), .D(n_622), .Y(n_472) );
OAI221xp5_ASAP7_75t_SL g473 ( .A1(n_474), .A2(n_520), .B1(n_550), .B2(n_559), .C(n_563), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g706 ( .A(n_474), .B(n_707), .Y(n_706) );
OR2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_500), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_488), .Y(n_476) );
AND2x2_ASAP7_75t_L g569 ( .A(n_477), .B(n_489), .Y(n_569) );
INVx3_ASAP7_75t_L g577 ( .A(n_477), .Y(n_577) );
AND2x2_ASAP7_75t_L g631 ( .A(n_477), .B(n_503), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_477), .B(n_502), .Y(n_667) );
AND2x2_ASAP7_75t_L g725 ( .A(n_477), .B(n_587), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B(n_486), .Y(n_482) );
INVx2_ASAP7_75t_L g496 ( .A(n_485), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_486), .A2(n_496), .B(n_510), .C(n_511), .Y(n_509) );
AND2x2_ASAP7_75t_L g560 ( .A(n_488), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g574 ( .A(n_488), .B(n_503), .Y(n_574) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_489), .B(n_503), .Y(n_589) );
AND2x2_ASAP7_75t_L g601 ( .A(n_489), .B(n_577), .Y(n_601) );
OR2x2_ASAP7_75t_L g603 ( .A(n_489), .B(n_561), .Y(n_603) );
AND2x2_ASAP7_75t_L g638 ( .A(n_489), .B(n_561), .Y(n_638) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_489), .Y(n_683) );
INVx1_ASAP7_75t_L g691 ( .A(n_489), .Y(n_691) );
OAI21xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_494), .B(n_498), .Y(n_490) );
OAI221xp5_ASAP7_75t_L g608 ( .A1(n_500), .A2(n_609), .B1(n_613), .B2(n_617), .C(n_618), .Y(n_608) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g568 ( .A(n_501), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_513), .Y(n_501) );
INVx2_ASAP7_75t_L g567 ( .A(n_502), .Y(n_567) );
AND2x2_ASAP7_75t_L g620 ( .A(n_502), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g639 ( .A(n_502), .B(n_577), .Y(n_639) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g702 ( .A(n_503), .B(n_577), .Y(n_702) );
AND2x2_ASAP7_75t_L g624 ( .A(n_513), .B(n_569), .Y(n_624) );
OAI322xp33_ASAP7_75t_L g692 ( .A1(n_513), .A2(n_648), .A3(n_693), .B1(n_695), .B2(n_698), .C1(n_700), .C2(n_704), .Y(n_692) );
INVx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NOR2x1_ASAP7_75t_L g575 ( .A(n_514), .B(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g588 ( .A(n_514), .Y(n_588) );
AND2x2_ASAP7_75t_L g697 ( .A(n_514), .B(n_577), .Y(n_697) );
AND2x2_ASAP7_75t_L g729 ( .A(n_514), .B(n_601), .Y(n_729) );
OR2x2_ASAP7_75t_L g732 ( .A(n_514), .B(n_733), .Y(n_732) );
AND2x4_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
INVx1_ASAP7_75t_L g562 ( .A(n_515), .Y(n_562) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_533), .Y(n_521) );
INVx1_ASAP7_75t_L g745 ( .A(n_522), .Y(n_745) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
OR2x2_ASAP7_75t_L g552 ( .A(n_523), .B(n_540), .Y(n_552) );
INVx2_ASAP7_75t_L g585 ( .A(n_523), .Y(n_585) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g607 ( .A(n_524), .Y(n_607) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_524), .Y(n_615) );
OR2x2_ASAP7_75t_L g739 ( .A(n_524), .B(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g564 ( .A(n_533), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g604 ( .A(n_533), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g656 ( .A(n_533), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_540), .Y(n_533) );
AND2x2_ASAP7_75t_L g553 ( .A(n_534), .B(n_554), .Y(n_553) );
NOR2xp67_ASAP7_75t_L g611 ( .A(n_534), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g665 ( .A(n_534), .B(n_555), .Y(n_665) );
OR2x2_ASAP7_75t_L g673 ( .A(n_534), .B(n_607), .Y(n_673) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx2_ASAP7_75t_L g582 ( .A(n_535), .Y(n_582) );
AND2x2_ASAP7_75t_L g592 ( .A(n_535), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g616 ( .A(n_535), .B(n_540), .Y(n_616) );
AND2x2_ASAP7_75t_L g680 ( .A(n_535), .B(n_555), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_540), .B(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_540), .B(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g593 ( .A(n_540), .Y(n_593) );
INVx1_ASAP7_75t_L g598 ( .A(n_540), .Y(n_598) );
AND2x2_ASAP7_75t_L g610 ( .A(n_540), .B(n_611), .Y(n_610) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_540), .Y(n_688) );
INVx1_ASAP7_75t_L g740 ( .A(n_540), .Y(n_740) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .B(n_545), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_553), .Y(n_550) );
AND2x2_ASAP7_75t_L g717 ( .A(n_551), .B(n_626), .Y(n_717) );
INVx2_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g644 ( .A(n_553), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g743 ( .A(n_553), .B(n_678), .Y(n_743) );
INVx1_ASAP7_75t_L g565 ( .A(n_554), .Y(n_565) );
AND2x2_ASAP7_75t_L g591 ( .A(n_554), .B(n_585), .Y(n_591) );
BUFx2_ASAP7_75t_L g650 ( .A(n_554), .Y(n_650) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_555), .Y(n_571) );
INVx1_ASAP7_75t_L g581 ( .A(n_555), .Y(n_581) );
NOR2xp67_ASAP7_75t_L g719 ( .A(n_559), .B(n_566), .Y(n_719) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AOI32xp33_ASAP7_75t_L g563 ( .A1(n_560), .A2(n_564), .A3(n_566), .B1(n_568), .B2(n_570), .Y(n_563) );
AND2x2_ASAP7_75t_L g703 ( .A(n_560), .B(n_576), .Y(n_703) );
AND2x2_ASAP7_75t_L g741 ( .A(n_560), .B(n_639), .Y(n_741) );
INVx1_ASAP7_75t_L g621 ( .A(n_561), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_565), .B(n_627), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_566), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_566), .B(n_569), .Y(n_617) );
NAND2xp5_ASAP7_75t_SL g720 ( .A(n_566), .B(n_638), .Y(n_720) );
OR2x2_ASAP7_75t_L g734 ( .A(n_566), .B(n_603), .Y(n_734) );
INVx3_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g661 ( .A(n_567), .B(n_569), .Y(n_661) );
OR2x2_ASAP7_75t_L g670 ( .A(n_567), .B(n_657), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_569), .B(n_620), .Y(n_642) );
INVx2_ASAP7_75t_L g657 ( .A(n_571), .Y(n_657) );
OR2x2_ASAP7_75t_L g672 ( .A(n_571), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g687 ( .A(n_571), .B(n_688), .Y(n_687) );
A2O1A1Ixp33_ASAP7_75t_L g744 ( .A1(n_571), .A2(n_664), .B(n_745), .C(n_746), .Y(n_744) );
OAI321xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_578), .A3(n_583), .B1(n_586), .B2(n_590), .C(n_594), .Y(n_572) );
INVx1_ASAP7_75t_L g685 ( .A(n_573), .Y(n_685) );
NAND2x1p5_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
AND2x2_ASAP7_75t_L g696 ( .A(n_574), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g648 ( .A(n_576), .Y(n_648) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_577), .B(n_691), .Y(n_708) );
OAI221xp5_ASAP7_75t_L g715 ( .A1(n_578), .A2(n_716), .B1(n_718), .B2(n_720), .C(n_721), .Y(n_715) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
AND2x2_ASAP7_75t_L g653 ( .A(n_580), .B(n_627), .Y(n_653) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_581), .B(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g626 ( .A(n_582), .Y(n_626) );
A2O1A1Ixp33_ASAP7_75t_L g668 ( .A1(n_583), .A2(n_624), .B(n_669), .C(n_671), .Y(n_668) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g635 ( .A(n_585), .B(n_592), .Y(n_635) );
BUFx2_ASAP7_75t_L g645 ( .A(n_585), .Y(n_645) );
INVx1_ASAP7_75t_L g660 ( .A(n_585), .Y(n_660) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
OR2x2_ASAP7_75t_L g666 ( .A(n_588), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g749 ( .A(n_588), .Y(n_749) );
INVx1_ASAP7_75t_L g742 ( .A(n_589), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
AND2x2_ASAP7_75t_L g595 ( .A(n_591), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g699 ( .A(n_591), .B(n_616), .Y(n_699) );
INVx1_ASAP7_75t_L g628 ( .A(n_592), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_599), .B1(n_602), .B2(n_604), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_596), .B(n_712), .Y(n_711) );
INVxp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x4_ASAP7_75t_L g664 ( .A(n_597), .B(n_665), .Y(n_664) );
BUFx3_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_SL g627 ( .A(n_598), .B(n_607), .Y(n_627) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g619 ( .A(n_601), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g629 ( .A(n_603), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
OAI221xp5_ASAP7_75t_L g723 ( .A1(n_606), .A2(n_724), .B1(n_726), .B2(n_727), .C(n_728), .Y(n_723) );
INVx1_ASAP7_75t_L g612 ( .A(n_607), .Y(n_612) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_607), .Y(n_678) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_610), .B(n_729), .Y(n_728) );
OAI21xp5_ASAP7_75t_L g618 ( .A1(n_611), .A2(n_616), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_614), .B(n_624), .Y(n_721) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g690 ( .A(n_615), .Y(n_690) );
AND2x2_ASAP7_75t_L g649 ( .A(n_616), .B(n_650), .Y(n_649) );
INVx2_ASAP7_75t_L g738 ( .A(n_616), .Y(n_738) );
INVx1_ASAP7_75t_L g654 ( .A(n_619), .Y(n_654) );
INVx1_ASAP7_75t_L g709 ( .A(n_620), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_625), .B1(n_628), .B2(n_629), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_626), .B(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g694 ( .A(n_627), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g731 ( .A(n_627), .B(n_665), .Y(n_731) );
OR2x2_ASAP7_75t_L g704 ( .A(n_628), .B(n_657), .Y(n_704) );
INVx1_ASAP7_75t_L g643 ( .A(n_629), .Y(n_643) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_631), .B(n_682), .Y(n_681) );
NOR3xp33_ASAP7_75t_L g632 ( .A(n_633), .B(n_651), .C(n_662), .Y(n_632) );
OAI211xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_636), .B(n_640), .C(n_646), .Y(n_633) );
INVxp67_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g705 ( .A1(n_635), .A2(n_706), .B1(n_710), .B2(n_713), .C(n_715), .Y(n_705) );
INVx1_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
AND2x2_ASAP7_75t_L g647 ( .A(n_638), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g701 ( .A(n_638), .B(n_702), .Y(n_701) );
OAI211xp5_ASAP7_75t_L g686 ( .A1(n_639), .A2(n_687), .B(n_689), .C(n_691), .Y(n_686) );
INVx2_ASAP7_75t_L g733 ( .A(n_639), .Y(n_733) );
OAI21xp5_ASAP7_75t_SL g640 ( .A1(n_641), .A2(n_643), .B(n_644), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g712 ( .A(n_645), .B(n_665), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .Y(n_646) );
OAI21xp5_ASAP7_75t_SL g651 ( .A1(n_652), .A2(n_654), .B(n_655), .Y(n_651) );
INVxp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OAI21xp5_ASAP7_75t_SL g655 ( .A1(n_656), .A2(n_658), .B(n_661), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_656), .B(n_685), .Y(n_684) );
INVxp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_661), .B(n_748), .Y(n_747) );
OAI21xp33_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_666), .B(n_668), .Y(n_662) );
INVx1_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g689 ( .A(n_665), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND4x1_ASAP7_75t_L g674 ( .A(n_675), .B(n_705), .C(n_722), .D(n_744), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_692), .Y(n_675) );
OAI211xp5_ASAP7_75t_SL g676 ( .A1(n_677), .A2(n_681), .B(n_684), .C(n_686), .Y(n_676) );
OR2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_680), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_691), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_703), .Y(n_700) );
INVx1_ASAP7_75t_L g726 ( .A(n_701), .Y(n_726) );
INVx2_ASAP7_75t_SL g714 ( .A(n_702), .Y(n_714) );
OR2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g727 ( .A(n_712), .Y(n_727) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NOR2xp33_ASAP7_75t_SL g722 ( .A(n_723), .B(n_730), .Y(n_722) );
INVx1_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
OAI221xp5_ASAP7_75t_SL g730 ( .A1(n_731), .A2(n_732), .B1(n_734), .B2(n_735), .C(n_736), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_741), .B1(n_742), .B2(n_743), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g737 ( .A(n_738), .B(n_739), .Y(n_737) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g757 ( .A(n_751), .Y(n_757) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_760), .Y(n_759) );
endmodule