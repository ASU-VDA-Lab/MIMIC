module fake_jpeg_14158_n_514 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_514);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_514;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_10),
.B(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVxp33_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_8),
.B(n_12),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_57),
.Y(n_130)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_59),
.Y(n_157)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_60),
.Y(n_187)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_61),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_14),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_62),
.B(n_82),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_63),
.Y(n_170)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_65),
.Y(n_185)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

CKINVDCx6p67_ASAP7_75t_R g125 ( 
.A(n_66),
.Y(n_125)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_67),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_68),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_69),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_71),
.Y(n_148)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_72),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_76),
.Y(n_161)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_79),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_26),
.B(n_14),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_81),
.B(n_86),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_0),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_47),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_83),
.Y(n_140)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_84),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_85),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_26),
.B(n_0),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_88),
.Y(n_168)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_89),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_45),
.B(n_13),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_90),
.B(n_100),
.Y(n_159)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_91),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_92),
.Y(n_176)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

BUFx12f_ASAP7_75t_SL g186 ( 
.A(n_93),
.Y(n_186)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

AOI21xp33_ASAP7_75t_L g96 ( 
.A1(n_45),
.A2(n_1),
.B(n_2),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_103),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_97),
.Y(n_179)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_98),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_99),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_49),
.B(n_12),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_21),
.Y(n_101)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_35),
.Y(n_102)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_37),
.B(n_2),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_21),
.Y(n_104)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

INVx11_ASAP7_75t_L g193 ( 
.A(n_106),
.Y(n_193)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_19),
.Y(n_107)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_107),
.Y(n_182)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_19),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_114),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_41),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_110),
.B(n_116),
.Y(n_198)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_111),
.B(n_112),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_21),
.Y(n_112)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_20),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_113),
.B(n_119),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_18),
.Y(n_114)
);

AND2x4_ASAP7_75t_L g115 ( 
.A(n_32),
.B(n_12),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_115),
.B(n_122),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_41),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_41),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_117),
.B(n_118),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_20),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_49),
.B(n_2),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_120),
.B(n_3),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_46),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_22),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_46),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_86),
.A2(n_25),
.B(n_53),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_123),
.B(n_126),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_103),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_118),
.A2(n_32),
.B1(n_55),
.B2(n_25),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_129),
.A2(n_138),
.B1(n_142),
.B2(n_173),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_59),
.A2(n_32),
.B1(n_21),
.B2(n_50),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_60),
.A2(n_55),
.B1(n_53),
.B2(n_50),
.Y(n_142)
);

NOR4xp25_ASAP7_75t_L g149 ( 
.A(n_81),
.B(n_52),
.C(n_24),
.D(n_29),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_149),
.B(n_154),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_152),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_83),
.B(n_52),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_66),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_155),
.B(n_169),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_115),
.A2(n_22),
.B1(n_42),
.B2(n_48),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_158),
.A2(n_190),
.B1(n_173),
.B2(n_189),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_114),
.B(n_34),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_112),
.B(n_34),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_171),
.B(n_177),
.Y(n_273)
);

O2A1O1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_115),
.A2(n_48),
.B(n_42),
.C(n_30),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_175),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_73),
.A2(n_30),
.B1(n_29),
.B2(n_27),
.Y(n_173)
);

INVx6_ASAP7_75t_SL g174 ( 
.A(n_121),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_174),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_85),
.B(n_27),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_87),
.B(n_24),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_178),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_97),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_180),
.A2(n_181),
.B1(n_184),
.B2(n_189),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_99),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_120),
.A2(n_68),
.B1(n_69),
.B2(n_65),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_183),
.A2(n_138),
.B1(n_142),
.B2(n_202),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_102),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_63),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_70),
.A2(n_39),
.B1(n_9),
.B2(n_11),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_191),
.A2(n_200),
.B1(n_140),
.B2(n_172),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_110),
.B(n_11),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_195),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_117),
.B(n_39),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_190),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_116),
.A2(n_39),
.B1(n_80),
.B2(n_71),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_76),
.B(n_81),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_204),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_167),
.A2(n_124),
.B1(n_133),
.B2(n_129),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_205),
.A2(n_209),
.B1(n_231),
.B2(n_234),
.Y(n_277)
);

BUFx12f_ASAP7_75t_L g207 ( 
.A(n_132),
.Y(n_207)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_207),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_211),
.A2(n_213),
.B1(n_239),
.B2(n_271),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_136),
.B(n_159),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_214),
.B(n_216),
.Y(n_275)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_130),
.Y(n_215)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_215),
.Y(n_284)
);

AO22x1_ASAP7_75t_SL g216 ( 
.A1(n_199),
.A2(n_156),
.B1(n_143),
.B2(n_136),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_217),
.Y(n_316)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_218),
.Y(n_297)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_132),
.Y(n_219)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_219),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_131),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_220),
.Y(n_289)
);

OA22x2_ASAP7_75t_L g221 ( 
.A1(n_183),
.A2(n_179),
.B1(n_197),
.B2(n_144),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_221),
.Y(n_321)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_176),
.Y(n_223)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_223),
.Y(n_313)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_128),
.Y(n_224)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_224),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_225),
.A2(n_232),
.B1(n_222),
.B2(n_210),
.Y(n_285)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_226),
.Y(n_288)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_160),
.Y(n_227)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_227),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_134),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_228),
.B(n_251),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_146),
.B(n_158),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_229),
.B(n_233),
.Y(n_311)
);

OA22x2_ASAP7_75t_L g230 ( 
.A1(n_147),
.A2(n_131),
.B1(n_137),
.B2(n_184),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_230),
.A2(n_240),
.B1(n_256),
.B2(n_261),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_196),
.A2(n_161),
.B1(n_148),
.B2(n_135),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_150),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_196),
.A2(n_148),
.B1(n_161),
.B2(n_135),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_139),
.B(n_192),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_235),
.B(n_244),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_203),
.Y(n_236)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_236),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_193),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_237),
.B(n_241),
.Y(n_309)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_141),
.Y(n_238)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_238),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_180),
.A2(n_181),
.B1(n_201),
.B2(n_170),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_153),
.A2(n_137),
.B1(n_186),
.B2(n_187),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_193),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_166),
.Y(n_242)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_242),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_141),
.B(n_168),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_243),
.B(n_266),
.C(n_216),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_163),
.B(n_168),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_162),
.Y(n_245)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_245),
.Y(n_310)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_247),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_163),
.B(n_162),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_248),
.B(n_252),
.Y(n_325)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_166),
.Y(n_249)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_249),
.Y(n_320)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_185),
.Y(n_250)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_250),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_186),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_185),
.B(n_201),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_194),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_253),
.B(n_254),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_127),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_194),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_255),
.B(n_260),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_153),
.A2(n_187),
.B1(n_157),
.B2(n_203),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_164),
.A2(n_145),
.B1(n_125),
.B2(n_151),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_257),
.A2(n_258),
.B1(n_236),
.B2(n_262),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_164),
.A2(n_145),
.B1(n_125),
.B2(n_157),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_176),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_259),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_127),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_165),
.A2(n_176),
.B1(n_125),
.B2(n_127),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_165),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_262),
.B(n_272),
.Y(n_301)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_165),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_263),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_193),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_264),
.B(n_207),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_136),
.B(n_159),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_126),
.A2(n_136),
.B1(n_103),
.B2(n_191),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_270),
.A2(n_229),
.B(n_211),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_153),
.A2(n_35),
.B1(n_31),
.B2(n_73),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_153),
.A2(n_35),
.B1(n_31),
.B2(n_73),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_235),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_274),
.B(n_276),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_268),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_278),
.A2(n_220),
.B1(n_226),
.B2(n_247),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_214),
.B(n_266),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_279),
.B(n_292),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_280),
.B(n_304),
.Y(n_326)
);

MAJx2_ASAP7_75t_L g283 ( 
.A(n_211),
.B(n_210),
.C(n_233),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_283),
.B(n_315),
.C(n_219),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_285),
.A2(n_287),
.B1(n_295),
.B2(n_280),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_225),
.A2(n_210),
.B1(n_212),
.B2(n_209),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_243),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_291),
.B(n_294),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_246),
.B(n_267),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_243),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_269),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_298),
.B(n_305),
.Y(n_358)
);

A2O1A1Ixp33_ASAP7_75t_L g302 ( 
.A1(n_216),
.A2(n_270),
.B(n_273),
.C(n_265),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_230),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_244),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_206),
.A2(n_265),
.B1(n_252),
.B2(n_221),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_306),
.A2(n_307),
.B1(n_277),
.B2(n_295),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_221),
.A2(n_248),
.B1(n_230),
.B2(n_208),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_208),
.B(n_218),
.C(n_215),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_236),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_317),
.B(n_281),
.Y(n_364)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_323),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_291),
.B(n_221),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_327),
.Y(n_391)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_324),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_330),
.B(n_352),
.Y(n_376)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_293),
.Y(n_331)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_331),
.Y(n_367)
);

NOR2x1_ASAP7_75t_L g332 ( 
.A(n_275),
.B(n_287),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_332),
.A2(n_335),
.B(n_339),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_312),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_333),
.B(n_345),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_305),
.B(n_325),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_334),
.B(n_338),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_307),
.A2(n_306),
.B1(n_321),
.B2(n_304),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_337),
.A2(n_348),
.B1(n_353),
.B2(n_355),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_325),
.B(n_230),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_275),
.B(n_263),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_293),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_303),
.Y(n_341)
);

MAJx2_ASAP7_75t_L g342 ( 
.A(n_283),
.B(n_242),
.C(n_249),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_342),
.B(n_344),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_274),
.B(n_250),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_343),
.B(n_354),
.Y(n_373)
);

O2A1O1Ixp33_ASAP7_75t_SL g345 ( 
.A1(n_321),
.A2(n_253),
.B(n_255),
.C(n_207),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_277),
.A2(n_217),
.B1(n_259),
.B2(n_223),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_346),
.A2(n_289),
.B1(n_316),
.B2(n_300),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_347),
.A2(n_357),
.B1(n_361),
.B2(n_327),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_309),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_349),
.Y(n_384)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_303),
.Y(n_350)
);

FAx1_ASAP7_75t_SL g352 ( 
.A(n_311),
.B(n_279),
.CI(n_319),
.CON(n_352),
.SN(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_311),
.A2(n_319),
.B1(n_285),
.B2(n_278),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_324),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_294),
.A2(n_302),
.B1(n_315),
.B2(n_282),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_301),
.A2(n_296),
.B1(n_276),
.B2(n_314),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_299),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_359),
.B(n_362),
.Y(n_383)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_322),
.Y(n_360)
);

NAND3xp33_ASAP7_75t_L g379 ( 
.A(n_360),
.B(n_288),
.C(n_318),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_301),
.A2(n_290),
.B1(n_292),
.B2(n_281),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_290),
.B(n_310),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_299),
.B(n_310),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_363),
.B(n_320),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_364),
.Y(n_377)
);

INVx13_ASAP7_75t_L g365 ( 
.A(n_331),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_365),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_366),
.A2(n_368),
.B1(n_372),
.B2(n_386),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_338),
.A2(n_316),
.B1(n_289),
.B2(n_300),
.Y(n_372)
);

AND2x6_ASAP7_75t_L g374 ( 
.A(n_352),
.B(n_308),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_374),
.B(n_380),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_348),
.A2(n_316),
.B1(n_284),
.B2(n_297),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_375),
.A2(n_387),
.B1(n_361),
.B2(n_357),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_336),
.B(n_351),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_378),
.B(n_286),
.Y(n_418)
);

HB1xp67_ASAP7_75t_SL g411 ( 
.A(n_379),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_363),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_332),
.A2(n_288),
.B(n_318),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_385),
.A2(n_339),
.B(n_356),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_347),
.A2(n_284),
.B1(n_320),
.B2(n_297),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_353),
.A2(n_335),
.B1(n_334),
.B2(n_355),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_388),
.B(n_389),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_352),
.B(n_313),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_362),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_390),
.B(n_392),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_343),
.B(n_333),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_384),
.Y(n_394)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_394),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_382),
.B(n_326),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_395),
.B(n_406),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_398),
.B(n_381),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_369),
.A2(n_330),
.B(n_332),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_401),
.A2(n_417),
.B(n_373),
.Y(n_436)
);

AO21x2_ASAP7_75t_L g402 ( 
.A1(n_385),
.A2(n_345),
.B(n_327),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_402),
.A2(n_404),
.B1(n_381),
.B2(n_386),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_380),
.B(n_358),
.Y(n_403)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_403),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_371),
.A2(n_326),
.B1(n_344),
.B2(n_345),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_405),
.A2(n_408),
.B1(n_414),
.B2(n_372),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_382),
.B(n_326),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_370),
.B(n_342),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_407),
.B(n_409),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_371),
.A2(n_328),
.B1(n_349),
.B2(n_339),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_366),
.B(n_342),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_388),
.Y(n_410)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_410),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_387),
.B(n_336),
.C(n_340),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_412),
.B(n_418),
.Y(n_423)
);

XNOR2x1_ASAP7_75t_L g413 ( 
.A(n_389),
.B(n_341),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_413),
.B(n_419),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_375),
.A2(n_350),
.B1(n_359),
.B2(n_354),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_384),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_415),
.B(n_377),
.Y(n_424)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_367),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_416),
.B(n_377),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_369),
.A2(n_313),
.B(n_329),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_370),
.B(n_286),
.Y(n_419)
);

NOR4xp25_ASAP7_75t_L g420 ( 
.A(n_403),
.B(n_390),
.C(n_392),
.D(n_391),
.Y(n_420)
);

NOR3xp33_ASAP7_75t_SL g446 ( 
.A(n_420),
.B(n_410),
.C(n_396),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_422),
.Y(n_444)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_424),
.Y(n_448)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_425),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_399),
.B(n_383),
.Y(n_426)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_426),
.Y(n_454)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_428),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_412),
.B(n_378),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_429),
.B(n_437),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_399),
.B(n_383),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_433),
.B(n_434),
.Y(n_450)
);

INVx6_ASAP7_75t_L g434 ( 
.A(n_411),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_417),
.B(n_376),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_435),
.A2(n_436),
.B(n_439),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_393),
.B(n_376),
.Y(n_437)
);

AND2x6_ASAP7_75t_L g440 ( 
.A(n_393),
.B(n_374),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_440),
.A2(n_402),
.B1(n_404),
.B2(n_401),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_407),
.B(n_374),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_441),
.B(n_405),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g442 ( 
.A(n_408),
.B(n_373),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_442),
.A2(n_398),
.B(n_396),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_432),
.B(n_395),
.C(n_406),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_445),
.B(n_447),
.C(n_457),
.Y(n_461)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_446),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_432),
.B(n_409),
.C(n_419),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_449),
.B(n_456),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_453),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_455),
.A2(n_435),
.B(n_436),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_438),
.B(n_413),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_438),
.B(n_402),
.Y(n_457)
);

FAx1_ASAP7_75t_L g458 ( 
.A(n_422),
.B(n_402),
.CI(n_397),
.CON(n_458),
.SN(n_458)
);

A2O1A1Ixp33_ASAP7_75t_SL g463 ( 
.A1(n_458),
.A2(n_425),
.B(n_442),
.C(n_420),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_431),
.B(n_400),
.C(n_367),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_459),
.B(n_445),
.C(n_447),
.Y(n_467)
);

INVx11_ASAP7_75t_L g462 ( 
.A(n_450),
.Y(n_462)
);

INVx11_ASAP7_75t_L g482 ( 
.A(n_462),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_463),
.A2(n_455),
.B(n_439),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_444),
.A2(n_435),
.B1(n_442),
.B2(n_427),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_467),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_460),
.B(n_423),
.Y(n_469)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_469),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_457),
.B(n_459),
.C(n_449),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_470),
.B(n_441),
.C(n_456),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_451),
.B(n_424),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_471),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_444),
.A2(n_427),
.B1(n_430),
.B2(n_426),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_472),
.A2(n_474),
.B(n_454),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_473),
.A2(n_452),
.B(n_448),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_443),
.A2(n_430),
.B1(n_433),
.B2(n_440),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_477),
.B(n_481),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_478),
.B(n_479),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_467),
.B(n_443),
.C(n_452),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_480),
.B(n_484),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_461),
.B(n_431),
.C(n_421),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_461),
.B(n_421),
.C(n_400),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_485),
.B(n_470),
.C(n_468),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_476),
.B(n_451),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_486),
.B(n_488),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_483),
.B(n_465),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_492),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_485),
.B(n_466),
.C(n_474),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_482),
.A2(n_462),
.B1(n_479),
.B2(n_473),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_493),
.B(n_494),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_475),
.A2(n_434),
.B1(n_458),
.B2(n_463),
.Y(n_494)
);

AOI21x1_ASAP7_75t_L g495 ( 
.A1(n_491),
.A2(n_480),
.B(n_446),
.Y(n_495)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_495),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_487),
.A2(n_482),
.B(n_477),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_496),
.B(n_497),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_492),
.Y(n_497)
);

NOR2xp67_ASAP7_75t_L g498 ( 
.A(n_490),
.B(n_481),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_498),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_500),
.B(n_489),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_502),
.B(n_506),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_497),
.B(n_490),
.C(n_463),
.Y(n_506)
);

OAI21xp33_ASAP7_75t_L g507 ( 
.A1(n_503),
.A2(n_499),
.B(n_504),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_507),
.B(n_509),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_505),
.B(n_501),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_508),
.Y(n_510)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_510),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_512),
.A2(n_511),
.B(n_505),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_513),
.B(n_472),
.Y(n_514)
);


endmodule