module fake_jpeg_26048_n_223 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_223);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_223;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_220;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_40),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_1),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_37),
.B(n_23),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_48),
.Y(n_75)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_53),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_40),
.B1(n_23),
.B2(n_18),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_47),
.A2(n_54),
.B1(n_17),
.B2(n_22),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_32),
.B1(n_31),
.B2(n_20),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_32),
.B1(n_31),
.B2(n_20),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_55),
.A2(n_17),
.B(n_22),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_30),
.B1(n_16),
.B2(n_25),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_56),
.A2(n_57),
.B1(n_16),
.B2(n_25),
.Y(n_87)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_30),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_38),
.Y(n_80)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_65),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_L g113 ( 
.A1(n_64),
.A2(n_94),
.B(n_27),
.Y(n_113)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_38),
.C(n_39),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_74),
.C(n_91),
.Y(n_107)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_69),
.Y(n_118)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_72),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_34),
.B1(n_57),
.B2(n_49),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_22),
.B1(n_17),
.B2(n_24),
.Y(n_98)
);

MAJx2_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_39),
.C(n_38),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_77),
.Y(n_105)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_82),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_93),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_26),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_81),
.B(n_84),
.Y(n_106)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_26),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_86),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_52),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_85),
.B(n_88),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_21),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_87),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_51),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_89),
.Y(n_119)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_92),
.B1(n_17),
.B2(n_24),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_36),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_66),
.A2(n_36),
.B1(n_21),
.B2(n_22),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_96),
.A2(n_98),
.B1(n_115),
.B2(n_116),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_1),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_103),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_2),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_3),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_4),
.Y(n_108)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_113),
.A2(n_68),
.B(n_90),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_87),
.A2(n_27),
.B1(n_6),
.B2(n_7),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_64),
.A2(n_27),
.B1(n_6),
.B2(n_7),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_62),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_120),
.A2(n_106),
.B1(n_101),
.B2(n_75),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_112),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_123),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_67),
.Y(n_123)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_74),
.Y(n_124)
);

A2O1A1O1Ixp25_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_104),
.B(n_103),
.C(n_100),
.D(n_95),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_81),
.B(n_93),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_125),
.A2(n_131),
.B(n_136),
.Y(n_145)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_127),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_119),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_132),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_96),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_116),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_119),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_140),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_79),
.Y(n_134)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

NOR2x1_ASAP7_75t_SL g136 ( 
.A(n_107),
.B(n_92),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_78),
.C(n_68),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_97),
.C(n_12),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_120),
.A2(n_69),
.B1(n_70),
.B2(n_10),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_139),
.A2(n_118),
.B1(n_10),
.B2(n_97),
.Y(n_155)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_10),
.B(n_11),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_142),
.A2(n_11),
.B(n_13),
.Y(n_162)
);

AO22x1_ASAP7_75t_SL g143 ( 
.A1(n_136),
.A2(n_115),
.B1(n_109),
.B2(n_98),
.Y(n_143)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_161),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_108),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_149),
.Y(n_177)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_152),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_95),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_148),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_129),
.A2(n_118),
.B(n_97),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_154),
.A2(n_159),
.B(n_162),
.Y(n_170)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_158),
.B(n_132),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_141),
.B(n_140),
.Y(n_159)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_167),
.B(n_169),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_146),
.B(n_126),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_160),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_171),
.A2(n_175),
.B(n_176),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_159),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_174),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_173),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_154),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_145),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_145),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_147),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_153),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_184),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_170),
.A2(n_159),
.B(n_150),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_164),
.Y(n_200)
);

INVxp33_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_186),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_152),
.C(n_157),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_171),
.C(n_170),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_165),
.A2(n_128),
.B1(n_139),
.B2(n_121),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_149),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_191),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_144),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_194),
.Y(n_207)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_190),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_167),
.C(n_177),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_198),
.C(n_184),
.Y(n_205)
);

NOR3xp33_ASAP7_75t_SL g199 ( 
.A(n_189),
.B(n_131),
.C(n_162),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_199),
.A2(n_122),
.B1(n_164),
.B2(n_165),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_172),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_201),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_202),
.A2(n_203),
.B(n_181),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_204),
.B(n_131),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_208),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_199),
.A2(n_182),
.B1(n_130),
.B2(n_155),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_207),
.A2(n_183),
.B(n_198),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_211),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_210),
.A2(n_202),
.B1(n_206),
.B2(n_133),
.Y(n_215)
);

AOI31xp67_ASAP7_75t_L g212 ( 
.A1(n_203),
.A2(n_143),
.A3(n_188),
.B(n_185),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_143),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_135),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_216),
.A2(n_214),
.B(n_142),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_213),
.C(n_192),
.Y(n_217)
);

NOR3xp33_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_197),
.C(n_191),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_218),
.A2(n_219),
.B(n_135),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_220),
.A2(n_221),
.B(n_197),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_192),
.B(n_137),
.Y(n_223)
);


endmodule