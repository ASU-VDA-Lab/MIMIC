module fake_jpeg_229_n_129 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_7),
.B(n_3),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_26),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_29),
.B(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_31)
);

AO22x1_ASAP7_75t_SL g48 ( 
.A1(n_31),
.A2(n_40),
.B1(n_24),
.B2(n_16),
.Y(n_48)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_32),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_23),
.A2(n_26),
.B1(n_14),
.B2(n_22),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_38),
.B1(n_43),
.B2(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_10),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_34),
.B(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_19),
.B(n_8),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_13),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_2),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_45),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_15),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_40)
);

CKINVDCx9p33_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_13),
.A2(n_5),
.B1(n_27),
.B2(n_17),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_27),
.B1(n_25),
.B2(n_17),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_45),
.B1(n_42),
.B2(n_46),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_24),
.B(n_18),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_12),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_20),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_52),
.Y(n_87)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_51),
.A2(n_69),
.B1(n_57),
.B2(n_49),
.Y(n_86)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_55),
.B(n_66),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_12),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_56),
.B(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_12),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_62),
.B(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_29),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_71),
.B1(n_50),
.B2(n_67),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_31),
.B(n_40),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_47),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_47),
.A2(n_37),
.B1(n_42),
.B2(n_36),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_34),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_57),
.Y(n_85)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_61),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_72),
.Y(n_95)
);

MAJx2_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_68),
.C(n_59),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_83),
.C(n_88),
.Y(n_96)
);

OA21x2_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_48),
.B(n_65),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_76),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_68),
.B(n_53),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_48),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_86),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_52),
.C(n_61),
.Y(n_83)
);

OA22x2_ASAP7_75t_SL g84 ( 
.A1(n_58),
.A2(n_64),
.B1(n_66),
.B2(n_68),
.Y(n_84)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

FAx1_ASAP7_75t_SL g92 ( 
.A(n_73),
.B(n_49),
.CI(n_76),
.CON(n_92),
.SN(n_92)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_87),
.B(n_74),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_93),
.B(n_94),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_75),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_96),
.B(n_97),
.Y(n_108)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_75),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_99),
.Y(n_103)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_74),
.B1(n_79),
.B2(n_87),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_101),
.A2(n_89),
.B1(n_96),
.B2(n_91),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_87),
.B(n_84),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_109),
.B(n_91),
.Y(n_112)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_104),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_99),
.B1(n_89),
.B2(n_98),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_116),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_109),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_113),
.C(n_115),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_112),
.A2(n_107),
.B(n_103),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_92),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_106),
.B(n_92),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_119),
.C(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_105),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_72),
.C(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

AOI321xp33_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_113),
.A3(n_121),
.B1(n_111),
.B2(n_115),
.C(n_109),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_124),
.C(n_86),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_121),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_125),
.A2(n_126),
.B1(n_101),
.B2(n_102),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_127),
.B(n_102),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_83),
.Y(n_129)
);


endmodule