module real_jpeg_7203_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_1),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_1),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_1),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_1),
.Y(n_204)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_1),
.Y(n_208)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_1),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_2),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_2),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_2),
.A2(n_47),
.B1(n_132),
.B2(n_220),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_2),
.A2(n_132),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_3),
.Y(n_84)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_3),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_3),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_4),
.A2(n_97),
.B1(n_101),
.B2(n_104),
.Y(n_96)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_4),
.Y(n_104)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_6),
.A2(n_35),
.B1(n_38),
.B2(n_42),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_6),
.A2(n_42),
.B1(n_267),
.B2(n_269),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_6),
.A2(n_42),
.B1(n_86),
.B2(n_283),
.Y(n_282)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_7),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_7),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_7),
.Y(n_155)
);

INVx8_ASAP7_75t_L g262 ( 
.A(n_7),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_7),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_8),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_8),
.B(n_53),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_8),
.A2(n_69),
.B1(n_241),
.B2(n_243),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_8),
.B(n_118),
.C(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_8),
.B(n_23),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_8),
.B(n_92),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_8),
.B(n_138),
.Y(n_288)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_10),
.Y(n_79)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_10),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g177 ( 
.A(n_10),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_11),
.A2(n_82),
.B1(n_85),
.B2(n_86),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_11),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_11),
.A2(n_85),
.B1(n_225),
.B2(n_228),
.Y(n_224)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_12),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_12),
.Y(n_118)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_12),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_13),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_13),
.A2(n_29),
.B1(n_51),
.B2(n_135),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_13),
.A2(n_51),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_13),
.A2(n_51),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_14),
.A2(n_124),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_14),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_234),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_232),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_163),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_18),
.B(n_163),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_107),
.C(n_139),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_19),
.A2(n_20),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_67),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_21),
.B(n_68),
.C(n_80),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_34),
.B(n_43),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_22),
.A2(n_34),
.B1(n_55),
.B2(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_22),
.B(n_45),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_23),
.B(n_56),
.Y(n_55)
);

AO22x2_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_26),
.B1(n_29),
.B2(n_31),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_26),
.Y(n_247)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_26),
.Y(n_268)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_27),
.Y(n_130)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_28),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_28),
.Y(n_147)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_28),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_30),
.Y(n_113)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_30),
.Y(n_227)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_30),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_30),
.Y(n_271)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_33),
.Y(n_151)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_54),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI32xp33_ASAP7_75t_L g140 ( 
.A1(n_47),
.A2(n_129),
.A3(n_141),
.B1(n_144),
.B2(n_145),
.Y(n_140)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_50),
.Y(n_311)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_54),
.A2(n_308),
.B(n_313),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_60),
.B1(n_63),
.B2(n_65),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_59),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_61),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_62),
.Y(n_180)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_80),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_69),
.B(n_182),
.Y(n_181)
);

OAI21xp33_ASAP7_75t_SL g206 ( 
.A1(n_69),
.A2(n_181),
.B(n_207),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_69),
.A2(n_185),
.B(n_259),
.Y(n_279)
);

OAI21xp33_ASAP7_75t_SL g308 ( 
.A1(n_69),
.A2(n_309),
.B(n_312),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_71),
.B(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_72),
.B(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_72)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_75),
.Y(n_170)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_78),
.Y(n_205)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_91),
.B1(n_96),
.B2(n_105),
.Y(n_80)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_81),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_82),
.Y(n_254)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx8_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_84),
.Y(n_258)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_91),
.B(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_91),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_91),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_96),
.Y(n_186)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_100),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_101),
.B(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_107),
.B(n_139),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_128),
.B(n_133),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_108),
.A2(n_133),
.B(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_108),
.A2(n_120),
.B1(n_128),
.B2(n_266),
.Y(n_305)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_109),
.B(n_134),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_120),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_114),
.B1(n_117),
.B2(n_119),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI22x1_ASAP7_75t_L g120 ( 
.A1(n_117),
.A2(n_121),
.B1(n_124),
.B2(n_126),
.Y(n_120)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_120),
.A2(n_224),
.B(n_230),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_120),
.A2(n_230),
.B(n_266),
.Y(n_265)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_127),
.Y(n_192)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_127),
.Y(n_250)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_138),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_152),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_140),
.B(n_152),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVxp33_ASAP7_75t_L g312 ( 
.A(n_144),
.Y(n_312)
);

NAND2xp33_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B(n_156),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_154),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_156),
.A2(n_282),
.B(n_285),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_157),
.B(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_196),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_164)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_183),
.B2(n_184),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI32xp33_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_171),
.A3(n_173),
.B1(n_175),
.B2(n_181),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_189),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_185),
.A2(n_253),
.B(n_259),
.Y(n_252)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_193),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_217),
.B2(n_231),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_206),
.B(n_209),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_200)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_223),
.Y(n_217)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AO21x1_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_316),
.B(n_321),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_300),
.B(n_315),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_274),
.B(n_299),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_251),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_238),
.B(n_251),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_245),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_239),
.A2(n_245),
.B1(n_246),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_239),
.Y(n_297)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_263),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_252),
.B(n_264),
.C(n_273),
.Y(n_301)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_253),
.Y(n_293)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_272),
.B2(n_273),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_290),
.B(n_298),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_280),
.B(n_289),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_288),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_288),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_296),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_296),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_302),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_314),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_306),
.C(n_314),
.Y(n_317)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_317),
.B(n_318),
.Y(n_321)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);


endmodule