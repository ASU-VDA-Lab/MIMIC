module real_aes_16192_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_733;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_0), .Y(n_551) );
AND2x4_ASAP7_75t_L g841 ( .A(n_1), .B(n_842), .Y(n_841) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_2), .A2(n_4), .B1(n_253), .B2(n_254), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_3), .A2(n_23), .B1(n_153), .B2(n_234), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_5), .A2(n_53), .B1(n_161), .B2(n_190), .Y(n_189) );
BUFx3_ASAP7_75t_L g585 ( .A(n_6), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g123 ( .A1(n_7), .A2(n_13), .B1(n_124), .B2(n_126), .Y(n_123) );
INVx1_ASAP7_75t_L g842 ( .A(n_8), .Y(n_842) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_9), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_10), .B(n_159), .Y(n_599) );
OR2x2_ASAP7_75t_L g105 ( .A(n_11), .B(n_33), .Y(n_105) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_12), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_14), .B(n_195), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g826 ( .A(n_15), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_16), .B(n_168), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_17), .A2(n_85), .B1(n_195), .B2(n_234), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g856 ( .A(n_18), .Y(n_856) );
OAI22xp5_ASAP7_75t_L g108 ( .A1(n_19), .A2(n_59), .B1(n_109), .B2(n_110), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_19), .Y(n_109) );
INVx1_ASAP7_75t_L g851 ( .A(n_20), .Y(n_851) );
OAI21x1_ASAP7_75t_L g136 ( .A1(n_21), .A2(n_49), .B(n_137), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_22), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_24), .B(n_153), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_25), .B(n_129), .Y(n_209) );
INVx4_ASAP7_75t_R g177 ( .A(n_26), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g852 ( .A(n_27), .Y(n_852) );
AO32x2_ASAP7_75t_L g510 ( .A1(n_28), .A2(n_147), .A3(n_148), .B1(n_511), .B2(n_514), .Y(n_510) );
AO32x1_ASAP7_75t_L g615 ( .A1(n_28), .A2(n_147), .A3(n_148), .B1(n_511), .B2(n_514), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_29), .B(n_153), .Y(n_216) );
INVx1_ASAP7_75t_L g258 ( .A(n_30), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_SL g231 ( .A1(n_31), .A2(n_124), .B(n_128), .C(n_232), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_32), .A2(n_46), .B1(n_124), .B2(n_131), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_34), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_35), .A2(n_52), .B1(n_153), .B2(n_178), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_36), .A2(n_90), .B1(n_131), .B2(n_234), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_37), .B(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_38), .B(n_523), .Y(n_527) );
INVx1_ASAP7_75t_L g213 ( .A(n_39), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_40), .B(n_124), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_41), .A2(n_68), .B1(n_131), .B2(n_536), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_42), .Y(n_151) );
INVx2_ASAP7_75t_L g840 ( .A(n_43), .Y(n_840) );
BUFx3_ASAP7_75t_L g104 ( .A(n_44), .Y(n_104) );
INVx1_ASAP7_75t_L g835 ( .A(n_44), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_45), .B(n_529), .Y(n_528) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_47), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_48), .A2(n_84), .B1(n_124), .B2(n_131), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_50), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g576 ( .A(n_51), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_54), .A2(n_78), .B1(n_197), .B2(n_523), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_55), .Y(n_142) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_56), .A2(n_82), .B1(n_195), .B2(n_234), .Y(n_581) );
INVx1_ASAP7_75t_L g137 ( .A(n_57), .Y(n_137) );
AND2x4_ASAP7_75t_L g139 ( .A(n_58), .B(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g110 ( .A(n_59), .Y(n_110) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_60), .A2(n_89), .B1(n_131), .B2(n_251), .Y(n_250) );
AO22x1_ASAP7_75t_L g193 ( .A1(n_61), .A2(n_73), .B1(n_194), .B2(n_196), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_62), .B(n_234), .Y(n_598) );
INVx1_ASAP7_75t_L g140 ( .A(n_63), .Y(n_140) );
AND2x2_ASAP7_75t_L g235 ( .A(n_64), .B(n_147), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_65), .B(n_147), .Y(n_604) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_66), .A2(n_161), .B(n_188), .C(n_550), .Y(n_549) );
NAND3xp33_ASAP7_75t_L g603 ( .A(n_67), .B(n_234), .C(n_602), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_69), .B(n_161), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_70), .Y(n_226) );
AND2x2_ASAP7_75t_L g552 ( .A(n_71), .B(n_182), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g539 ( .A(n_72), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_74), .B(n_153), .Y(n_152) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_75), .A2(n_95), .B1(n_195), .B2(n_197), .Y(n_574) );
INVx2_ASAP7_75t_L g129 ( .A(n_76), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_77), .B(n_154), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_79), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_80), .B(n_147), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g546 ( .A(n_81), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_83), .B(n_135), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_86), .B(n_602), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_87), .A2(n_99), .B1(n_131), .B2(n_178), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_88), .B(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_91), .B(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g501 ( .A(n_92), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_92), .B(n_834), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_93), .B(n_168), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g171 ( .A1(n_94), .A2(n_133), .B(n_161), .C(n_172), .Y(n_171) );
AND2x2_ASAP7_75t_L g181 ( .A(n_96), .B(n_182), .Y(n_181) );
NAND2xp33_ASAP7_75t_L g158 ( .A(n_97), .B(n_159), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_98), .Y(n_561) );
AOI211xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_829), .B(n_843), .C(n_864), .Y(n_100) );
OAI22xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_106), .B1(n_826), .B2(n_827), .Y(n_101) );
BUFx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g828 ( .A(n_103), .B(n_500), .Y(n_828) );
NOR2x1_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
INVx1_ASAP7_75t_L g836 ( .A(n_105), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_108), .B1(n_111), .B2(n_825), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g825 ( .A(n_111), .Y(n_825) );
AOI22x1_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_498), .B1(n_502), .B2(n_822), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
XNOR2x1_ASAP7_75t_L g849 ( .A(n_113), .B(n_850), .Y(n_849) );
AND2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_407), .Y(n_113) );
NOR3xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_323), .C(n_354), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_289), .Y(n_115) );
AOI211x1_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_201), .B(n_244), .C(n_275), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_165), .Y(n_118) );
AND2x2_ASAP7_75t_L g430 ( .A(n_119), .B(n_305), .Y(n_430) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_144), .Y(n_119) );
INVx1_ASAP7_75t_L g315 ( .A(n_120), .Y(n_315) );
OR2x2_ASAP7_75t_L g436 ( .A(n_120), .B(n_287), .Y(n_436) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g272 ( .A(n_121), .B(n_145), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_121), .B(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g304 ( .A(n_121), .Y(n_304) );
OR2x2_ASAP7_75t_L g335 ( .A(n_121), .B(n_166), .Y(n_335) );
AND2x2_ASAP7_75t_L g349 ( .A(n_121), .B(n_166), .Y(n_349) );
AND2x2_ASAP7_75t_L g386 ( .A(n_121), .B(n_342), .Y(n_386) );
AO31x2_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_134), .A3(n_138), .B(n_141), .Y(n_121) );
OAI22x1_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_127), .B1(n_130), .B2(n_132), .Y(n_122) );
INVx4_ASAP7_75t_L g126 ( .A(n_124), .Y(n_126) );
INVx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_125), .Y(n_131) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_125), .Y(n_153) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_125), .Y(n_159) );
INVx1_ASAP7_75t_L g161 ( .A(n_125), .Y(n_161) );
INVx1_ASAP7_75t_L g173 ( .A(n_125), .Y(n_173) );
INVx1_ASAP7_75t_L g178 ( .A(n_125), .Y(n_178) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_125), .Y(n_195) );
INVx1_ASAP7_75t_L g197 ( .A(n_125), .Y(n_197) );
INVx1_ASAP7_75t_L g228 ( .A(n_125), .Y(n_228) );
INVx2_ASAP7_75t_L g234 ( .A(n_125), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g150 ( .A1(n_126), .A2(n_151), .B(n_152), .C(n_154), .Y(n_150) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_127), .A2(n_187), .B1(n_239), .B2(n_240), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_127), .A2(n_132), .B1(n_250), .B2(n_252), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_127), .A2(n_527), .B(n_528), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_127), .A2(n_187), .B1(n_535), .B2(n_537), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_127), .A2(n_572), .B1(n_573), .B2(n_574), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_127), .A2(n_128), .B1(n_581), .B2(n_582), .Y(n_580) );
INVx6_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_128), .A2(n_158), .B(n_160), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_128), .B(n_193), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g288 ( .A1(n_128), .A2(n_186), .B(n_193), .C(n_199), .Y(n_288) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_128), .A2(n_230), .B1(n_512), .B2(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_128), .A2(n_598), .B(n_599), .Y(n_597) );
BUFx8_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g133 ( .A(n_129), .Y(n_133) );
INVx2_ASAP7_75t_L g156 ( .A(n_129), .Y(n_156) );
INVx1_ASAP7_75t_L g212 ( .A(n_129), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_131), .B(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g253 ( .A(n_131), .Y(n_253) );
INVx2_ASAP7_75t_L g525 ( .A(n_131), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_132), .B(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g548 ( .A(n_133), .Y(n_548) );
INVx1_ASAP7_75t_SL g573 ( .A(n_133), .Y(n_573) );
INVx2_ASAP7_75t_L g595 ( .A(n_134), .Y(n_595) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g143 ( .A(n_135), .Y(n_143) );
INVx2_ASAP7_75t_L g169 ( .A(n_135), .Y(n_169) );
OAI21xp33_ASAP7_75t_L g199 ( .A1(n_135), .A2(n_191), .B(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_136), .Y(n_148) );
INVx2_ASAP7_75t_L g180 ( .A(n_138), .Y(n_180) );
BUFx10_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx10_ASAP7_75t_L g164 ( .A(n_139), .Y(n_164) );
INVx1_ASAP7_75t_L g200 ( .A(n_139), .Y(n_200) );
INVx1_ASAP7_75t_L g256 ( .A(n_139), .Y(n_256) );
AO31x2_ASAP7_75t_L g532 ( .A1(n_139), .A2(n_533), .A3(n_534), .B(n_538), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
INVx2_ASAP7_75t_L g182 ( .A(n_143), .Y(n_182) );
BUFx2_ASAP7_75t_L g222 ( .A(n_143), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_143), .B(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_143), .B(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_143), .B(n_576), .Y(n_575) );
BUFx2_ASAP7_75t_L g266 ( .A(n_144), .Y(n_266) );
AND2x2_ASAP7_75t_L g317 ( .A(n_144), .B(n_183), .Y(n_317) );
AND2x2_ASAP7_75t_L g460 ( .A(n_144), .B(n_166), .Y(n_460) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
BUFx3_ASAP7_75t_L g284 ( .A(n_145), .Y(n_284) );
AND2x2_ASAP7_75t_L g303 ( .A(n_145), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g340 ( .A(n_145), .Y(n_340) );
AND2x2_ASAP7_75t_L g364 ( .A(n_145), .B(n_166), .Y(n_364) );
NAND2x1p5_ASAP7_75t_L g145 ( .A(n_146), .B(n_149), .Y(n_145) );
NOR2x1_ASAP7_75t_L g162 ( .A(n_147), .B(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g241 ( .A(n_147), .Y(n_241) );
INVx4_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x2_ASAP7_75t_L g217 ( .A(n_148), .B(n_164), .Y(n_217) );
INVx2_ASAP7_75t_SL g519 ( .A(n_148), .Y(n_519) );
BUFx3_ASAP7_75t_L g533 ( .A(n_148), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_148), .B(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g558 ( .A(n_148), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_148), .B(n_584), .Y(n_583) );
OAI21x1_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_157), .B(n_162), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_153), .B(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g536 ( .A(n_153), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_153), .A2(n_178), .B1(n_546), .B2(n_547), .Y(n_545) );
INVx2_ASAP7_75t_SL g154 ( .A(n_155), .Y(n_154) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_155), .A2(n_564), .B1(n_565), .B2(n_566), .Y(n_563) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx3_ASAP7_75t_L g188 ( .A(n_156), .Y(n_188) );
OAI22xp33_ASAP7_75t_L g176 ( .A1(n_159), .A2(n_177), .B1(n_178), .B2(n_179), .Y(n_176) );
INVx2_ASAP7_75t_L g251 ( .A(n_159), .Y(n_251) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AO31x2_ASAP7_75t_L g237 ( .A1(n_164), .A2(n_238), .A3(n_241), .B(n_242), .Y(n_237) );
OAI21x1_ASAP7_75t_L g559 ( .A1(n_164), .A2(n_560), .B(n_563), .Y(n_559) );
AOI31xp67_ASAP7_75t_L g579 ( .A1(n_164), .A2(n_241), .A3(n_580), .B(n_583), .Y(n_579) );
OAI21x1_ASAP7_75t_L g596 ( .A1(n_164), .A2(n_597), .B(n_600), .Y(n_596) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_165), .Y(n_264) );
AND2x2_ASAP7_75t_L g325 ( .A(n_165), .B(n_314), .Y(n_325) );
INVx2_ASAP7_75t_L g457 ( .A(n_165), .Y(n_457) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_183), .Y(n_165) );
INVx1_ASAP7_75t_L g262 ( .A(n_166), .Y(n_262) );
AND2x4_ASAP7_75t_L g274 ( .A(n_166), .B(n_184), .Y(n_274) );
INVx2_ASAP7_75t_L g342 ( .A(n_166), .Y(n_342) );
AO21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_170), .B(n_181), .Y(n_166) );
AOI21x1_ASAP7_75t_L g542 ( .A1(n_167), .A2(n_543), .B(n_552), .Y(n_542) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_175), .B(n_180), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
INVx2_ASAP7_75t_L g190 ( .A(n_173), .Y(n_190) );
INVx1_ASAP7_75t_L g565 ( .A(n_178), .Y(n_565) );
AND2x2_ASAP7_75t_L g341 ( .A(n_183), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g348 ( .A(n_183), .Y(n_348) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g426 ( .A(n_184), .B(n_342), .Y(n_426) );
AOI21x1_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_192), .B(n_198), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
OAI21x1_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_189), .B(n_191), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_187), .A2(n_215), .B(n_216), .Y(n_214) );
AOI21x1_ASAP7_75t_L g521 ( .A1(n_187), .A2(n_522), .B(n_524), .Y(n_521) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVxp67_ASAP7_75t_SL g194 ( .A(n_195), .Y(n_194) );
INVx3_ASAP7_75t_L g529 ( .A(n_195), .Y(n_529) );
OAI21xp33_ASAP7_75t_SL g208 ( .A1(n_196), .A2(n_209), .B(n_210), .Y(n_208) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_197), .B(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_200), .A2(n_224), .B(n_231), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_200), .A2(n_544), .B(n_549), .Y(n_543) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_203), .B(n_218), .Y(n_202) );
OR2x2_ASAP7_75t_L g331 ( .A(n_203), .B(n_219), .Y(n_331) );
AND2x2_ASAP7_75t_L g469 ( .A(n_203), .B(n_413), .Y(n_469) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x4_ASAP7_75t_L g246 ( .A(n_204), .B(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g351 ( .A(n_204), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_204), .B(n_293), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_204), .B(n_269), .Y(n_406) );
INVx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g263 ( .A(n_205), .Y(n_263) );
AND2x2_ASAP7_75t_L g279 ( .A(n_205), .B(n_280), .Y(n_279) );
NAND2x1p5_ASAP7_75t_SL g292 ( .A(n_205), .B(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g300 ( .A(n_205), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_205), .B(n_269), .Y(n_371) );
AND2x2_ASAP7_75t_L g419 ( .A(n_205), .B(n_248), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_205), .B(n_247), .Y(n_462) );
BUFx2_ASAP7_75t_L g481 ( .A(n_205), .Y(n_481) );
AND2x4_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
OAI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_214), .B(n_217), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
BUFx4f_ASAP7_75t_L g230 ( .A(n_212), .Y(n_230) );
INVx1_ASAP7_75t_L g602 ( .A(n_212), .Y(n_602) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
OR2x2_ASAP7_75t_L g265 ( .A(n_219), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g378 ( .A(n_219), .Y(n_378) );
OR2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_236), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_220), .B(n_248), .Y(n_281) );
INVx2_ASAP7_75t_L g293 ( .A(n_220), .Y(n_293) );
AND2x2_ASAP7_75t_L g329 ( .A(n_220), .B(n_237), .Y(n_329) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g269 ( .A(n_221), .Y(n_269) );
AOI21x1_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_235), .Y(n_221) );
AO31x2_ASAP7_75t_L g248 ( .A1(n_222), .A2(n_249), .A3(n_255), .B(n_257), .Y(n_248) );
OAI21xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_227), .B(n_230), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
INVx2_ASAP7_75t_L g254 ( .A(n_228), .Y(n_254) );
O2A1O1Ixp5_ASAP7_75t_L g560 ( .A1(n_230), .A2(n_254), .B(n_561), .C(n_562), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
INVx2_ASAP7_75t_SL g523 ( .A(n_234), .Y(n_523) );
INVx1_ASAP7_75t_L g353 ( .A(n_236), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_236), .B(n_248), .Y(n_370) );
INVx2_ASAP7_75t_SL g236 ( .A(n_237), .Y(n_236) );
BUFx2_ASAP7_75t_L g280 ( .A(n_237), .Y(n_280) );
OR2x2_ASAP7_75t_L g312 ( .A(n_237), .B(n_248), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_237), .B(n_248), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_265), .B1(n_267), .B2(n_271), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_259), .B1(n_263), .B2(n_264), .Y(n_245) );
INVx2_ASAP7_75t_L g270 ( .A(n_246), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_246), .B(n_329), .Y(n_343) );
AND2x2_ASAP7_75t_L g377 ( .A(n_246), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g295 ( .A(n_248), .Y(n_295) );
INVx1_ASAP7_75t_L g301 ( .A(n_248), .Y(n_301) );
AO31x2_ASAP7_75t_L g570 ( .A1(n_255), .A2(n_533), .A3(n_571), .B(n_575), .Y(n_570) );
INVx2_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
INVx2_ASAP7_75t_SL g514 ( .A(n_256), .Y(n_514) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g435 ( .A(n_261), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g316 ( .A(n_262), .Y(n_316) );
AND3x1_ASAP7_75t_L g420 ( .A(n_262), .B(n_283), .C(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g376 ( .A(n_263), .Y(n_376) );
AND2x4_ASAP7_75t_L g412 ( .A(n_263), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g450 ( .A(n_266), .Y(n_450) );
INVx1_ASAP7_75t_L g454 ( .A(n_267), .Y(n_454) );
OR2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
OR2x2_ASAP7_75t_L g427 ( .A(n_268), .B(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_SL g475 ( .A(n_268), .Y(n_475) );
INVxp67_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g375 ( .A(n_269), .B(n_353), .Y(n_375) );
AND2x2_ASAP7_75t_L g417 ( .A(n_269), .B(n_284), .Y(n_417) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_269), .Y(n_421) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_272), .B(n_273), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_L g336 ( .A1(n_272), .A2(n_273), .B(n_337), .C(n_343), .Y(n_336) );
NAND2x1_ASAP7_75t_L g380 ( .A(n_272), .B(n_381), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_272), .B(n_430), .Y(n_476) );
INVx3_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_274), .B(n_303), .Y(n_322) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_277), .B(n_282), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVx2_ASAP7_75t_L g298 ( .A(n_280), .Y(n_298) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_281), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_282), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
AND2x2_ASAP7_75t_L g332 ( .A(n_283), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_283), .B(n_349), .Y(n_396) );
NAND2x1p5_ASAP7_75t_L g402 ( .A(n_283), .B(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_283), .B(n_341), .Y(n_497) );
INVx3_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx2_ASAP7_75t_L g480 ( .A(n_284), .Y(n_480) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g306 ( .A(n_287), .Y(n_306) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_302), .B(n_307), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_296), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
OAI33xp33_ASAP7_75t_L g356 ( .A1(n_292), .A2(n_297), .A3(n_357), .B1(n_358), .B2(n_360), .B3(n_361), .Y(n_356) );
OR2x2_ASAP7_75t_L g488 ( .A(n_292), .B(n_312), .Y(n_488) );
INVx2_ASAP7_75t_L g490 ( .A(n_292), .Y(n_490) );
INVx1_ASAP7_75t_L g311 ( .A(n_293), .Y(n_311) );
OR2x2_ASAP7_75t_L g352 ( .A(n_293), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
INVx1_ASAP7_75t_L g360 ( .A(n_297), .Y(n_360) );
NOR3xp33_ASAP7_75t_L g478 ( .A(n_297), .B(n_479), .C(n_481), .Y(n_478) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_298), .B(n_438), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_298), .B(n_462), .Y(n_466) );
AND2x4_ASAP7_75t_L g495 ( .A(n_298), .B(n_496), .Y(n_495) );
INVxp67_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g321 ( .A(n_300), .Y(n_321) );
OR2x2_ASAP7_75t_L g327 ( .A(n_300), .B(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g440 ( .A(n_300), .B(n_375), .Y(n_440) );
INVx1_ASAP7_75t_L g496 ( .A(n_300), .Y(n_496) );
AND2x4_ASAP7_75t_SL g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx1_ASAP7_75t_L g319 ( .A(n_303), .Y(n_319) );
INVx1_ASAP7_75t_L g362 ( .A(n_304), .Y(n_362) );
AND2x2_ASAP7_75t_L g403 ( .A(n_304), .B(n_306), .Y(n_403) );
INVx1_ASAP7_75t_L g443 ( .A(n_305), .Y(n_443) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g334 ( .A(n_306), .B(n_335), .Y(n_334) );
OAI22xp33_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_313), .B1(n_320), .B2(n_322), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx2_ASAP7_75t_L g399 ( .A(n_312), .Y(n_399) );
INVx2_ASAP7_75t_L g413 ( .A(n_312), .Y(n_413) );
AOI211xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_316), .B(n_317), .C(n_318), .Y(n_313) );
INVx1_ASAP7_75t_L g357 ( .A(n_314), .Y(n_357) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_315), .B(n_340), .Y(n_442) );
OR2x2_ASAP7_75t_L g458 ( .A(n_315), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g471 ( .A(n_315), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_317), .B(n_385), .Y(n_446) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g323 ( .A(n_324), .B(n_344), .Y(n_323) );
AOI221xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_326), .B1(n_330), .B2(n_332), .C(n_336), .Y(n_324) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OAI32xp33_ASAP7_75t_L g493 ( .A1(n_327), .A2(n_424), .A3(n_442), .B1(n_494), .B2(n_497), .Y(n_493) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g463 ( .A(n_329), .Y(n_463) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OAI21xp5_ASAP7_75t_L g344 ( .A1(n_332), .A2(n_345), .B(n_350), .Y(n_344) );
NAND2x1_ASAP7_75t_L g492 ( .A(n_333), .B(n_480), .Y(n_492) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g367 ( .A(n_335), .Y(n_367) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
AND2x2_ASAP7_75t_L g486 ( .A(n_339), .B(n_367), .Y(n_486) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g434 ( .A(n_340), .Y(n_434) );
INVx2_ASAP7_75t_L g387 ( .A(n_341), .Y(n_387) );
INVx2_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
AND2x2_ASAP7_75t_L g363 ( .A(n_347), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g382 ( .A(n_348), .Y(n_382) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NAND4xp25_ASAP7_75t_L g354 ( .A(n_355), .B(n_372), .C(n_383), .D(n_394), .Y(n_354) );
AOI22xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_363), .B1(n_365), .B2(n_368), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_357), .A2(n_485), .B1(n_487), .B2(n_488), .Y(n_484) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g467 ( .A(n_362), .B(n_426), .Y(n_467) );
AND2x2_ASAP7_75t_L g470 ( .A(n_364), .B(n_471), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_365), .A2(n_384), .B1(n_388), .B2(n_391), .Y(n_383) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
OR2x2_ASAP7_75t_L g405 ( .A(n_370), .B(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g389 ( .A(n_371), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g400 ( .A(n_371), .Y(n_400) );
OAI21xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_377), .B(n_379), .Y(n_372) );
O2A1O1Ixp33_ASAP7_75t_L g477 ( .A1(n_373), .A2(n_478), .B(n_482), .C(n_484), .Y(n_477) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
INVxp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g452 ( .A(n_375), .Y(n_452) );
AND2x4_ASAP7_75t_L g445 ( .A(n_378), .B(n_419), .Y(n_445) );
INVx2_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
OAI21xp33_ASAP7_75t_L g410 ( .A1(n_385), .A2(n_411), .B(n_414), .Y(n_410) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g416 ( .A(n_386), .B(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_386), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g392 ( .A(n_390), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_392), .A2(n_423), .B1(n_427), .B2(n_429), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_397), .B1(n_401), .B2(n_404), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_399), .Y(n_415) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_472), .Y(n_407) );
NAND4xp25_ASAP7_75t_L g408 ( .A(n_409), .B(n_431), .C(n_447), .D(n_464), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_422), .Y(n_409) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g474 ( .A(n_412), .B(n_475), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_416), .B1(n_418), .B2(n_420), .Y(n_414) );
INVxp67_ASAP7_75t_L g438 ( .A(n_418), .Y(n_438) );
BUFx2_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g428 ( .A(n_419), .Y(n_428) );
AND2x2_ASAP7_75t_L g451 ( .A(n_419), .B(n_452), .Y(n_451) );
INVx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_437), .B(n_439), .Y(n_431) );
NOR2x1_ASAP7_75t_L g432 ( .A(n_433), .B(n_435), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OR2x6_ASAP7_75t_L g456 ( .A(n_434), .B(n_457), .Y(n_456) );
INVx3_ASAP7_75t_L g453 ( .A(n_435), .Y(n_453) );
OAI32xp33_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .A3(n_443), .B1(n_444), .B2(n_446), .Y(n_439) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AOI221xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_451), .B1(n_453), .B2(n_454), .C(n_455), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_458), .B(n_461), .Y(n_455) );
INVx2_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
OR2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
NOR2x1_ASAP7_75t_L g464 ( .A(n_465), .B(n_468), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
INVx1_ASAP7_75t_L g487 ( .A(n_466), .Y(n_487) );
INVx1_ASAP7_75t_L g483 ( .A(n_467), .Y(n_483) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
OAI211xp5_ASAP7_75t_SL g472 ( .A1(n_473), .A2(n_476), .B(n_477), .C(n_489), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVxp67_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
AOI21xp33_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_491), .B(n_493), .Y(n_489) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_499), .Y(n_498) );
BUFx8_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g824 ( .A(n_500), .Y(n_824) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx2_ASAP7_75t_L g848 ( .A(n_501), .Y(n_848) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NOR2x1p5_ASAP7_75t_L g503 ( .A(n_504), .B(n_730), .Y(n_503) );
NAND4xp75_ASAP7_75t_L g504 ( .A(n_505), .B(n_627), .C(n_661), .D(n_710), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_553), .B(n_586), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_515), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g706 ( .A(n_509), .Y(n_706) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g591 ( .A(n_510), .B(n_517), .Y(n_591) );
AND2x4_ASAP7_75t_L g622 ( .A(n_510), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g643 ( .A(n_510), .Y(n_643) );
OAI21x1_ASAP7_75t_L g520 ( .A1(n_514), .A2(n_521), .B(n_526), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_515), .B(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_531), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_516), .B(n_657), .Y(n_734) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_516), .Y(n_761) );
OR2x2_ASAP7_75t_L g810 ( .A(n_516), .B(n_614), .Y(n_810) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g626 ( .A(n_517), .Y(n_626) );
INVx3_ASAP7_75t_L g634 ( .A(n_517), .Y(n_634) );
OR2x2_ASAP7_75t_L g642 ( .A(n_517), .B(n_643), .Y(n_642) );
OR2x2_ASAP7_75t_L g670 ( .A(n_517), .B(n_640), .Y(n_670) );
INVx1_ASAP7_75t_L g681 ( .A(n_517), .Y(n_681) );
AND2x2_ASAP7_75t_L g702 ( .A(n_517), .B(n_643), .Y(n_702) );
INVxp67_ASAP7_75t_L g726 ( .A(n_517), .Y(n_726) );
BUFx2_ASAP7_75t_L g770 ( .A(n_517), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_517), .B(n_532), .Y(n_779) );
AND2x2_ASAP7_75t_L g786 ( .A(n_517), .B(n_787), .Y(n_786) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
OAI21x1_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B(n_530), .Y(n_518) );
OAI21xp5_ASAP7_75t_L g600 ( .A1(n_525), .A2(n_601), .B(n_603), .Y(n_600) );
AND2x2_ASAP7_75t_L g644 ( .A(n_531), .B(n_645), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g798 ( .A1(n_531), .A2(n_556), .B1(n_760), .B2(n_799), .Y(n_798) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_540), .Y(n_531) );
OR2x2_ASAP7_75t_L g614 ( .A(n_532), .B(n_615), .Y(n_614) );
INVx3_ASAP7_75t_L g623 ( .A(n_532), .Y(n_623) );
AND2x2_ASAP7_75t_L g635 ( .A(n_532), .B(n_615), .Y(n_635) );
AND2x2_ASAP7_75t_L g693 ( .A(n_532), .B(n_541), .Y(n_693) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g590 ( .A(n_541), .Y(n_590) );
INVx1_ASAP7_75t_L g684 ( .A(n_541), .Y(n_684) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_541), .Y(n_787) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g640 ( .A(n_542), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_545), .B(n_548), .Y(n_544) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_568), .Y(n_554) );
AND2x2_ASAP7_75t_L g741 ( .A(n_555), .B(n_687), .Y(n_741) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AOI32xp33_ASAP7_75t_L g771 ( .A1(n_556), .A2(n_664), .A3(n_738), .B1(n_772), .B2(n_774), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_556), .B(n_801), .Y(n_800) );
INVx2_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
OR2x2_ASAP7_75t_L g593 ( .A(n_557), .B(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g610 ( .A(n_557), .B(n_570), .Y(n_610) );
BUFx2_ASAP7_75t_L g629 ( .A(n_557), .Y(n_629) );
INVx1_ASAP7_75t_L g676 ( .A(n_557), .Y(n_676) );
AND2x2_ASAP7_75t_L g709 ( .A(n_557), .B(n_688), .Y(n_709) );
OA21x2_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B(n_567), .Y(n_557) );
OA21x2_ASAP7_75t_L g655 ( .A1(n_558), .A2(n_559), .B(n_567), .Y(n_655) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g592 ( .A(n_569), .B(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g797 ( .A(n_569), .B(n_681), .Y(n_797) );
INVx1_ASAP7_75t_L g801 ( .A(n_569), .Y(n_801) );
OR2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_577), .Y(n_569) );
INVx2_ASAP7_75t_L g625 ( .A(n_570), .Y(n_625) );
AND2x2_ASAP7_75t_L g649 ( .A(n_570), .B(n_608), .Y(n_649) );
AND2x2_ASAP7_75t_L g660 ( .A(n_570), .B(n_655), .Y(n_660) );
INVx1_ASAP7_75t_L g667 ( .A(n_570), .Y(n_667) );
AND2x2_ASAP7_75t_L g675 ( .A(n_570), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g688 ( .A(n_570), .Y(n_688) );
AND2x2_ASAP7_75t_L g754 ( .A(n_570), .B(n_577), .Y(n_754) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g618 ( .A(n_578), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g608 ( .A(n_579), .Y(n_608) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_585), .Y(n_584) );
OAI221xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_592), .B1(n_605), .B2(n_611), .C(n_616), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OAI21xp5_ASAP7_75t_L g737 ( .A1(n_588), .A2(n_738), .B(n_741), .Y(n_737) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
AND2x4_ASAP7_75t_L g813 ( .A(n_589), .B(n_613), .Y(n_813) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x4_ASAP7_75t_L g657 ( .A(n_590), .B(n_623), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_591), .B(n_692), .Y(n_691) );
BUFx2_ASAP7_75t_L g722 ( .A(n_591), .Y(n_722) );
OR2x2_ASAP7_75t_L g666 ( .A(n_593), .B(n_667), .Y(n_666) );
OR2x2_ASAP7_75t_L g728 ( .A(n_593), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g799 ( .A(n_593), .Y(n_799) );
AND2x2_ASAP7_75t_L g607 ( .A(n_594), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g756 ( .A(n_594), .B(n_655), .Y(n_756) );
OAI21xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B(n_604), .Y(n_594) );
OAI21x1_ASAP7_75t_L g619 ( .A1(n_595), .A2(n_596), .B(n_604), .Y(n_619) );
OAI221xp5_ASAP7_75t_L g636 ( .A1(n_605), .A2(n_637), .B1(n_638), .B2(n_647), .C(n_656), .Y(n_636) );
OAI221xp5_ASAP7_75t_L g732 ( .A1(n_605), .A2(n_720), .B1(n_733), .B2(n_735), .C(n_737), .Y(n_732) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
AND2x2_ASAP7_75t_L g659 ( .A(n_607), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g672 ( .A(n_608), .B(n_655), .Y(n_672) );
INVx2_ASAP7_75t_L g678 ( .A(n_608), .Y(n_678) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OAI221xp5_ASAP7_75t_L g742 ( .A1(n_611), .A2(n_743), .B1(n_748), .B2(n_752), .C(n_757), .Y(n_742) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g794 ( .A(n_614), .B(n_764), .Y(n_794) );
INVx1_ASAP7_75t_L g646 ( .A(n_615), .Y(n_646) );
INVx1_ASAP7_75t_L g683 ( .A(n_615), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_620), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g632 ( .A(n_618), .Y(n_632) );
OR2x2_ASAP7_75t_L g695 ( .A(n_618), .B(n_631), .Y(n_695) );
INVx2_ASAP7_75t_L g708 ( .A(n_618), .Y(n_708) );
INVx2_ASAP7_75t_L g653 ( .A(n_619), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_624), .Y(n_620) );
INVx3_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
BUFx2_ASAP7_75t_L g658 ( .A(n_622), .Y(n_658) );
AND2x4_ASAP7_75t_L g664 ( .A(n_622), .B(n_665), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_622), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g738 ( .A(n_622), .B(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g815 ( .A(n_622), .B(n_770), .Y(n_815) );
AND2x2_ASAP7_75t_L g639 ( .A(n_623), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g701 ( .A(n_623), .Y(n_701) );
INVx1_ASAP7_75t_L g760 ( .A(n_623), .Y(n_760) );
OR2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
INVx2_ASAP7_75t_SL g631 ( .A(n_625), .Y(n_631) );
AND2x2_ASAP7_75t_L g673 ( .A(n_625), .B(n_652), .Y(n_673) );
AND2x2_ASAP7_75t_L g747 ( .A(n_626), .B(n_701), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_633), .B(n_636), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx1_ASAP7_75t_L g713 ( .A(n_629), .Y(n_713) );
AND2x2_ASAP7_75t_L g780 ( .A(n_629), .B(n_708), .Y(n_780) );
AND2x2_ASAP7_75t_L g795 ( .A(n_629), .B(n_754), .Y(n_795) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
INVx2_ASAP7_75t_L g749 ( .A(n_631), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_631), .B(n_756), .Y(n_766) );
OAI33xp33_ASAP7_75t_L g803 ( .A1(n_631), .A2(n_705), .A3(n_773), .B1(n_804), .B2(n_805), .B3(n_806), .Y(n_803) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_634), .B(n_640), .Y(n_764) );
AND2x2_ASAP7_75t_L g792 ( .A(n_635), .B(n_740), .Y(n_792) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_641), .B(n_644), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g665 ( .A(n_640), .Y(n_665) );
INVx1_ASAP7_75t_L g740 ( .A(n_640), .Y(n_740) );
OAI32xp33_ASAP7_75t_L g685 ( .A1(n_641), .A2(n_666), .A3(n_686), .B1(n_689), .B2(n_691), .Y(n_685) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g720 ( .A(n_642), .B(n_665), .Y(n_720) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g698 ( .A(n_646), .Y(n_698) );
INVx2_ASAP7_75t_L g746 ( .A(n_646), .Y(n_746) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x4_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
INVx2_ASAP7_75t_L g729 ( .A(n_649), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_650), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g789 ( .A(n_650), .B(n_736), .Y(n_789) );
INVx2_ASAP7_75t_L g820 ( .A(n_650), .Y(n_820) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g735 ( .A(n_651), .B(n_736), .Y(n_735) );
NAND2x1p5_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
AND2x2_ASAP7_75t_L g677 ( .A(n_652), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g719 ( .A(n_653), .Y(n_719) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI21xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_658), .B(n_659), .Y(n_656) );
INVx2_ASAP7_75t_L g727 ( .A(n_657), .Y(n_727) );
AND2x2_ASAP7_75t_L g711 ( .A(n_658), .B(n_712), .Y(n_711) );
NOR3x1_ASAP7_75t_L g661 ( .A(n_662), .B(n_685), .C(n_694), .Y(n_661) );
OAI21xp5_ASAP7_75t_SL g662 ( .A1(n_663), .A2(n_666), .B(n_668), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g806 ( .A(n_665), .B(n_807), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_667), .B(n_718), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_671), .B1(n_674), .B2(n_679), .Y(n_668) );
INVx3_ASAP7_75t_L g703 ( .A(n_670), .Y(n_703) );
AND2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVxp67_ASAP7_75t_L g716 ( .A(n_672), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_672), .B(n_751), .Y(n_750) );
AND2x4_ASAP7_75t_L g674 ( .A(n_675), .B(n_677), .Y(n_674) );
AND2x2_ASAP7_75t_L g817 ( .A(n_675), .B(n_708), .Y(n_817) );
AND2x2_ASAP7_75t_L g687 ( .A(n_678), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g736 ( .A(n_678), .Y(n_736) );
INVx1_ASAP7_75t_L g773 ( .A(n_678), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_678), .B(n_719), .Y(n_807) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NAND2x1p5_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
INVx1_ASAP7_75t_L g804 ( .A(n_682), .Y(n_804) );
AND2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx1_ASAP7_75t_L g690 ( .A(n_684), .Y(n_690) );
AND2x2_ASAP7_75t_L g816 ( .A(n_687), .B(n_756), .Y(n_816) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
BUFx2_ASAP7_75t_L g724 ( .A(n_693), .Y(n_724) );
AND2x2_ASAP7_75t_L g821 ( .A(n_693), .B(n_702), .Y(n_821) );
OAI22xp33_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B1(n_704), .B2(n_707), .Y(n_694) );
AOI211xp5_ASAP7_75t_SL g696 ( .A1(n_697), .A2(n_699), .B(n_702), .C(n_703), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OR2x2_ASAP7_75t_L g778 ( .A(n_698), .B(n_779), .Y(n_778) );
INVxp67_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVxp33_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
AND2x2_ASAP7_75t_L g712 ( .A(n_708), .B(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g790 ( .A(n_709), .B(n_751), .Y(n_790) );
INVx1_ASAP7_75t_L g805 ( .A(n_709), .Y(n_805) );
NOR3xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_714), .C(n_721), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_720), .Y(n_714) );
OR2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g751 ( .A(n_719), .Y(n_751) );
O2A1O1Ixp33_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B(n_725), .C(n_728), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_722), .A2(n_815), .B1(n_816), .B2(n_817), .Y(n_814) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OR2x2_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_782), .Y(n_730) );
NOR3xp33_ASAP7_75t_SL g731 ( .A(n_732), .B(n_742), .C(n_767), .Y(n_731) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_738), .A2(n_777), .B1(n_780), .B2(n_781), .Y(n_776) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_747), .Y(n_744) );
AND2x2_ASAP7_75t_L g762 ( .A(n_745), .B(n_763), .Y(n_762) );
AND2x4_ASAP7_75t_L g785 ( .A(n_745), .B(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OR2x2_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
INVx1_ASAP7_75t_L g781 ( .A(n_750), .Y(n_781) );
OR2x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_755), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_756), .B(n_773), .Y(n_775) );
OAI21xp5_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_762), .B(n_765), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_759), .B(n_761), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g818 ( .A1(n_762), .A2(n_817), .B1(n_819), .B2(n_821), .Y(n_818) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
OAI21xp33_ASAP7_75t_SL g767 ( .A1(n_768), .A2(n_771), .B(n_776), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_769), .B(n_813), .Y(n_812) );
BUFx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g808 ( .A(n_779), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_781), .A2(n_803), .B1(n_808), .B2(n_809), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_811), .Y(n_782) );
OAI211xp5_ASAP7_75t_SL g783 ( .A1(n_784), .A2(n_788), .B(n_791), .C(n_802), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
NOR2x1_ASAP7_75t_L g788 ( .A(n_789), .B(n_790), .Y(n_788) );
O2A1O1Ixp5_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_793), .B(n_795), .C(n_796), .Y(n_791) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_794), .A2(n_797), .B1(n_798), .B2(n_800), .Y(n_796) );
OAI211xp5_ASAP7_75t_L g811 ( .A1(n_805), .A2(n_812), .B(n_814), .C(n_818), .Y(n_811) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx8_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
BUFx12f_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_830), .B(n_837), .Y(n_829) );
INVx3_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
CKINVDCx8_ASAP7_75t_R g831 ( .A(n_832), .Y(n_831) );
INVx5_ASAP7_75t_L g855 ( .A(n_832), .Y(n_855) );
INVx3_ASAP7_75t_L g869 ( .A(n_832), .Y(n_869) );
AND2x6_ASAP7_75t_SL g832 ( .A(n_833), .B(n_836), .Y(n_832) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
HB1xp67_ASAP7_75t_L g847 ( .A(n_835), .Y(n_847) );
AND3x2_ASAP7_75t_L g846 ( .A(n_836), .B(n_847), .C(n_848), .Y(n_846) );
NAND2xp5_ASAP7_75t_SL g837 ( .A(n_838), .B(n_841), .Y(n_837) );
BUFx2_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
NOR2xp33_ASAP7_75t_L g861 ( .A(n_839), .B(n_862), .Y(n_861) );
INVx3_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_840), .B(n_869), .Y(n_868) );
INVx2_ASAP7_75t_SL g863 ( .A(n_841), .Y(n_863) );
AOI21xp33_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_853), .B(n_857), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_845), .B(n_849), .Y(n_844) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
XOR2xp5_ASAP7_75t_L g850 ( .A(n_851), .B(n_852), .Y(n_850) );
NOR2xp33_ASAP7_75t_L g864 ( .A(n_852), .B(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_855), .B(n_856), .Y(n_854) );
CKINVDCx20_ASAP7_75t_R g857 ( .A(n_858), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g858 ( .A(n_859), .Y(n_858) );
INVx4_ASAP7_75t_SL g859 ( .A(n_860), .Y(n_859) );
BUFx3_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
OR2x4_ASAP7_75t_L g867 ( .A(n_862), .B(n_868), .Y(n_867) );
BUFx2_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
INVx4_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
BUFx3_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
endmodule