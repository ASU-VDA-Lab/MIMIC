module fake_jpeg_29266_n_102 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_102);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_35),
.Y(n_43)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_48),
.Y(n_57)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_49),
.A2(n_44),
.B1(n_39),
.B2(n_43),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_41),
.B1(n_33),
.B2(n_43),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_53),
.B1(n_58),
.B2(n_59),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_33),
.B1(n_41),
.B2(n_37),
.Y(n_53)
);

AO21x1_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_47),
.B(n_18),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_39),
.B1(n_42),
.B2(n_34),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_42),
.B1(n_34),
.B2(n_40),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_36),
.B1(n_1),
.B2(n_2),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_47),
.C(n_16),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_10),
.C(n_12),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_63),
.A2(n_52),
.B1(n_8),
.B2(n_9),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_0),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_70),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_13),
.B1(n_14),
.B2(n_19),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_59),
.B1(n_54),
.B2(n_50),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_68),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_3),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_69),
.B(n_7),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_4),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_12),
.B(n_13),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_52),
.B1(n_55),
.B2(n_22),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_72),
.A2(n_76),
.B1(n_78),
.B2(n_81),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_72),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_77),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_68),
.B1(n_67),
.B2(n_63),
.Y(n_78)
);

NOR3xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_20),
.C(n_23),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_61),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_85),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_65),
.Y(n_85)
);

NAND3xp33_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_88),
.C(n_24),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_74),
.A2(n_64),
.B(n_26),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_88),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_90),
.B(n_83),
.Y(n_93)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_92),
.C(n_77),
.Y(n_96)
);

XNOR2x1_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_95),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_95),
.B(n_86),
.C(n_87),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_78),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_94),
.C(n_82),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_73),
.Y(n_101)
);

OAI222xp33_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.C1(n_31),
.C2(n_32),
.Y(n_102)
);


endmodule