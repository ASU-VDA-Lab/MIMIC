module fake_netlist_5_804_n_617 (n_91, n_82, n_122, n_10, n_24, n_124, n_86, n_83, n_61, n_90, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_105, n_80, n_4, n_125, n_35, n_73, n_17, n_92, n_19, n_120, n_30, n_5, n_33, n_14, n_84, n_23, n_29, n_79, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_617);

input n_91;
input n_82;
input n_122;
input n_10;
input n_24;
input n_124;
input n_86;
input n_83;
input n_61;
input n_90;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_30;
input n_5;
input n_33;
input n_14;
input n_84;
input n_23;
input n_29;
input n_79;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_617;

wire n_137;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_611;
wire n_444;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_418;
wire n_248;
wire n_136;
wire n_146;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_408;
wire n_376;
wire n_503;
wire n_127;
wire n_235;
wire n_226;
wire n_605;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_483;
wire n_544;
wire n_155;
wire n_552;
wire n_547;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_139;
wire n_280;
wire n_590;
wire n_378;
wire n_551;
wire n_581;
wire n_382;
wire n_554;
wire n_254;
wire n_583;
wire n_302;
wire n_265;
wire n_526;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_455;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_606;
wire n_559;
wire n_275;
wire n_252;
wire n_295;
wire n_133;
wire n_330;
wire n_508;
wire n_506;
wire n_610;
wire n_509;
wire n_568;
wire n_147;
wire n_373;
wire n_307;
wire n_439;
wire n_150;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_134;
wire n_191;
wire n_587;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_320;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_132;
wire n_546;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_152;
wire n_540;
wire n_317;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_131;
wire n_192;
wire n_600;
wire n_223;
wire n_392;
wire n_158;
wire n_138;
wire n_264;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_347;
wire n_169;
wire n_550;
wire n_522;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_459;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_386;
wire n_578;
wire n_344;
wire n_287;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_415;
wire n_141;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_336;
wire n_584;
wire n_591;
wire n_145;
wire n_521;
wire n_614;
wire n_337;
wire n_430;
wire n_313;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_140;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_613;
wire n_241;
wire n_357;
wire n_598;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_144;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_129;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_309;
wire n_512;
wire n_462;
wire n_130;
wire n_322;
wire n_567;
wire n_258;
wire n_151;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_474;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_489;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_365;
wire n_176;
wire n_557;
wire n_182;
wire n_143;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_180;
wire n_560;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_572;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_269;
wire n_529;
wire n_128;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_135;
wire n_126;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_426;
wire n_565;
wire n_520;
wire n_409;
wire n_589;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_541;
wire n_391;
wire n_434;
wire n_539;
wire n_175;
wire n_538;
wire n_262;
wire n_238;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_324;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_424;
wire n_256;
wire n_305;
wire n_533;
wire n_278;

OR2x2_ASAP7_75t_L g126 ( 
.A(n_6),
.B(n_43),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_17),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_70),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_5),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_118),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_99),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_76),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_8),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_22),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_71),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_81),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_124),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_89),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_80),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_100),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_84),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_2),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_58),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_42),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_41),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_20),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_69),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_25),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_105),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_83),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_49),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_3),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_14),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_103),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_50),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_74),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_110),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_123),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_37),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_2),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_30),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_38),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_5),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_120),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_56),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_31),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_113),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_77),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_102),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_40),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_9),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_28),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_39),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_0),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_0),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_45),
.Y(n_184)
);

NOR2xp67_ASAP7_75t_L g185 ( 
.A(n_87),
.B(n_46),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_95),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_109),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_63),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_108),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_93),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_36),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_16),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_130),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_149),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_1),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_R g196 ( 
.A1(n_179),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_4),
.Y(n_197)
);

OAI21x1_ASAP7_75t_L g198 ( 
.A1(n_143),
.A2(n_57),
.B(n_119),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

AND2x4_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_6),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

OAI21x1_ASAP7_75t_L g205 ( 
.A1(n_181),
.A2(n_55),
.B(n_117),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_165),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_157),
.B(n_7),
.Y(n_208)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

AOI22x1_ASAP7_75t_SL g210 ( 
.A1(n_136),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_210)
);

CKINVDCx11_ASAP7_75t_R g211 ( 
.A(n_168),
.Y(n_211)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_128),
.Y(n_213)
);

OAI22x1_ASAP7_75t_R g214 ( 
.A1(n_163),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_163),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_132),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_127),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_189),
.Y(n_219)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_129),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_131),
.Y(n_223)
);

OA21x2_ASAP7_75t_L g224 ( 
.A1(n_135),
.A2(n_13),
.B(n_15),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_164),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_164),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_139),
.B(n_144),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_145),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_146),
.Y(n_229)
);

AND2x4_ASAP7_75t_L g230 ( 
.A(n_150),
.B(n_27),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_151),
.Y(n_231)
);

AND2x4_ASAP7_75t_L g232 ( 
.A(n_162),
.B(n_29),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_172),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_173),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_176),
.Y(n_235)
);

CKINVDCx11_ASAP7_75t_R g236 ( 
.A(n_178),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_216),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_221),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_199),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_230),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_236),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_212),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_222),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_222),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_223),
.Y(n_252)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_223),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_223),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_230),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_223),
.Y(n_256)
);

NAND3xp33_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_126),
.C(n_192),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_232),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_202),
.B(n_147),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_234),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_229),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_197),
.B(n_178),
.Y(n_263)
);

OR2x6_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_185),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_206),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_229),
.Y(n_266)
);

AOI21x1_ASAP7_75t_L g267 ( 
.A1(n_227),
.A2(n_191),
.B(n_184),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_229),
.Y(n_268)
);

AND3x2_ASAP7_75t_L g269 ( 
.A(n_203),
.B(n_219),
.C(n_208),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_229),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_204),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_213),
.B(n_134),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_235),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_232),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_212),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_203),
.B(n_166),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_236),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_204),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_212),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_218),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_235),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_235),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_202),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_209),
.B(n_167),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_235),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_217),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_260),
.B(n_193),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_245),
.B(n_255),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_245),
.B(n_220),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_260),
.B(n_226),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_239),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_257),
.B(n_225),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_245),
.B(n_255),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_239),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_263),
.B(n_209),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_255),
.B(n_220),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_259),
.B(n_220),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_238),
.B(n_207),
.Y(n_298)
);

NOR3xp33_ASAP7_75t_L g299 ( 
.A(n_238),
.B(n_208),
.C(n_211),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_264),
.A2(n_215),
.B1(n_133),
.B2(n_142),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_259),
.B(n_274),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_280),
.Y(n_302)
);

NOR2xp67_ASAP7_75t_SL g303 ( 
.A(n_274),
.B(n_224),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_244),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_228),
.Y(n_305)
);

BUFx6f_ASAP7_75t_SL g306 ( 
.A(n_264),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_244),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_265),
.Y(n_308)
);

BUFx8_ASAP7_75t_L g309 ( 
.A(n_271),
.Y(n_309)
);

NAND3xp33_ASAP7_75t_L g310 ( 
.A(n_271),
.B(n_195),
.C(n_233),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_269),
.B(n_276),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_283),
.B(n_140),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_278),
.B(n_194),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_278),
.B(n_194),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_264),
.B(n_195),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_241),
.B(n_137),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_249),
.B(n_224),
.Y(n_317)
);

NAND2xp33_ASAP7_75t_L g318 ( 
.A(n_249),
.B(n_138),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_284),
.B(n_141),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_279),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_237),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_264),
.B(n_148),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_237),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_285),
.B(n_152),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_265),
.Y(n_325)
);

AO221x1_ASAP7_75t_L g326 ( 
.A1(n_237),
.A2(n_196),
.B1(n_224),
.B2(n_214),
.C(n_210),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_279),
.B(n_153),
.Y(n_327)
);

NAND3xp33_ASAP7_75t_L g328 ( 
.A(n_258),
.B(n_154),
.C(n_155),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_285),
.B(n_156),
.Y(n_329)
);

AOI221xp5_ASAP7_75t_L g330 ( 
.A1(n_240),
.A2(n_175),
.B1(n_158),
.B2(n_177),
.C(n_188),
.Y(n_330)
);

OR2x6_ASAP7_75t_L g331 ( 
.A(n_275),
.B(n_205),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_247),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_247),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_275),
.B(n_180),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_253),
.B(n_187),
.Y(n_335)
);

BUFx5_ASAP7_75t_L g336 ( 
.A(n_242),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_237),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_237),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_261),
.B(n_186),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_253),
.B(n_174),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_253),
.B(n_169),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_267),
.B(n_161),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_240),
.B(n_198),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_248),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_248),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_320),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_330),
.B(n_267),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_334),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_288),
.B(n_282),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_302),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_304),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_317),
.A2(n_282),
.B(n_281),
.Y(n_352)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_345),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_293),
.B(n_250),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g355 ( 
.A1(n_315),
.A2(n_281),
.B1(n_251),
.B2(n_273),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_301),
.A2(n_273),
.B(n_270),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_342),
.A2(n_254),
.B(n_270),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_311),
.A2(n_290),
.B1(n_292),
.B2(n_322),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_313),
.B(n_251),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_289),
.A2(n_268),
.B(n_266),
.Y(n_360)
);

AOI21x1_ASAP7_75t_L g361 ( 
.A1(n_303),
.A2(n_268),
.B(n_266),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_307),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_314),
.B(n_211),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_312),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_343),
.A2(n_252),
.B(n_262),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_345),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_308),
.B(n_277),
.Y(n_367)
);

NAND3xp33_ASAP7_75t_L g368 ( 
.A(n_310),
.B(n_242),
.C(n_243),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_325),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_295),
.B(n_277),
.Y(n_370)
);

O2A1O1Ixp5_ASAP7_75t_L g371 ( 
.A1(n_305),
.A2(n_262),
.B(n_256),
.C(n_254),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_332),
.Y(n_372)
);

AOI21x1_ASAP7_75t_L g373 ( 
.A1(n_296),
.A2(n_256),
.B(n_252),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_297),
.A2(n_243),
.B(n_32),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_336),
.B(n_33),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_316),
.A2(n_34),
.B(n_35),
.Y(n_376)
);

A2O1A1Ixp33_ASAP7_75t_L g377 ( 
.A1(n_286),
.A2(n_246),
.B(n_47),
.C(n_48),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_333),
.Y(n_378)
);

AO21x2_ASAP7_75t_L g379 ( 
.A1(n_324),
.A2(n_44),
.B(n_51),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_309),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_291),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_336),
.B(n_52),
.Y(n_382)
);

OR2x6_ASAP7_75t_L g383 ( 
.A(n_298),
.B(n_246),
.Y(n_383)
);

AO21x1_ASAP7_75t_L g384 ( 
.A1(n_319),
.A2(n_53),
.B(n_54),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_327),
.B(n_59),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_329),
.A2(n_60),
.B(n_61),
.Y(n_386)
);

BUFx4f_ASAP7_75t_L g387 ( 
.A(n_344),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_331),
.A2(n_65),
.B(n_66),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_287),
.B(n_67),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_336),
.B(n_72),
.Y(n_390)
);

A2O1A1Ixp33_ASAP7_75t_L g391 ( 
.A1(n_300),
.A2(n_73),
.B(n_75),
.C(n_78),
.Y(n_391)
);

CKINVDCx8_ASAP7_75t_R g392 ( 
.A(n_326),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_294),
.Y(n_393)
);

A2O1A1Ixp33_ASAP7_75t_L g394 ( 
.A1(n_300),
.A2(n_79),
.B(n_82),
.C(n_85),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_306),
.A2(n_86),
.B1(n_88),
.B2(n_90),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_R g396 ( 
.A(n_318),
.B(n_94),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_335),
.B(n_341),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_340),
.A2(n_96),
.B(n_97),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_328),
.B(n_98),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_365),
.A2(n_347),
.B(n_352),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_358),
.B(n_323),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_392),
.B(n_306),
.Y(n_402)
);

OAI21x1_ASAP7_75t_L g403 ( 
.A1(n_361),
.A2(n_337),
.B(n_321),
.Y(n_403)
);

A2O1A1Ixp33_ASAP7_75t_L g404 ( 
.A1(n_389),
.A2(n_299),
.B(n_339),
.C(n_338),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_350),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_363),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_348),
.B(n_309),
.Y(n_407)
);

A2O1A1Ixp33_ASAP7_75t_L g408 ( 
.A1(n_397),
.A2(n_101),
.B(n_104),
.C(n_106),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_351),
.B(n_107),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_387),
.B(n_111),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_365),
.A2(n_112),
.B(n_115),
.Y(n_411)
);

A2O1A1Ixp33_ASAP7_75t_L g412 ( 
.A1(n_388),
.A2(n_116),
.B(n_122),
.C(n_369),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_371),
.A2(n_349),
.B(n_354),
.Y(n_413)
);

AO31x2_ASAP7_75t_L g414 ( 
.A1(n_384),
.A2(n_391),
.A3(n_394),
.B(n_382),
.Y(n_414)
);

OAI21x1_ASAP7_75t_L g415 ( 
.A1(n_356),
.A2(n_357),
.B(n_360),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_359),
.A2(n_353),
.B(n_387),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_353),
.A2(n_375),
.B(n_390),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_362),
.B(n_378),
.Y(n_418)
);

OAI21x1_ASAP7_75t_L g419 ( 
.A1(n_381),
.A2(n_355),
.B(n_393),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_346),
.Y(n_420)
);

AOI221xp5_ASAP7_75t_SL g421 ( 
.A1(n_385),
.A2(n_399),
.B1(n_377),
.B2(n_374),
.C(n_398),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_367),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_372),
.Y(n_423)
);

AOI21xp33_ASAP7_75t_L g424 ( 
.A1(n_370),
.A2(n_364),
.B(n_383),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_368),
.A2(n_386),
.B(n_376),
.Y(n_425)
);

O2A1O1Ixp5_ASAP7_75t_L g426 ( 
.A1(n_395),
.A2(n_379),
.B(n_396),
.C(n_366),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_383),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_366),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_383),
.B(n_380),
.Y(n_429)
);

AOI21x1_ASAP7_75t_L g430 ( 
.A1(n_379),
.A2(n_303),
.B(n_361),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_351),
.Y(n_431)
);

AO31x2_ASAP7_75t_L g432 ( 
.A1(n_384),
.A2(n_315),
.A3(n_358),
.B(n_391),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_351),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_351),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_431),
.B(n_434),
.Y(n_435)
);

NAND2x1p5_ASAP7_75t_L g436 ( 
.A(n_405),
.B(n_410),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_L g437 ( 
.A1(n_433),
.A2(n_423),
.B1(n_411),
.B2(n_418),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_422),
.B(n_400),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_419),
.Y(n_439)
);

INVx8_ASAP7_75t_L g440 ( 
.A(n_405),
.Y(n_440)
);

AO21x2_ASAP7_75t_L g441 ( 
.A1(n_425),
.A2(n_413),
.B(n_411),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_401),
.Y(n_442)
);

OAI21x1_ASAP7_75t_L g443 ( 
.A1(n_415),
.A2(n_403),
.B(n_417),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_422),
.B(n_424),
.Y(n_444)
);

BUFx2_ASAP7_75t_SL g445 ( 
.A(n_420),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_405),
.B(n_416),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_406),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_428),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_427),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_404),
.B(n_429),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_402),
.B(n_407),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_409),
.Y(n_452)
);

OA21x2_ASAP7_75t_L g453 ( 
.A1(n_421),
.A2(n_412),
.B(n_426),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_421),
.Y(n_454)
);

AO21x2_ASAP7_75t_L g455 ( 
.A1(n_408),
.A2(n_414),
.B(n_432),
.Y(n_455)
);

NOR2x1_ASAP7_75t_L g456 ( 
.A(n_432),
.B(n_414),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_432),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_414),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_422),
.B(n_358),
.Y(n_459)
);

AOI21x1_ASAP7_75t_L g460 ( 
.A1(n_430),
.A2(n_401),
.B(n_373),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_459),
.B(n_442),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_435),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_439),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_437),
.A2(n_459),
.B1(n_452),
.B2(n_444),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_446),
.B(n_450),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_447),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_438),
.B(n_450),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_458),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_457),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_454),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_456),
.Y(n_471)
);

CKINVDCx14_ASAP7_75t_R g472 ( 
.A(n_447),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_460),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_446),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_446),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_453),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_445),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_L g478 ( 
.A1(n_444),
.A2(n_450),
.B1(n_451),
.B2(n_441),
.Y(n_478)
);

OA21x2_ASAP7_75t_L g479 ( 
.A1(n_443),
.A2(n_441),
.B(n_455),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_455),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_453),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_441),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_468),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_474),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_467),
.B(n_436),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_465),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_463),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_478),
.B(n_449),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_463),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_461),
.B(n_451),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_474),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_462),
.A2(n_436),
.B1(n_449),
.B2(n_448),
.Y(n_492)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_475),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_466),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_472),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_467),
.B(n_440),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_461),
.B(n_440),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_468),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_469),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_465),
.B(n_440),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_469),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_473),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_462),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_477),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_470),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_465),
.B(n_475),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_465),
.B(n_440),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_470),
.B(n_464),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_482),
.B(n_480),
.Y(n_509)
);

INVxp67_ASAP7_75t_SL g510 ( 
.A(n_471),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_471),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_482),
.B(n_480),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_505),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_499),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_506),
.B(n_479),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_503),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_502),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_499),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_483),
.B(n_501),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_498),
.B(n_479),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_490),
.B(n_476),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_509),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_508),
.B(n_476),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_509),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_510),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_511),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_485),
.B(n_479),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_485),
.B(n_479),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_486),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_484),
.B(n_493),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_487),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_494),
.B(n_481),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_491),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_514),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_527),
.B(n_528),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_513),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_521),
.B(n_508),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_527),
.B(n_512),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_514),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_518),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_518),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_528),
.B(n_493),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_516),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_515),
.B(n_491),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_532),
.B(n_504),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_533),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_525),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_526),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_547),
.B(n_524),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_548),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_546),
.B(n_525),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_536),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_543),
.A2(n_488),
.B1(n_486),
.B2(n_497),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_535),
.B(n_515),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_535),
.B(n_524),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_534),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_539),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_539),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_L g559 ( 
.A1(n_545),
.A2(n_492),
.B(n_488),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_557),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_558),
.Y(n_561)
);

BUFx2_ASAP7_75t_SL g562 ( 
.A(n_549),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_553),
.A2(n_537),
.B1(n_523),
.B2(n_530),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_549),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_555),
.B(n_554),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_550),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_560),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_561),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_566),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_563),
.A2(n_559),
.B(n_553),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_563),
.A2(n_564),
.B1(n_552),
.B2(n_562),
.Y(n_571)
);

OAI22xp33_ASAP7_75t_L g572 ( 
.A1(n_566),
.A2(n_551),
.B1(n_552),
.B2(n_486),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_567),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_571),
.B(n_565),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_568),
.B(n_556),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_570),
.B(n_572),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_SL g577 ( 
.A1(n_569),
.A2(n_495),
.B(n_556),
.Y(n_577)
);

OAI32xp33_ASAP7_75t_L g578 ( 
.A1(n_571),
.A2(n_541),
.A3(n_540),
.B1(n_534),
.B2(n_542),
.Y(n_578)
);

AOI21xp33_ASAP7_75t_SL g579 ( 
.A1(n_576),
.A2(n_574),
.B(n_578),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_575),
.B(n_538),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_580),
.Y(n_581)
);

NOR3xp33_ASAP7_75t_L g582 ( 
.A(n_579),
.B(n_573),
.C(n_500),
.Y(n_582)
);

NAND4xp25_ASAP7_75t_L g583 ( 
.A(n_582),
.B(n_577),
.C(n_497),
.D(n_496),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_581),
.B(n_538),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_581),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_584),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_585),
.B(n_529),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_583),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_586),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_588),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_587),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_590),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_589),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_591),
.B(n_542),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_589),
.Y(n_595)
);

AOI21xp33_ASAP7_75t_L g596 ( 
.A1(n_595),
.A2(n_500),
.B(n_507),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_595),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_592),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_593),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_L g600 ( 
.A1(n_597),
.A2(n_594),
.B(n_496),
.Y(n_600)
);

AO21x2_ASAP7_75t_L g601 ( 
.A1(n_599),
.A2(n_519),
.B(n_507),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_598),
.B(n_519),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_596),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_597),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_604),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_603),
.A2(n_507),
.B1(n_529),
.B2(n_544),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_600),
.A2(n_529),
.B1(n_486),
.B2(n_531),
.Y(n_607)
);

AOI221xp5_ASAP7_75t_L g608 ( 
.A1(n_602),
.A2(n_522),
.B1(n_520),
.B2(n_487),
.C(n_489),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_605),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_606),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_SL g611 ( 
.A1(n_607),
.A2(n_601),
.B1(n_486),
.B2(n_522),
.Y(n_611)
);

OAI21x1_ASAP7_75t_L g612 ( 
.A1(n_608),
.A2(n_489),
.B(n_530),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_609),
.B(n_517),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_610),
.B(n_544),
.Y(n_614)
);

INVxp67_ASAP7_75t_L g615 ( 
.A(n_611),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_614),
.B(n_612),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_616),
.A2(n_615),
.B(n_613),
.Y(n_617)
);


endmodule