module fake_ibex_149_n_620 (n_85, n_84, n_64, n_3, n_73, n_65, n_103, n_95, n_55, n_63, n_98, n_29, n_106, n_2, n_76, n_8, n_67, n_9, n_38, n_37, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_48, n_57, n_59, n_28, n_39, n_5, n_62, n_71, n_93, n_13, n_61, n_14, n_0, n_94, n_12, n_42, n_77, n_88, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_22, n_4, n_33, n_30, n_6, n_100, n_72, n_26, n_34, n_97, n_102, n_15, n_24, n_52, n_99, n_105, n_1, n_25, n_36, n_104, n_41, n_45, n_18, n_89, n_83, n_32, n_53, n_107, n_50, n_11, n_92, n_101, n_96, n_68, n_79, n_81, n_35, n_31, n_56, n_23, n_91, n_54, n_19, n_620);

input n_85;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_103;
input n_95;
input n_55;
input n_63;
input n_98;
input n_29;
input n_106;
input n_2;
input n_76;
input n_8;
input n_67;
input n_9;
input n_38;
input n_37;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_48;
input n_57;
input n_59;
input n_28;
input n_39;
input n_5;
input n_62;
input n_71;
input n_93;
input n_13;
input n_61;
input n_14;
input n_0;
input n_94;
input n_12;
input n_42;
input n_77;
input n_88;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_22;
input n_4;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_34;
input n_97;
input n_102;
input n_15;
input n_24;
input n_52;
input n_99;
input n_105;
input n_1;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_50;
input n_11;
input n_92;
input n_101;
input n_96;
input n_68;
input n_79;
input n_81;
input n_35;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_620;

wire n_151;
wire n_599;
wire n_507;
wire n_540;
wire n_395;
wire n_171;
wire n_529;
wire n_389;
wire n_204;
wire n_274;
wire n_387;
wire n_130;
wire n_177;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_124;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_350;
wire n_601;
wire n_610;
wire n_165;
wire n_452;
wire n_255;
wire n_175;
wire n_586;
wire n_398;
wire n_125;
wire n_304;
wire n_191;
wire n_593;
wire n_153;
wire n_545;
wire n_583;
wire n_194;
wire n_249;
wire n_334;
wire n_312;
wire n_578;
wire n_478;
wire n_239;
wire n_134;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_216;
wire n_421;
wire n_475;
wire n_166;
wire n_163;
wire n_500;
wire n_542;
wire n_114;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_556;
wire n_189;
wire n_498;
wire n_317;
wire n_280;
wire n_340;
wire n_375;
wire n_187;
wire n_154;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_144;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_113;
wire n_561;
wire n_117;
wire n_417;
wire n_471;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_210;
wire n_348;
wire n_220;
wire n_481;
wire n_243;
wire n_287;
wire n_497;
wire n_228;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_426;
wire n_323;
wire n_469;
wire n_598;
wire n_143;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_333;
wire n_110;
wire n_306;
wire n_400;
wire n_550;
wire n_169;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_127;
wire n_121;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_120;
wire n_168;
wire n_526;
wire n_155;
wire n_315;
wire n_441;
wire n_604;
wire n_122;
wire n_523;
wire n_116;
wire n_614;
wire n_370;
wire n_431;
wire n_574;
wire n_289;
wire n_515;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_136;
wire n_261;
wire n_521;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_437;
wire n_602;
wire n_355;
wire n_474;
wire n_281;
wire n_594;
wire n_407;
wire n_490;
wire n_568;
wire n_448;
wire n_595;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_126;
wire n_585;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_141;
wire n_487;
wire n_222;
wire n_186;
wire n_524;
wire n_349;
wire n_454;
wire n_295;
wire n_331;
wire n_576;
wire n_230;
wire n_185;
wire n_388;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_167;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_618;
wire n_514;
wire n_139;
wire n_488;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_129;
wire n_613;
wire n_267;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_347;
wire n_473;
wire n_445;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_137;
wire n_338;
wire n_173;
wire n_477;
wire n_363;
wire n_402;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_401;
wire n_553;
wire n_554;
wire n_305;
wire n_307;
wire n_192;
wire n_140;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_365;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_516;
wire n_548;
wire n_567;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_562;
wire n_564;
wire n_506;
wire n_546;
wire n_199;
wire n_592;
wire n_495;
wire n_410;
wire n_308;
wire n_463;
wire n_411;
wire n_135;
wire n_520;
wire n_512;
wire n_615;
wire n_283;
wire n_397;
wire n_366;
wire n_111;
wire n_322;
wire n_227;
wire n_499;
wire n_115;
wire n_248;
wire n_451;
wire n_190;
wire n_138;
wire n_409;
wire n_582;
wire n_238;
wire n_214;
wire n_579;
wire n_332;
wire n_517;
wire n_211;
wire n_218;
wire n_314;
wire n_563;
wire n_132;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_535;
wire n_382;
wire n_502;
wire n_532;
wire n_405;
wire n_415;
wire n_597;
wire n_285;
wire n_288;
wire n_247;
wire n_320;
wire n_379;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_148;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_118;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_264;
wire n_198;
wire n_616;
wire n_217;
wire n_324;
wire n_391;
wire n_537;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_303;
wire n_362;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_501;
wire n_266;
wire n_294;
wire n_112;
wire n_485;
wire n_284;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_119;
wire n_361;
wire n_455;
wire n_419;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_311;
wire n_406;
wire n_606;
wire n_197;
wire n_528;
wire n_181;
wire n_131;
wire n_123;
wire n_260;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_572;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_252;
wire n_396;
wire n_149;
wire n_489;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_159;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_160;
wire n_184;
wire n_492;
wire n_232;
wire n_380;
wire n_559;
wire n_425;

INVxp67_ASAP7_75t_SL g110 ( 
.A(n_62),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_78),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_27),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_15),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_42),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_102),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_7),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_31),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_50),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_34),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_1),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_3),
.Y(n_128)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

INVxp33_ASAP7_75t_SL g130 ( 
.A(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_1),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

INVxp33_ASAP7_75t_SL g133 ( 
.A(n_4),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_91),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_73),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_20),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_49),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_17),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_39),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_32),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_55),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_11),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_43),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_22),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_63),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_23),
.Y(n_149)
);

INVxp67_ASAP7_75t_SL g150 ( 
.A(n_40),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_57),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_52),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_14),
.Y(n_153)
);

INVxp67_ASAP7_75t_SL g154 ( 
.A(n_24),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_16),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_37),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_67),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_54),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_76),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_58),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_3),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_88),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_28),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_101),
.B(n_66),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_103),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_21),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_48),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_6),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_30),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_97),
.Y(n_174)
);

INVxp33_ASAP7_75t_SL g175 ( 
.A(n_26),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_47),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

NOR2xp67_ASAP7_75t_L g178 ( 
.A(n_13),
.B(n_105),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_86),
.Y(n_179)
);

INVxp67_ASAP7_75t_SL g180 ( 
.A(n_71),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_0),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_69),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_11),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_77),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_100),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_29),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_80),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_84),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_5),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_144),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_122),
.B(n_0),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_129),
.B(n_2),
.Y(n_194)
);

OA21x2_ASAP7_75t_L g195 ( 
.A1(n_153),
.A2(n_44),
.B(n_96),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_117),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_129),
.B(n_2),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_171),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_145),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_127),
.B(n_4),
.Y(n_204)
);

CKINVDCx8_ASAP7_75t_R g205 ( 
.A(n_121),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_145),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_128),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_137),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_131),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_159),
.B(n_5),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_137),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_169),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_111),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_114),
.B(n_6),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_158),
.B(n_7),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_169),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_112),
.B(n_115),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_116),
.B(n_119),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_120),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_123),
.B(n_8),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_113),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_124),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_125),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_132),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_136),
.B(n_8),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_138),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_139),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_140),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_141),
.Y(n_233)
);

AND2x4_ASAP7_75t_L g234 ( 
.A(n_142),
.B(n_9),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_147),
.Y(n_235)
);

AND2x4_ASAP7_75t_L g236 ( 
.A(n_148),
.B(n_149),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_155),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_156),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_157),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_162),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_161),
.B(n_9),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_164),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_165),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_168),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_170),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_173),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_174),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_133),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_177),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_182),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_133),
.Y(n_251)
);

NAND2xp33_ASAP7_75t_SL g252 ( 
.A(n_113),
.B(n_118),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_184),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_118),
.A2(n_135),
.B1(n_143),
.B2(n_186),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_188),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_185),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_187),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_110),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_150),
.B(n_10),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_126),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_135),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_154),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_130),
.B(n_10),
.Y(n_263)
);

AND2x4_ASAP7_75t_L g264 ( 
.A(n_180),
.B(n_12),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_134),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_151),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_160),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_179),
.B(n_12),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_166),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_178),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_175),
.B(n_18),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_202),
.B(n_172),
.Y(n_272)
);

NAND2xp33_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_186),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_194),
.A2(n_172),
.B1(n_152),
.B2(n_143),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_L g275 ( 
.A1(n_248),
.A2(n_152),
.B1(n_19),
.B2(n_25),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_33),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_194),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_192),
.B(n_41),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_234),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_234),
.A2(n_45),
.B1(n_46),
.B2(n_51),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_56),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_265),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_197),
.B(n_59),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_211),
.A2(n_60),
.B1(n_64),
.B2(n_65),
.Y(n_284)
);

NOR2xp67_ASAP7_75t_L g285 ( 
.A(n_240),
.B(n_70),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_201),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_238),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_238),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_258),
.B(n_75),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_236),
.B(n_79),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_238),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_238),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_82),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_253),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_221),
.A2(n_83),
.B(n_87),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_208),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_236),
.B(n_89),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_236),
.B(n_94),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_210),
.Y(n_299)
);

AO22x2_ASAP7_75t_L g300 ( 
.A1(n_264),
.A2(n_204),
.B1(n_210),
.B2(n_262),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_266),
.B(n_262),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_212),
.A2(n_264),
.B1(n_244),
.B2(n_249),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_217),
.B(n_237),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_251),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_215),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_264),
.A2(n_193),
.B1(n_263),
.B2(n_241),
.Y(n_306)
);

INVx8_ASAP7_75t_L g307 ( 
.A(n_268),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_215),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_223),
.B(n_226),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_260),
.B(n_205),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_260),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_260),
.B(n_216),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_231),
.B(n_233),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_225),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_232),
.B(n_245),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_190),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_205),
.B(n_239),
.Y(n_317)
);

OR2x6_ASAP7_75t_L g318 ( 
.A(n_254),
.B(n_259),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_243),
.B(n_257),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_268),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_247),
.B(n_255),
.Y(n_321)
);

AO22x2_ASAP7_75t_L g322 ( 
.A1(n_270),
.A2(n_252),
.B1(n_214),
.B2(n_209),
.Y(n_322)
);

INVx5_ASAP7_75t_L g323 ( 
.A(n_246),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_261),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_246),
.B(n_255),
.Y(n_325)
);

NOR3xp33_ASAP7_75t_L g326 ( 
.A(n_252),
.B(n_263),
.C(n_229),
.Y(n_326)
);

XOR2x2_ASAP7_75t_L g327 ( 
.A(n_261),
.B(n_222),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g328 ( 
.A1(n_207),
.A2(n_242),
.B1(n_228),
.B2(n_256),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_218),
.A2(n_241),
.B1(n_219),
.B2(n_224),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_246),
.B(n_255),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_271),
.B(n_256),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_218),
.B(n_219),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_200),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_227),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_227),
.B(n_250),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_230),
.B(n_235),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_191),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_213),
.B(n_220),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_L g339 ( 
.A(n_203),
.B(n_206),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_196),
.B(n_198),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_213),
.B(n_196),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_199),
.A2(n_194),
.B1(n_210),
.B2(n_133),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_195),
.Y(n_343)
);

NAND2xp33_ASAP7_75t_SL g344 ( 
.A(n_195),
.B(n_194),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_195),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_248),
.A2(n_251),
.B1(n_194),
.B2(n_202),
.Y(n_346)
);

INVx8_ASAP7_75t_L g347 ( 
.A(n_202),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_202),
.B(n_269),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_202),
.B(n_269),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_202),
.B(n_269),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_202),
.B(n_269),
.Y(n_351)
);

NAND3xp33_ASAP7_75t_SL g352 ( 
.A(n_263),
.B(n_118),
.C(n_113),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_202),
.B(n_269),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_202),
.B(n_269),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_340),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_327),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_348),
.B(n_351),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_347),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_347),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_299),
.B(n_304),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_353),
.B(n_279),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_345),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_336),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_300),
.A2(n_346),
.B1(n_342),
.B2(n_306),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_316),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_325),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_347),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_354),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_312),
.B(n_329),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_329),
.B(n_332),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_316),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_334),
.Y(n_372)
);

A2O1A1Ixp33_ASAP7_75t_L g373 ( 
.A1(n_335),
.A2(n_344),
.B(n_306),
.C(n_309),
.Y(n_373)
);

BUFx2_ASAP7_75t_SL g374 ( 
.A(n_314),
.Y(n_374)
);

NAND2xp33_ASAP7_75t_L g375 ( 
.A(n_290),
.B(n_297),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_342),
.A2(n_302),
.B1(n_274),
.B2(n_318),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_307),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_337),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_303),
.B(n_315),
.Y(n_379)
);

AO22x1_ASAP7_75t_L g380 ( 
.A1(n_324),
.A2(n_272),
.B1(n_311),
.B2(n_273),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_330),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_L g382 ( 
.A1(n_322),
.A2(n_301),
.B1(n_319),
.B2(n_307),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_333),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_318),
.A2(n_322),
.B1(n_328),
.B2(n_313),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_341),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_339),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_323),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_307),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_323),
.Y(n_389)
);

BUFx12f_ASAP7_75t_L g390 ( 
.A(n_318),
.Y(n_390)
);

AO22x1_ASAP7_75t_L g391 ( 
.A1(n_275),
.A2(n_298),
.B1(n_352),
.B2(n_282),
.Y(n_391)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_317),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g393 ( 
.A(n_310),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_276),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_278),
.Y(n_395)
);

OR2x6_ASAP7_75t_L g396 ( 
.A(n_331),
.B(n_283),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_321),
.B(n_289),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_338),
.Y(n_398)
);

AND3x1_ASAP7_75t_SL g399 ( 
.A(n_287),
.B(n_294),
.C(n_292),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_285),
.B(n_343),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_285),
.B(n_281),
.Y(n_401)
);

CKINVDCx6p67_ASAP7_75t_R g402 ( 
.A(n_288),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_280),
.B(n_293),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_R g404 ( 
.A(n_277),
.B(n_284),
.Y(n_404)
);

BUFx4_ASAP7_75t_SL g405 ( 
.A(n_291),
.Y(n_405)
);

INVx4_ASAP7_75t_L g406 ( 
.A(n_296),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_305),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_295),
.B(n_308),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_286),
.B(n_320),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_348),
.B(n_269),
.Y(n_410)
);

BUFx4f_ASAP7_75t_L g411 ( 
.A(n_347),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_L g412 ( 
.A1(n_326),
.A2(n_300),
.B1(n_286),
.B2(n_234),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_347),
.Y(n_413)
);

OR2x6_ASAP7_75t_L g414 ( 
.A(n_307),
.B(n_347),
.Y(n_414)
);

OAI21x1_ASAP7_75t_L g415 ( 
.A1(n_343),
.A2(n_276),
.B(n_290),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_L g416 ( 
.A1(n_326),
.A2(n_300),
.B1(n_286),
.B2(n_234),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_327),
.Y(n_417)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_347),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_340),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_349),
.B(n_350),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_363),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_385),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_398),
.Y(n_423)
);

BUFx8_ASAP7_75t_SL g424 ( 
.A(n_390),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_367),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_375),
.A2(n_403),
.B(n_401),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_374),
.Y(n_427)
);

BUFx8_ASAP7_75t_L g428 ( 
.A(n_359),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_355),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_401),
.A2(n_400),
.B(n_397),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_379),
.B(n_357),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_357),
.Y(n_432)
);

OR2x6_ASAP7_75t_SL g433 ( 
.A(n_376),
.B(n_356),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_414),
.B(n_379),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_369),
.B(n_418),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_358),
.Y(n_436)
);

INVx2_ASAP7_75t_SL g437 ( 
.A(n_411),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_419),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_414),
.B(n_358),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_366),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_410),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_413),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_377),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_405),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_394),
.A2(n_361),
.B(n_415),
.Y(n_445)
);

INVx3_ASAP7_75t_SL g446 ( 
.A(n_414),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_378),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_360),
.B(n_376),
.Y(n_448)
);

NOR2xp67_ASAP7_75t_L g449 ( 
.A(n_364),
.B(n_392),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_383),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_388),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_365),
.Y(n_452)
);

INVx5_ASAP7_75t_L g453 ( 
.A(n_362),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_370),
.A2(n_369),
.B1(n_412),
.B2(n_416),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_373),
.A2(n_382),
.B1(n_384),
.B2(n_395),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_362),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_409),
.B(n_420),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_371),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_368),
.B(n_380),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g460 ( 
.A1(n_384),
.A2(n_404),
.B1(n_393),
.B2(n_386),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_417),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_372),
.B(n_381),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_391),
.B(n_396),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_389),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_396),
.B(n_389),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_402),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_387),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_408),
.B(n_406),
.Y(n_468)
);

OR2x6_ASAP7_75t_L g469 ( 
.A(n_406),
.B(n_399),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_407),
.A2(n_375),
.B(n_344),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_379),
.B(n_357),
.Y(n_471)
);

INVx3_ASAP7_75t_SL g472 ( 
.A(n_414),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_369),
.B(n_304),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_379),
.B(n_357),
.Y(n_474)
);

A2O1A1Ixp33_ASAP7_75t_L g475 ( 
.A1(n_370),
.A2(n_373),
.B(n_379),
.C(n_363),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_431),
.B(n_471),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_448),
.A2(n_454),
.B1(n_473),
.B2(n_441),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_474),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_432),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_429),
.B(n_438),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_427),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_434),
.B(n_421),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_422),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_422),
.A2(n_423),
.B1(n_475),
.B2(n_440),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_453),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_436),
.B(n_433),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_466),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_428),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_457),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_428),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_435),
.B(n_449),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_442),
.B(n_443),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_455),
.A2(n_460),
.B1(n_459),
.B2(n_463),
.Y(n_493)
);

AO31x2_ASAP7_75t_L g494 ( 
.A1(n_445),
.A2(n_426),
.A3(n_470),
.B(n_430),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_456),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_452),
.Y(n_496)
);

INVx6_ASAP7_75t_SL g497 ( 
.A(n_469),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_451),
.Y(n_498)
);

OR2x6_ASAP7_75t_L g499 ( 
.A(n_439),
.B(n_437),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_468),
.A2(n_469),
.B1(n_453),
.B2(n_439),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_465),
.B(n_464),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_447),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_467),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_462),
.Y(n_504)
);

BUFx4f_ASAP7_75t_SL g505 ( 
.A(n_446),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_472),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_444),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_425),
.B(n_458),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_461),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_L g510 ( 
.A1(n_450),
.A2(n_370),
.B1(n_448),
.B2(n_454),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_424),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_431),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_431),
.B(n_471),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_431),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_431),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_431),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_431),
.B(n_471),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_431),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_513),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_478),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_478),
.Y(n_521)
);

OR2x2_ASAP7_75t_L g522 ( 
.A(n_476),
.B(n_514),
.Y(n_522)
);

NOR2x1_ASAP7_75t_SL g523 ( 
.A(n_518),
.B(n_512),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_517),
.B(n_512),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_517),
.B(n_515),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_515),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_518),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_516),
.B(n_514),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_483),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_483),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_482),
.B(n_489),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_477),
.A2(n_493),
.B1(n_510),
.B2(n_484),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_492),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_477),
.B(n_510),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_494),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_496),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_479),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_493),
.B(n_480),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_505),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_495),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_488),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_530),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_522),
.B(n_486),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_SL g544 ( 
.A1(n_532),
.A2(n_500),
.B1(n_505),
.B2(n_490),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_522),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_524),
.B(n_491),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_524),
.B(n_485),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_528),
.Y(n_548)
);

OR2x6_ASAP7_75t_L g549 ( 
.A(n_519),
.B(n_495),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_528),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_534),
.A2(n_497),
.B1(n_504),
.B2(n_509),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_537),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_519),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_536),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_531),
.B(n_501),
.Y(n_555)
);

OR2x2_ASAP7_75t_SL g556 ( 
.A(n_520),
.B(n_526),
.Y(n_556)
);

INVx5_ASAP7_75t_L g557 ( 
.A(n_540),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_536),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_SL g559 ( 
.A(n_539),
.B(n_488),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_534),
.A2(n_497),
.B1(n_499),
.B2(n_498),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_525),
.B(n_485),
.Y(n_561)
);

NAND3xp33_ASAP7_75t_L g562 ( 
.A(n_535),
.B(n_503),
.C(n_502),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_542),
.A2(n_523),
.B(n_529),
.Y(n_563)
);

O2A1O1Ixp33_ASAP7_75t_SL g564 ( 
.A1(n_562),
.A2(n_520),
.B(n_521),
.C(n_526),
.Y(n_564)
);

OR2x6_ASAP7_75t_L g565 ( 
.A(n_553),
.B(n_539),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_554),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_545),
.B(n_533),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_555),
.B(n_531),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_558),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_548),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_546),
.B(n_521),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_542),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_550),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_546),
.B(n_527),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_552),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_543),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_572),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_571),
.B(n_561),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_575),
.Y(n_579)
);

CKINVDCx16_ASAP7_75t_R g580 ( 
.A(n_565),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_566),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_567),
.B(n_556),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_576),
.B(n_544),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_574),
.B(n_568),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_568),
.B(n_551),
.Y(n_585)
);

NOR2x1_ASAP7_75t_L g586 ( 
.A(n_565),
.B(n_511),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_578),
.B(n_569),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_584),
.B(n_570),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_580),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_583),
.B(n_573),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_579),
.B(n_563),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_581),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_582),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_583),
.B(n_563),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_577),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_SL g596 ( 
.A1(n_594),
.A2(n_586),
.B(n_585),
.Y(n_596)
);

NAND4xp25_ASAP7_75t_L g597 ( 
.A(n_590),
.B(n_585),
.C(n_560),
.D(n_559),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_592),
.Y(n_598)
);

NAND4xp25_ASAP7_75t_L g599 ( 
.A(n_590),
.B(n_481),
.C(n_538),
.D(n_508),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_593),
.B(n_535),
.Y(n_600)
);

NAND3xp33_ASAP7_75t_SL g601 ( 
.A(n_589),
.B(n_511),
.C(n_487),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_SL g602 ( 
.A(n_587),
.B(n_487),
.Y(n_602)
);

NAND4xp75_ASAP7_75t_L g603 ( 
.A(n_591),
.B(n_538),
.C(n_561),
.D(n_547),
.Y(n_603)
);

AOI221xp5_ASAP7_75t_L g604 ( 
.A1(n_596),
.A2(n_588),
.B1(n_595),
.B2(n_541),
.C(n_564),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_598),
.B(n_595),
.Y(n_605)
);

NOR2x1_ASAP7_75t_L g606 ( 
.A(n_601),
.B(n_565),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_SL g607 ( 
.A1(n_602),
.A2(n_553),
.B(n_523),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_599),
.A2(n_506),
.B(n_497),
.Y(n_608)
);

OAI22xp33_ASAP7_75t_L g609 ( 
.A1(n_597),
.A2(n_553),
.B1(n_549),
.B2(n_557),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_600),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_605),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_610),
.Y(n_612)
);

NOR2x1_ASAP7_75t_L g613 ( 
.A(n_606),
.B(n_603),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_611),
.B(n_604),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_612),
.B(n_609),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_614),
.B(n_613),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_616),
.Y(n_617)
);

NOR2x1_ASAP7_75t_SL g618 ( 
.A(n_617),
.B(n_608),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_618),
.Y(n_619)
);

AOI221xp5_ASAP7_75t_L g620 ( 
.A1(n_619),
.A2(n_615),
.B1(n_507),
.B2(n_506),
.C(n_607),
.Y(n_620)
);


endmodule