module fake_jpeg_522_n_687 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_687);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_687;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_15),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_7),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_59),
.Y(n_144)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_9),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_61),
.B(n_64),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g149 ( 
.A(n_62),
.Y(n_149)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_63),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_9),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_65),
.B(n_76),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_66),
.Y(n_141)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_68),
.Y(n_156)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_70),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_71),
.Y(n_159)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_73),
.Y(n_175)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_40),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_75),
.B(n_80),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_34),
.B(n_9),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_77),
.Y(n_184)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_78),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_79),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_40),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_40),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_81),
.B(n_86),
.Y(n_146)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_83),
.Y(n_208)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_84),
.Y(n_188)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_85),
.Y(n_195)
);

NOR2xp67_ASAP7_75t_L g86 ( 
.A(n_23),
.B(n_9),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_87),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_42),
.B(n_43),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_88),
.B(n_121),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_89),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_91),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_92),
.Y(n_225)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_94),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_95),
.Y(n_215)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_96),
.Y(n_161)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_97),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_50),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_98),
.B(n_105),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_100),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_22),
.B(n_26),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_101),
.B(n_119),
.Y(n_166)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_102),
.Y(n_183)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_103),
.Y(n_211)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_104),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_50),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_106),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_107),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_30),
.Y(n_108)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_108),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_38),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_50),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_110),
.B(n_116),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_111),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_112),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_30),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

INVx4_ASAP7_75t_SL g114 ( 
.A(n_47),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_30),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g212 ( 
.A(n_115),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_31),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_117),
.B(n_124),
.Y(n_173)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_118),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_22),
.B(n_18),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_23),
.Y(n_120)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_120),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_19),
.B(n_8),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_38),
.Y(n_122)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_122),
.Y(n_222)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_23),
.Y(n_123)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_41),
.Y(n_124)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_47),
.Y(n_125)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_31),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_126),
.B(n_127),
.Y(n_187)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_41),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_128),
.Y(n_199)
);

AND2x6_ASAP7_75t_L g129 ( 
.A(n_47),
.B(n_10),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_129),
.B(n_130),
.Y(n_189)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_61),
.B(n_37),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_132),
.B(n_193),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_114),
.A2(n_62),
.B1(n_38),
.B2(n_47),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g249 ( 
.A1(n_135),
.A2(n_142),
.B1(n_221),
.B2(n_197),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_72),
.B(n_58),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_139),
.B(n_182),
.Y(n_233)
);

BUFx24_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

BUFx4f_ASAP7_75t_SL g279 ( 
.A(n_140),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_62),
.A2(n_27),
.B1(n_54),
.B2(n_45),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_67),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_145),
.B(n_176),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_31),
.B1(n_54),
.B2(n_45),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_151),
.A2(n_197),
.B1(n_35),
.B2(n_37),
.Y(n_236)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

INVx4_ASAP7_75t_SL g253 ( 
.A(n_160),
.Y(n_253)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_68),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_165),
.Y(n_288)
);

BUFx12_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g260 ( 
.A(n_168),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_91),
.Y(n_174)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_174),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_78),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_70),
.Y(n_177)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_177),
.Y(n_235)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_118),
.Y(n_178)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_178),
.Y(n_244)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_100),
.Y(n_181)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_181),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_93),
.B(n_26),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_107),
.B(n_128),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_210),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_66),
.Y(n_193)
);

BUFx12_ASAP7_75t_L g196 ( 
.A(n_92),
.Y(n_196)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_196),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_71),
.A2(n_27),
.B1(n_54),
.B2(n_45),
.Y(n_197)
);

BUFx24_ASAP7_75t_L g198 ( 
.A(n_107),
.Y(n_198)
);

INVx11_ASAP7_75t_L g275 ( 
.A(n_198),
.Y(n_275)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_120),
.Y(n_202)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_202),
.Y(n_230)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_125),
.Y(n_203)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_96),
.Y(n_205)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_205),
.Y(n_294)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_97),
.Y(n_206)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_206),
.Y(n_303)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_123),
.Y(n_207)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_207),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_111),
.B(n_24),
.Y(n_210)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_73),
.Y(n_214)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_214),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_79),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_216),
.B(n_223),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_111),
.B(n_24),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_149),
.Y(n_234)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_83),
.Y(n_218)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_218),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_109),
.B(n_27),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_220),
.B(n_112),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_104),
.A2(n_27),
.B1(n_54),
.B2(n_45),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_87),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_182),
.A2(n_122),
.B1(n_44),
.B2(n_57),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_227),
.A2(n_249),
.B1(n_267),
.B2(n_283),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_189),
.A2(n_90),
.B1(n_115),
.B2(n_113),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_228),
.A2(n_236),
.B1(n_300),
.B2(n_306),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_187),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_229),
.B(n_238),
.Y(n_365)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_141),
.Y(n_232)
);

INVx5_ASAP7_75t_L g335 ( 
.A(n_232),
.Y(n_335)
);

OAI21xp33_ASAP7_75t_L g360 ( 
.A1(n_234),
.A2(n_258),
.B(n_272),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_141),
.Y(n_237)
);

INVx5_ASAP7_75t_L g349 ( 
.A(n_237),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_156),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_138),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_239),
.B(n_241),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_156),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_173),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_242),
.B(n_264),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_159),
.Y(n_245)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_245),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_159),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_246),
.Y(n_318)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_180),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_248),
.Y(n_333)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_175),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_250),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_149),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_251),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_146),
.A2(n_19),
.B1(n_56),
.B2(n_46),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_252),
.A2(n_262),
.B1(n_289),
.B2(n_302),
.Y(n_350)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_200),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_254),
.Y(n_312)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_194),
.Y(n_256)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_256),
.Y(n_332)
);

AND2x2_ASAP7_75t_SL g257 ( 
.A(n_139),
.B(n_128),
.Y(n_257)
);

XNOR2x1_ASAP7_75t_SL g352 ( 
.A(n_257),
.B(n_273),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_166),
.B(n_28),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_175),
.Y(n_259)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_259),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_144),
.A2(n_28),
.B1(n_33),
.B2(n_36),
.Y(n_262)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_204),
.Y(n_263)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_263),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_140),
.Y(n_264)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_194),
.Y(n_265)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_265),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_134),
.A2(n_37),
.B1(n_44),
.B2(n_57),
.Y(n_267)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_225),
.Y(n_268)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_268),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_191),
.B(n_112),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_269),
.B(n_280),
.Y(n_328)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_225),
.Y(n_270)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_270),
.Y(n_310)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_157),
.Y(n_271)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_271),
.Y(n_311)
);

AND2x2_ASAP7_75t_SL g273 ( 
.A(n_171),
.B(n_35),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_158),
.Y(n_274)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_274),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_204),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_276),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_190),
.Y(n_277)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_277),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_188),
.B(n_108),
.C(n_99),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_278),
.B(n_304),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_155),
.Y(n_280)
);

NAND2x1p5_ASAP7_75t_L g281 ( 
.A(n_184),
.B(n_35),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_281),
.A2(n_167),
.B(n_199),
.Y(n_317)
);

INVx8_ASAP7_75t_L g282 ( 
.A(n_180),
.Y(n_282)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_282),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_170),
.A2(n_44),
.B1(n_57),
.B2(n_31),
.Y(n_283)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_158),
.Y(n_286)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_286),
.Y(n_344)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_195),
.Y(n_287)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_287),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_211),
.A2(n_56),
.B1(n_33),
.B2(n_46),
.Y(n_289)
);

AOI21xp33_ASAP7_75t_L g290 ( 
.A1(n_136),
.A2(n_32),
.B(n_36),
.Y(n_290)
);

AOI32xp33_ASAP7_75t_L g358 ( 
.A1(n_290),
.A2(n_168),
.A3(n_196),
.B1(n_140),
.B2(n_198),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_164),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_291),
.B(n_292),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_132),
.B(n_95),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_220),
.A2(n_94),
.B1(n_89),
.B2(n_32),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_293),
.A2(n_167),
.B1(n_199),
.B2(n_180),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_133),
.B(n_11),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_295),
.B(n_297),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_174),
.Y(n_297)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_208),
.Y(n_298)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_298),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_143),
.B(n_11),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_299),
.B(n_301),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_142),
.A2(n_32),
.B1(n_55),
.B2(n_2),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_153),
.B(n_10),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_221),
.A2(n_10),
.B1(n_17),
.B2(n_16),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_183),
.B(n_7),
.C(n_16),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_147),
.B(n_5),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_305),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_135),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_306)
);

OAI32xp33_ASAP7_75t_L g308 ( 
.A1(n_255),
.A2(n_179),
.A3(n_161),
.B1(n_154),
.B2(n_201),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_308),
.B(n_361),
.Y(n_400)
);

OAI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_233),
.A2(n_222),
.B1(n_150),
.B2(n_163),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_313),
.A2(n_346),
.B1(n_265),
.B2(n_279),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_281),
.B(n_148),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_316),
.B(n_325),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_317),
.A2(n_196),
.B(n_296),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_247),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_320),
.B(n_358),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_281),
.B(n_148),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_233),
.A2(n_185),
.B1(n_186),
.B2(n_137),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_326),
.A2(n_356),
.B1(n_339),
.B2(n_346),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_228),
.A2(n_185),
.B1(n_208),
.B2(n_209),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_327),
.A2(n_339),
.B1(n_364),
.B2(n_279),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_330),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_226),
.B(n_131),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_334),
.B(n_272),
.C(n_304),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_273),
.B(n_172),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_337),
.B(n_338),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_273),
.B(n_172),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_300),
.A2(n_209),
.B1(n_213),
.B2(n_152),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_305),
.B(n_222),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_345),
.B(n_353),
.Y(n_384)
);

OAI22x1_ASAP7_75t_L g346 ( 
.A1(n_249),
.A2(n_224),
.B1(n_162),
.B2(n_212),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_257),
.B(n_186),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_267),
.A2(n_137),
.B1(n_215),
.B2(n_213),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_257),
.B(n_215),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_359),
.B(n_362),
.Y(n_397)
);

OA22x2_ASAP7_75t_L g361 ( 
.A1(n_227),
.A2(n_219),
.B1(n_163),
.B2(n_162),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_278),
.B(n_212),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_235),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_363),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_266),
.A2(n_219),
.B1(n_169),
.B2(n_152),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_294),
.Y(n_366)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_366),
.Y(n_390)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_294),
.Y(n_367)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_367),
.Y(n_401)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_303),
.Y(n_368)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_368),
.Y(n_403)
);

OAI22xp33_ASAP7_75t_SL g435 ( 
.A1(n_370),
.A2(n_394),
.B1(n_230),
.B2(n_331),
.Y(n_435)
);

INVx13_ASAP7_75t_L g371 ( 
.A(n_355),
.Y(n_371)
);

CKINVDCx14_ASAP7_75t_R g446 ( 
.A(n_371),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_322),
.A2(n_249),
.B1(n_293),
.B2(n_283),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_372),
.A2(n_386),
.B1(n_398),
.B2(n_404),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_326),
.A2(n_306),
.B1(n_288),
.B2(n_275),
.Y(n_373)
);

OAI21xp33_ASAP7_75t_SL g419 ( 
.A1(n_373),
.A2(n_382),
.B(n_361),
.Y(n_419)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_307),
.Y(n_374)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_374),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g375 ( 
.A(n_315),
.Y(n_375)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_375),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_377),
.B(n_399),
.Y(n_427)
);

OAI32xp33_ASAP7_75t_L g378 ( 
.A1(n_316),
.A2(n_303),
.A3(n_261),
.B1(n_284),
.B2(n_285),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_378),
.B(n_367),
.Y(n_433)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_307),
.Y(n_381)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_381),
.Y(n_440)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_311),
.A2(n_288),
.B1(n_275),
.B2(n_256),
.Y(n_382)
);

AND2x6_ASAP7_75t_L g383 ( 
.A(n_334),
.B(n_279),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_383),
.B(n_395),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_348),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g423 ( 
.A1(n_385),
.A2(n_388),
.B1(n_391),
.B2(n_315),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_322),
.A2(n_314),
.B1(n_325),
.B2(n_362),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_324),
.B(n_240),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_387),
.Y(n_431)
);

INVx13_ASAP7_75t_L g388 ( 
.A(n_355),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_328),
.B(n_251),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_389),
.Y(n_450)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_335),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_392),
.Y(n_451)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_335),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_393),
.B(n_406),
.Y(n_424)
);

AND2x6_ASAP7_75t_L g395 ( 
.A(n_352),
.B(n_198),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_327),
.A2(n_169),
.B1(n_298),
.B2(n_232),
.Y(n_398)
);

AND2x2_ASAP7_75t_SL g399 ( 
.A(n_352),
.B(n_286),
.Y(n_399)
);

NAND2x1_ASAP7_75t_L g402 ( 
.A(n_317),
.B(n_274),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_402),
.A2(n_412),
.B(n_361),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_353),
.A2(n_250),
.B1(n_263),
.B2(n_259),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_359),
.A2(n_237),
.B1(n_245),
.B2(n_276),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_405),
.A2(n_415),
.B1(n_360),
.B2(n_351),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_336),
.Y(n_406)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_315),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_407),
.B(n_408),
.Y(n_436)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_351),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_366),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_409),
.B(n_347),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_319),
.B(n_244),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_410),
.B(n_414),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_311),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_411),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_337),
.A2(n_270),
.B(n_268),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_341),
.B(n_296),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_413),
.B(n_347),
.C(n_365),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_343),
.B(n_231),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_341),
.A2(n_338),
.B1(n_350),
.B2(n_342),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_321),
.A2(n_231),
.B1(n_271),
.B2(n_246),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_416),
.A2(n_349),
.B1(n_318),
.B2(n_253),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_417),
.A2(n_344),
.B(n_323),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_418),
.A2(n_434),
.B(n_447),
.Y(n_463)
);

BUFx5_ASAP7_75t_L g462 ( 
.A(n_419),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_369),
.A2(n_329),
.B1(n_345),
.B2(n_308),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_421),
.A2(n_435),
.B1(n_455),
.B2(n_391),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_423),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_425),
.B(n_428),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_417),
.A2(n_361),
.B(n_336),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_429),
.A2(n_402),
.B(n_400),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_430),
.B(n_442),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_369),
.B(n_368),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_432),
.B(n_449),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_433),
.B(n_438),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_SL g434 ( 
.A1(n_379),
.A2(n_331),
.B1(n_309),
.B2(n_332),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_415),
.B(n_312),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_386),
.A2(n_354),
.B1(n_348),
.B2(n_340),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_441),
.A2(n_370),
.B1(n_416),
.B2(n_375),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_413),
.B(n_357),
.Y(n_442)
);

AO22x1_ASAP7_75t_L g443 ( 
.A1(n_400),
.A2(n_323),
.B1(n_344),
.B2(n_310),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_443),
.B(n_445),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_377),
.B(n_310),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_453),
.C(n_399),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_397),
.B(n_309),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_397),
.B(n_354),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_448),
.B(n_458),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_384),
.B(n_376),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_384),
.B(n_376),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_452),
.B(n_456),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_399),
.B(n_363),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_400),
.A2(n_340),
.B1(n_349),
.B2(n_318),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_414),
.B(n_332),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_457),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_402),
.B(n_403),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_460),
.B(n_404),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_461),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_464),
.A2(n_455),
.B1(n_443),
.B2(n_441),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_465),
.A2(n_475),
.B1(n_385),
.B2(n_393),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_445),
.B(n_380),
.Y(n_466)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_466),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_458),
.B(n_394),
.Y(n_467)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_467),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_454),
.B(n_406),
.Y(n_468)
);

NAND3xp33_ASAP7_75t_L g522 ( 
.A(n_468),
.B(n_479),
.C(n_484),
.Y(n_522)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_425),
.Y(n_469)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_469),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_427),
.B(n_383),
.C(n_395),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_471),
.B(n_488),
.C(n_444),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_446),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_472),
.B(n_483),
.Y(n_502)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_448),
.Y(n_473)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_473),
.Y(n_497)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_422),
.Y(n_474)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_474),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_426),
.A2(n_372),
.B1(n_412),
.B2(n_379),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_451),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_476),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_418),
.A2(n_396),
.B(n_390),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_478),
.A2(n_480),
.B(n_496),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_454),
.B(n_409),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_429),
.A2(n_396),
.B(n_403),
.Y(n_480)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_422),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_450),
.B(n_390),
.Y(n_484)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_440),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_486),
.B(n_492),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_427),
.B(n_401),
.Y(n_488)
);

CKINVDCx16_ASAP7_75t_R g489 ( 
.A(n_424),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_489),
.B(n_424),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_431),
.B(n_401),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_490),
.B(n_491),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_456),
.B(n_408),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_446),
.Y(n_492)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_440),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_495),
.B(n_437),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_447),
.A2(n_385),
.B(n_371),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_499),
.B(n_529),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_488),
.B(n_442),
.C(n_453),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_500),
.B(n_501),
.C(n_506),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_488),
.B(n_430),
.C(n_438),
.Y(n_501)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_503),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_494),
.B(n_449),
.C(n_452),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_490),
.B(n_421),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g548 ( 
.A(n_508),
.B(n_512),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_494),
.B(n_432),
.C(n_420),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_510),
.B(n_513),
.C(n_460),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_481),
.A2(n_426),
.B1(n_420),
.B2(n_433),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_511),
.A2(n_518),
.B1(n_528),
.B2(n_477),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_479),
.B(n_487),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_494),
.B(n_428),
.C(n_439),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_487),
.B(n_439),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g563 ( 
.A(n_514),
.B(n_525),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_516),
.A2(n_527),
.B1(n_533),
.B2(n_459),
.Y(n_545)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_517),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_481),
.A2(n_443),
.B1(n_436),
.B2(n_437),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_484),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_519),
.B(n_531),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_466),
.B(n_392),
.Y(n_521)
);

CKINVDCx14_ASAP7_75t_R g541 ( 
.A(n_521),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_476),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_523),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_470),
.B(n_451),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_475),
.A2(n_398),
.B1(n_457),
.B2(n_405),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_465),
.A2(n_436),
.B1(n_451),
.B2(n_375),
.Y(n_528)
);

OA22x2_ASAP7_75t_L g530 ( 
.A1(n_459),
.A2(n_378),
.B1(n_407),
.B2(n_374),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_530),
.B(n_464),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_470),
.B(n_468),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_460),
.B(n_381),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_532),
.B(n_496),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_537),
.A2(n_528),
.B1(n_505),
.B2(n_526),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_523),
.Y(n_538)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_538),
.Y(n_570)
);

NOR3xp33_ASAP7_75t_SL g539 ( 
.A(n_520),
.B(n_471),
.C(n_467),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_539),
.B(n_549),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_540),
.B(n_547),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_506),
.B(n_489),
.Y(n_543)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_543),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_516),
.A2(n_485),
.B1(n_477),
.B2(n_461),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_544),
.A2(n_545),
.B1(n_550),
.B2(n_551),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_L g546 ( 
.A1(n_498),
.A2(n_478),
.B(n_480),
.Y(n_546)
);

INVxp33_ASAP7_75t_L g584 ( 
.A(n_546),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_532),
.B(n_501),
.Y(n_547)
);

NOR3xp33_ASAP7_75t_SL g549 ( 
.A(n_515),
.B(n_471),
.C(n_467),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_509),
.A2(n_485),
.B1(n_473),
.B2(n_493),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_509),
.A2(n_493),
.B1(n_469),
.B2(n_482),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_552),
.B(n_498),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_499),
.B(n_513),
.C(n_510),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_553),
.B(n_555),
.C(n_558),
.Y(n_571)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_502),
.Y(n_554)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_554),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_500),
.B(n_463),
.C(n_486),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_522),
.B(n_524),
.Y(n_557)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_557),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_529),
.B(n_463),
.C(n_495),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_559),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_511),
.B(n_491),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_560),
.B(n_518),
.Y(n_574)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_502),
.Y(n_561)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_561),
.Y(n_578)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_504),
.Y(n_562)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_562),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_527),
.A2(n_462),
.B1(n_492),
.B2(n_472),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_564),
.A2(n_566),
.B1(n_526),
.B2(n_507),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_515),
.A2(n_462),
.B1(n_483),
.B2(n_474),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_534),
.B(n_504),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_567),
.B(n_589),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_SL g602 ( 
.A(n_569),
.B(n_574),
.Y(n_602)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_565),
.Y(n_572)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_572),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_534),
.B(n_497),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_576),
.B(n_580),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_535),
.B(n_497),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_547),
.B(n_505),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_581),
.B(n_586),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_583),
.Y(n_608)
);

XNOR2x1_ASAP7_75t_SL g586 ( 
.A(n_552),
.B(n_462),
.Y(n_586)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_588),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_535),
.B(n_530),
.C(n_507),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_542),
.Y(n_590)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_590),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_563),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_591),
.A2(n_556),
.B1(n_548),
.B2(n_541),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_553),
.B(n_530),
.C(n_333),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_592),
.B(n_593),
.C(n_558),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g593 ( 
.A(n_540),
.B(n_555),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_575),
.B(n_536),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g630 ( 
.A(n_594),
.B(n_595),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g627 ( 
.A(n_596),
.B(n_333),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_SL g597 ( 
.A1(n_584),
.A2(n_546),
.B(n_559),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_SL g623 ( 
.A1(n_597),
.A2(n_603),
.B(n_612),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_568),
.B(n_576),
.C(n_593),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_598),
.B(n_600),
.Y(n_628)
);

XOR2x2_ASAP7_75t_L g599 ( 
.A(n_589),
.B(n_544),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_599),
.B(n_605),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_568),
.B(n_562),
.C(n_554),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_580),
.B(n_560),
.C(n_537),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_601),
.B(n_614),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_SL g603 ( 
.A1(n_584),
.A2(n_587),
.B(n_585),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_582),
.B(n_550),
.Y(n_605)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_570),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_611),
.B(n_613),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_SL g612 ( 
.A1(n_586),
.A2(n_549),
.B(n_539),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_578),
.B(n_566),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_571),
.B(n_551),
.C(n_564),
.Y(n_614)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_572),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_616),
.B(n_254),
.Y(n_631)
);

CKINVDCx16_ASAP7_75t_R g617 ( 
.A(n_594),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_617),
.B(n_618),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_598),
.B(n_571),
.C(n_592),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_603),
.B(n_577),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_619),
.B(n_621),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_610),
.B(n_573),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_596),
.B(n_581),
.C(n_574),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_622),
.B(n_624),
.C(n_601),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_614),
.B(n_569),
.C(n_579),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_600),
.B(n_565),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_SL g637 ( 
.A(n_625),
.B(n_627),
.Y(n_637)
);

XOR2xp5_ASAP7_75t_L g626 ( 
.A(n_599),
.B(n_530),
.Y(n_626)
);

XOR2xp5_ASAP7_75t_L g650 ( 
.A(n_626),
.B(n_212),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_631),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_608),
.A2(n_277),
.B1(n_248),
.B2(n_282),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_633),
.A2(n_606),
.B1(n_609),
.B2(n_613),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_606),
.B(n_243),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_634),
.B(n_616),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_SL g635 ( 
.A1(n_608),
.A2(n_388),
.B1(n_230),
.B2(n_243),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_SL g642 ( 
.A1(n_635),
.A2(n_609),
.B1(n_605),
.B2(n_253),
.Y(n_642)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_636),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_638),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_623),
.A2(n_612),
.B(n_597),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_639),
.B(n_641),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_632),
.B(n_611),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_642),
.A2(n_643),
.B1(n_648),
.B2(n_633),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g643 ( 
.A1(n_623),
.A2(n_607),
.B(n_604),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_644),
.B(n_650),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_618),
.B(n_615),
.C(n_602),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_646),
.B(n_622),
.C(n_627),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_620),
.A2(n_607),
.B(n_602),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_628),
.B(n_629),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_SL g653 ( 
.A(n_649),
.B(n_624),
.Y(n_653)
);

NAND2x1_ASAP7_75t_L g651 ( 
.A(n_620),
.B(n_260),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_651),
.B(n_635),
.Y(n_658)
);

OAI21x1_ASAP7_75t_L g664 ( 
.A1(n_653),
.A2(n_659),
.B(n_637),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_SL g654 ( 
.A1(n_645),
.A2(n_630),
.B(n_632),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_654),
.B(n_655),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_SL g669 ( 
.A1(n_658),
.A2(n_661),
.B1(n_650),
.B2(n_260),
.Y(n_669)
);

NOR2xp67_ASAP7_75t_L g659 ( 
.A(n_647),
.B(n_630),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g662 ( 
.A(n_644),
.B(n_626),
.C(n_260),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_662),
.B(n_648),
.Y(n_668)
);

BUFx24_ASAP7_75t_SL g663 ( 
.A(n_639),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_SL g666 ( 
.A(n_663),
.B(n_646),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_664),
.A2(n_5),
.B(n_15),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_666),
.B(n_670),
.Y(n_676)
);

AOI322xp5_ASAP7_75t_L g667 ( 
.A1(n_652),
.A2(n_641),
.A3(n_643),
.B1(n_636),
.B2(n_640),
.C1(n_642),
.C2(n_651),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_667),
.B(n_669),
.Y(n_674)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_668),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_660),
.A2(n_190),
.B1(n_11),
.B2(n_13),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_657),
.A2(n_656),
.B1(n_662),
.B2(n_655),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_SL g673 ( 
.A1(n_671),
.A2(n_672),
.B(n_4),
.Y(n_673)
);

AOI322xp5_ASAP7_75t_L g672 ( 
.A1(n_654),
.A2(n_5),
.A3(n_16),
.B1(n_15),
.B2(n_13),
.C1(n_4),
.C2(n_18),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_673),
.A2(n_675),
.B(n_677),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_665),
.A2(n_5),
.B(n_18),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_678),
.B(n_671),
.Y(n_679)
);

AOI31xp33_ASAP7_75t_L g683 ( 
.A1(n_679),
.A2(n_0),
.A3(n_1),
.B(n_2),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_674),
.Y(n_680)
);

AO21x2_ASAP7_75t_L g682 ( 
.A1(n_680),
.A2(n_676),
.B(n_669),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_682),
.B(n_683),
.Y(n_684)
);

XNOR2xp5_ASAP7_75t_L g685 ( 
.A(n_684),
.B(n_681),
.Y(n_685)
);

MAJIxp5_ASAP7_75t_L g686 ( 
.A(n_685),
.B(n_2),
.C(n_3),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_686),
.Y(n_687)
);


endmodule