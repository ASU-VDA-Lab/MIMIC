module fake_jpeg_23102_n_260 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_260);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_260;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_100;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx4f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx2_ASAP7_75t_SL g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_14),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_28),
.Y(n_49)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

CKINVDCx12_ASAP7_75t_R g41 ( 
.A(n_37),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_45),
.Y(n_79)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_18),
.B1(n_25),
.B2(n_16),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_49),
.B(n_17),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_50),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_17),
.B(n_22),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_27),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_30),
.Y(n_53)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_56),
.B(n_29),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_60),
.Y(n_92)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_66),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_25),
.B1(n_18),
.B2(n_26),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_52),
.B1(n_25),
.B2(n_46),
.Y(n_91)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_35),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_75),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_71),
.Y(n_100)
);

MAJx2_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_19),
.C(n_27),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_27),
.C(n_19),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_35),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_19),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_79),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_89),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_85),
.A2(n_88),
.B(n_33),
.Y(n_111)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_93),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_32),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_70),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_91),
.A2(n_95),
.B1(n_66),
.B2(n_60),
.Y(n_122)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_68),
.A2(n_33),
.B1(n_31),
.B2(n_44),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_98),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_68),
.A2(n_20),
.B(n_14),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_28),
.B(n_20),
.Y(n_105)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_43),
.C(n_42),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_102),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_35),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_34),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_76),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_74),
.Y(n_124)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_106),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_105),
.B(n_111),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_67),
.B1(n_96),
.B2(n_16),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_103),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_110),
.Y(n_136)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_120),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_16),
.B1(n_57),
.B2(n_72),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_114),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_31),
.B1(n_53),
.B2(n_76),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_116),
.A2(n_119),
.B1(n_91),
.B2(n_85),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_63),
.B1(n_74),
.B2(n_16),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_122),
.B1(n_90),
.B2(n_87),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_61),
.Y(n_118)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_88),
.A2(n_63),
.B1(n_78),
.B2(n_61),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_125),
.Y(n_132)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_101),
.B(n_24),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_97),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_105),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_88),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_133),
.Y(n_152)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_138),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_109),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_113),
.A2(n_82),
.B1(n_102),
.B2(n_90),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_140),
.A2(n_142),
.B1(n_144),
.B2(n_104),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_82),
.Y(n_141)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_100),
.B1(n_98),
.B2(n_72),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_34),
.B1(n_32),
.B2(n_58),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_34),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_148),
.Y(n_159)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_136),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_149),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g151 ( 
.A(n_130),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_153),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_136),
.Y(n_153)
);

AOI22x1_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_116),
.B1(n_111),
.B2(n_119),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_154),
.A2(n_138),
.B1(n_128),
.B2(n_133),
.Y(n_171)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_160),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_158),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_109),
.C(n_112),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_127),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_127),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_164),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_125),
.Y(n_162)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_167),
.Y(n_184)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_168),
.A2(n_148),
.B1(n_137),
.B2(n_135),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_109),
.C(n_110),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_145),
.Y(n_182)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_171),
.B(n_172),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_154),
.B(n_140),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_132),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_177),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_139),
.Y(n_176)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_131),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_179),
.A2(n_187),
.B(n_159),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_157),
.C(n_159),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_185),
.A2(n_144),
.B1(n_118),
.B2(n_165),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_130),
.B(n_135),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_154),
.A2(n_157),
.B1(n_168),
.B2(n_158),
.Y(n_189)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_108),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_24),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_29),
.C(n_21),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_183),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_193),
.B(n_194),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_65),
.C(n_123),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_203),
.C(n_204),
.Y(n_209)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_200),
.Y(n_207)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_201),
.A2(n_188),
.B1(n_179),
.B2(n_186),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_165),
.C(n_147),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_172),
.C(n_180),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_206),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_143),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_208),
.A2(n_14),
.B1(n_24),
.B2(n_3),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_197),
.A2(n_178),
.B1(n_190),
.B2(n_177),
.Y(n_210)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_175),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_213),
.C(n_218),
.Y(n_222)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_217),
.Y(n_230)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_22),
.C(n_21),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_24),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_219),
.B(n_1),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_58),
.C(n_32),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_202),
.C(n_20),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_215),
.A2(n_202),
.B1(n_195),
.B2(n_28),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_224),
.C(n_228),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_225),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_227),
.Y(n_236)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_214),
.A2(n_13),
.B1(n_12),
.B2(n_3),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_2),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_212),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_209),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_232),
.B(n_234),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_209),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_235),
.B(n_237),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_211),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_239),
.A2(n_2),
.B(n_4),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_2),
.C(n_3),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_240),
.B(n_6),
.Y(n_246)
);

AOI322xp5_ASAP7_75t_L g242 ( 
.A1(n_238),
.A2(n_230),
.A3(n_228),
.B1(n_224),
.B2(n_24),
.C1(n_8),
.C2(n_9),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_7),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_244),
.B(n_246),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_236),
.A2(n_6),
.B(n_7),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_239),
.B(n_9),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_24),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_23),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_250),
.Y(n_253)
);

OAI21x1_ASAP7_75t_L g255 ( 
.A1(n_251),
.A2(n_8),
.B(n_11),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_8),
.C(n_10),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_252),
.A2(n_243),
.B(n_11),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_254),
.A2(n_255),
.B(n_23),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_249),
.C(n_11),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_256),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_257),
.Y(n_259)
);

AO21x1_ASAP7_75t_L g260 ( 
.A1(n_259),
.A2(n_23),
.B(n_178),
.Y(n_260)
);


endmodule