module fake_jpeg_19700_n_327 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_37),
.Y(n_52)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_29),
.Y(n_48)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_17),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_49),
.B(n_18),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_29),
.B1(n_16),
.B2(n_26),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_51),
.B1(n_55),
.B2(n_35),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_29),
.B1(n_16),
.B2(n_26),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_16),
.B1(n_26),
.B2(n_31),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_37),
.B1(n_36),
.B2(n_38),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_56),
.A2(n_60),
.B1(n_37),
.B2(n_36),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_22),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_42),
.Y(n_70)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_18),
.B1(n_21),
.B2(n_32),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_58),
.A2(n_37),
.B1(n_36),
.B2(n_34),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_61),
.A2(n_66),
.B1(n_69),
.B2(n_72),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_63),
.B(n_68),
.Y(n_96)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_71),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_38),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_38),
.B1(n_35),
.B2(n_37),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_35),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_73),
.B(n_74),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_42),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_32),
.B1(n_21),
.B2(n_27),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_49),
.B(n_36),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_76),
.B(n_77),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_27),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_43),
.B1(n_40),
.B2(n_32),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_59),
.B1(n_53),
.B2(n_54),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_42),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_83),
.C(n_84),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_60),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_80),
.Y(n_115)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_82),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_42),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_51),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_56),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_90),
.A2(n_57),
.B1(n_40),
.B2(n_54),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_89),
.A2(n_57),
.B1(n_21),
.B2(n_46),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

AO22x2_ASAP7_75t_L g101 ( 
.A1(n_69),
.A2(n_79),
.B1(n_83),
.B2(n_73),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_79),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_25),
.C(n_43),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_114),
.C(n_116),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_59),
.B1(n_53),
.B2(n_43),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_103),
.A2(n_105),
.B1(n_82),
.B2(n_64),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_104),
.A2(n_107),
.B1(n_84),
.B2(n_44),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_71),
.A2(n_46),
.B1(n_54),
.B2(n_44),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_66),
.A2(n_54),
.B1(n_44),
.B2(n_42),
.Y(n_107)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_62),
.C(n_70),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_62),
.B(n_41),
.C(n_44),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

AOI21xp33_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_76),
.B(n_74),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_121),
.A2(n_101),
.B(n_109),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_115),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_123),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_68),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_112),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_124),
.B(n_131),
.Y(n_161)
);

AOI21x1_ASAP7_75t_L g181 ( 
.A1(n_125),
.A2(n_25),
.B(n_120),
.Y(n_181)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_129),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_83),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_130),
.Y(n_156)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_75),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_118),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_133),
.B(n_149),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_134),
.A2(n_141),
.B1(n_105),
.B2(n_109),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_24),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_143),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_140),
.B1(n_145),
.B2(n_147),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_119),
.C(n_92),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_142),
.C(n_116),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_95),
.A2(n_81),
.B1(n_90),
.B2(n_88),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_100),
.A2(n_111),
.B1(n_95),
.B2(n_92),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_91),
.C(n_86),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_98),
.B(n_91),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_100),
.A2(n_41),
.B1(n_30),
.B2(n_20),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_91),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_101),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_111),
.A2(n_41),
.B1(n_30),
.B2(n_20),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_106),
.A2(n_30),
.B1(n_20),
.B2(n_19),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_145),
.B1(n_104),
.B2(n_107),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_106),
.B(n_24),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_151),
.A2(n_23),
.B1(n_14),
.B2(n_13),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_152),
.B(n_153),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_128),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_154),
.B(n_166),
.Y(n_203)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_133),
.C(n_147),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_102),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_160),
.B(n_163),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_101),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_173),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_144),
.A2(n_101),
.B(n_110),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_165),
.A2(n_170),
.B(n_174),
.Y(n_207)
);

OAI31xp33_ASAP7_75t_L g167 ( 
.A1(n_125),
.A2(n_146),
.A3(n_122),
.B(n_127),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g213 ( 
.A1(n_167),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_213)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_103),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_179),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_130),
.A2(n_136),
.B(n_121),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_171),
.A2(n_180),
.B1(n_126),
.B2(n_1),
.Y(n_189)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_141),
.B(n_25),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_91),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_123),
.B(n_25),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_181),
.Y(n_204)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_124),
.Y(n_176)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_132),
.A2(n_94),
.B(n_19),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_177),
.A2(n_0),
.B(n_1),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_137),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_134),
.A2(n_99),
.B1(n_120),
.B2(n_31),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_99),
.Y(n_183)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_185),
.B(n_186),
.C(n_199),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_148),
.C(n_129),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_189),
.A2(n_197),
.B1(n_214),
.B2(n_156),
.Y(n_222)
);

OA21x2_ASAP7_75t_L g190 ( 
.A1(n_152),
.A2(n_25),
.B(n_28),
.Y(n_190)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_23),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_191),
.B(n_193),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_162),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_176),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_195),
.A2(n_153),
.B(n_210),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_31),
.C(n_28),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_31),
.C(n_28),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_2),
.C(n_3),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_23),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_165),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_209),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_157),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_208),
.A2(n_212),
.B1(n_151),
.B2(n_156),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_162),
.B(n_13),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_174),
.A2(n_169),
.B1(n_173),
.B2(n_166),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_174),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_167),
.A2(n_10),
.B(n_11),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_215),
.A2(n_220),
.B(n_239),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_198),
.B(n_164),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_221),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_195),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_222),
.Y(n_241)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_184),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_224),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_195),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_229),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_181),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_237),
.C(n_198),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_208),
.A2(n_178),
.B1(n_177),
.B2(n_182),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_228),
.A2(n_238),
.B1(n_227),
.B2(n_190),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_212),
.A2(n_172),
.B1(n_168),
.B2(n_175),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_0),
.Y(n_230)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_189),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_231)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_2),
.Y(n_233)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_233),
.Y(n_245)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_194),
.Y(n_235)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_2),
.Y(n_236)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_3),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_207),
.A2(n_8),
.B(n_5),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_217),
.A2(n_207),
.B1(n_185),
.B2(n_186),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_240),
.A2(n_246),
.B1(n_247),
.B2(n_225),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_226),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_217),
.A2(n_220),
.B1(n_215),
.B2(n_219),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_227),
.A2(n_233),
.B1(n_238),
.B2(n_236),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_196),
.C(n_199),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_252),
.C(n_254),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_205),
.C(n_202),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_204),
.C(n_200),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_216),
.B(n_201),
.Y(n_255)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_255),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_257),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_223),
.A2(n_190),
.B1(n_206),
.B2(n_187),
.Y(n_259)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_230),
.B(n_192),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_260),
.B(n_231),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_234),
.Y(n_261)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_256),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_263),
.Y(n_285)
);

BUFx12_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_268),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_244),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_241),
.A2(n_239),
.B(n_235),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_188),
.Y(n_269)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_245),
.A2(n_221),
.B1(n_229),
.B2(n_237),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_271),
.A2(n_276),
.B1(n_242),
.B2(n_247),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_250),
.B(n_234),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_272),
.B(n_273),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_250),
.B(n_204),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_274),
.B(n_277),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_251),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_249),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_266),
.A2(n_241),
.B(n_248),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_286),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_287),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_264),
.A2(n_243),
.B1(n_251),
.B2(n_242),
.Y(n_280)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_280),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_252),
.C(n_240),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_283),
.B(n_284),
.Y(n_295)
);

BUFx24_ASAP7_75t_SL g286 ( 
.A(n_275),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_254),
.Y(n_287)
);

MAJx2_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_258),
.C(n_253),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_265),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_263),
.B(n_258),
.C(n_253),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_292),
.B(n_269),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_289),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_298),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_279),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_297),
.C(n_299),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_271),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_262),
.C(n_268),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_249),
.C(n_265),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_288),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_269),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_303),
.A2(n_304),
.B(n_291),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_303),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_308),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_281),
.Y(n_306)
);

OAI21xp33_ASAP7_75t_L g316 ( 
.A1(n_306),
.A2(n_310),
.B(n_4),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_295),
.B(n_282),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_309),
.B(n_311),
.Y(n_315)
);

NOR2x1_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_243),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_300),
.B(n_4),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_313),
.B(n_4),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_310),
.A2(n_302),
.B1(n_297),
.B2(n_296),
.Y(n_314)
);

OAI321xp33_ASAP7_75t_L g320 ( 
.A1(n_314),
.A2(n_316),
.A3(n_317),
.B1(n_305),
.B2(n_7),
.C(n_8),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_5),
.Y(n_318)
);

AO21x2_ASAP7_75t_L g321 ( 
.A1(n_318),
.A2(n_6),
.B(n_7),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_320),
.A2(n_321),
.B(n_322),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_312),
.B(n_6),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_315),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_6),
.B(n_7),
.Y(n_327)
);


endmodule