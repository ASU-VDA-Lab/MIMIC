module real_jpeg_17611_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_560;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B(n_563),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_0),
.B(n_564),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_1),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_1),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_1),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_1),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_1),
.B(n_132),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_1),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_1),
.B(n_187),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_1),
.B(n_316),
.Y(n_315)
);

NAND2x1_ASAP7_75t_L g125 ( 
.A(n_2),
.B(n_53),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_2),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_2),
.B(n_160),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_2),
.B(n_184),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_2),
.B(n_212),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_2),
.B(n_287),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_2),
.B(n_361),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_2),
.B(n_132),
.Y(n_429)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_3),
.Y(n_132)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_3),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_3),
.Y(n_357)
);

BUFx5_ASAP7_75t_L g366 ( 
.A(n_3),
.Y(n_366)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_4),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_4),
.Y(n_147)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_4),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g372 ( 
.A(n_4),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_5),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_6),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_6),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_6),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_6),
.B(n_236),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_6),
.B(n_289),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_6),
.B(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_6),
.B(n_426),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_6),
.B(n_443),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_7),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_7),
.B(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_7),
.B(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_7),
.B(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_7),
.B(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_7),
.B(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_7),
.B(n_473),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_8),
.Y(n_106)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_8),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_8),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_8),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g414 ( 
.A(n_8),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_9),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_9),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_9),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_9),
.B(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_9),
.A2(n_13),
.B1(n_135),
.B2(n_138),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_9),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_9),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_9),
.B(n_149),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_9),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_10),
.B(n_66),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_10),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_10),
.B(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_10),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_10),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_10),
.B(n_252),
.Y(n_251)
);

AND2x2_ASAP7_75t_SL g282 ( 
.A(n_10),
.B(n_132),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_10),
.B(n_306),
.Y(n_305)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_11),
.Y(n_130)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_11),
.Y(n_156)
);

BUFx4f_ASAP7_75t_L g244 ( 
.A(n_11),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_11),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_12),
.B(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_12),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_12),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_12),
.B(n_132),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_12),
.B(n_557),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_13),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_13),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_13),
.B(n_285),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_13),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_13),
.B(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_13),
.B(n_414),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_13),
.B(n_418),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_13),
.B(n_450),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_14),
.Y(n_214)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_14),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_15),
.Y(n_162)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_15),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_15),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_15),
.Y(n_261)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_15),
.Y(n_318)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_15),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_16),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_16),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_16),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_16),
.B(n_151),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_16),
.B(n_232),
.Y(n_231)
);

INVxp33_ASAP7_75t_L g281 ( 
.A(n_16),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_16),
.B(n_312),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_16),
.B(n_364),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g559 ( 
.A(n_18),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_551),
.Y(n_20)
);

OAI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_114),
.B(n_550),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_71),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g550 ( 
.A(n_24),
.B(n_71),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_56),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_42),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_26),
.B(n_42),
.C(n_56),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.C(n_37),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_27),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_43)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_27),
.A2(n_32),
.B1(n_48),
.B2(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_SL g554 ( 
.A(n_27),
.B(n_44),
.C(n_50),
.Y(n_554)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_31),
.Y(n_176)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_31),
.Y(n_233)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_65),
.C(n_68),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_32),
.B(n_69),
.Y(n_108)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_36),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g285 ( 
.A(n_36),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_40),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_50),
.Y(n_42)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_44),
.A2(n_49),
.B1(n_556),
.B2(n_560),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_47),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_47),
.B(n_105),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_47),
.B(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_55),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_61),
.C(n_64),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_57),
.A2(n_58),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_63),
.Y(n_195)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

XOR2x1_ASAP7_75t_L g107 ( 
.A(n_65),
.B(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_68),
.A2(n_69),
.B1(n_104),
.B2(n_304),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_SL g100 ( 
.A(n_69),
.B(n_101),
.C(n_104),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_109),
.C(n_110),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_72),
.B(n_526),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_100),
.C(n_107),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_73),
.B(n_524),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_86),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_79),
.C(n_86),
.Y(n_109)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_84),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.C(n_96),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_87),
.A2(n_88),
.B1(n_92),
.B2(n_93),
.Y(n_515)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_91),
.Y(n_307)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx5_ASAP7_75t_L g412 ( 
.A(n_95),
.Y(n_412)
);

XNOR2x1_ASAP7_75t_L g514 ( 
.A(n_96),
.B(n_515),
.Y(n_514)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_100),
.B(n_107),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_101),
.B(n_519),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_104),
.A2(n_242),
.B1(n_245),
.B2(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_104),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_104),
.B(n_245),
.C(n_305),
.Y(n_520)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_106),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_109),
.B(n_110),
.Y(n_526)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21x1_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_508),
.B(n_545),
.Y(n_114)
);

AO21x2_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_331),
.B(n_505),
.Y(n_115)
);

NOR2xp67_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_297),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_264),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_118),
.B(n_264),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_190),
.Y(n_118)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_119),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_157),
.C(n_177),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_121),
.B(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_133),
.C(n_142),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_122),
.B(n_374),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_125),
.B(n_127),
.C(n_131),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_125),
.B(n_231),
.Y(n_322)
);

MAJx2_ASAP7_75t_L g516 ( 
.A(n_125),
.B(n_231),
.C(n_325),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_133),
.A2(n_134),
.B1(n_142),
.B2(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_134),
.A2(n_347),
.B(n_352),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx6_ASAP7_75t_L g423 ( 
.A(n_136),
.Y(n_423)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_137),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_141),
.Y(n_184)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_141),
.Y(n_351)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_142),
.Y(n_375)
);

MAJx2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_148),
.C(n_152),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_143),
.A2(n_144),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_143),
.A2(n_144),
.B1(n_152),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g323 ( 
.A(n_144),
.B(n_197),
.C(n_242),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_146),
.Y(n_312)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_148),
.B(n_277),
.Y(n_276)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_152),
.Y(n_278)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_154),
.B(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_156),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_157),
.A2(n_178),
.B1(n_179),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_157),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_169),
.C(n_172),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_158),
.B(n_292),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.C(n_166),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_159),
.A2(n_166),
.B1(n_344),
.B2(n_345),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_159),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_159),
.B(n_409),
.Y(n_408)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_163),
.B(n_343),
.Y(n_342)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_165),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_166),
.Y(n_345)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_169),
.A2(n_170),
.B1(n_172),
.B2(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_172),
.Y(n_293)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_180),
.B(n_182),
.C(n_186),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_185),
.B2(n_186),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_182),
.A2(n_183),
.B1(n_368),
.B2(n_369),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_183),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_183),
.Y(n_367)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_189),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_238),
.B1(n_262),
.B2(n_263),
.Y(n_190)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_191),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_226),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_192),
.B(n_227),
.C(n_228),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_202),
.C(n_215),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_193),
.B(n_202),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_194),
.B(n_197),
.C(n_199),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_201),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_197),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_197),
.A2(n_201),
.B1(n_242),
.B2(n_245),
.Y(n_241)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.C(n_210),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_203),
.A2(n_210),
.B1(n_211),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_203),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_205),
.B(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_209),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_210),
.B(n_387),
.C(n_389),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_210),
.A2(n_211),
.B1(n_387),
.B2(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2x2_ASAP7_75t_SL g270 ( 
.A(n_215),
.B(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_220),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_221),
.C(n_225),
.Y(n_237)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_225),
.Y(n_220)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_237),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_234),
.B2(n_235),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_230),
.B(n_235),
.C(n_237),
.Y(n_326)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_238),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_246),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_239),
.B(n_247),
.C(n_248),
.Y(n_327)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_242),
.Y(n_245)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_244),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_244),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_249),
.B(n_251),
.C(n_258),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_258),
.Y(n_250)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_262),
.B(n_329),
.C(n_330),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_270),
.C(n_272),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_266),
.A2(n_267),
.B1(n_270),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_270),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_273),
.B(n_335),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_291),
.C(n_294),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_274),
.B(n_340),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_279),
.C(n_283),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_276),
.B(n_398),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_279),
.B(n_283),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_280),
.B(n_282),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.C(n_288),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_284),
.A2(n_286),
.B1(n_383),
.B2(n_384),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_284),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_286),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_286),
.A2(n_384),
.B1(n_459),
.B2(n_460),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_286),
.B(n_455),
.C(n_459),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_288),
.B(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_291),
.B(n_294),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_297),
.A2(n_506),
.B(n_507),
.Y(n_505)
);

AND2x2_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_328),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_298),
.B(n_328),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_299),
.B(n_301),
.C(n_319),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_319),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_308),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_302),
.B(n_309),
.C(n_310),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_305),
.Y(n_302)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_313),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_311),
.B(n_314),
.C(n_315),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

INVx6_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_327),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_326),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_321),
.B(n_326),
.C(n_539),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_323),
.B1(n_324),
.B2(n_325),
.Y(n_321)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_322),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_323),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_327),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_401),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_337),
.C(n_376),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_334),
.B(n_338),
.Y(n_504)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_341),
.C(n_373),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_339),
.B(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_341),
.B(n_373),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_346),
.C(n_358),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_342),
.B(n_346),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_344),
.B(n_410),
.C(n_413),
.Y(n_434)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

INVx5_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_358),
.B(n_379),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_367),
.C(n_368),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g490 ( 
.A(n_359),
.B(n_491),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_363),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_360),
.B(n_363),
.Y(n_441)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_360),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_360),
.A2(n_448),
.B1(n_449),
.B2(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

NOR2x1_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_399),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_377),
.B(n_399),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_380),
.C(n_396),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_378),
.B(n_502),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_380),
.B(n_397),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_385),
.C(n_394),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_381),
.B(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_386),
.B(n_395),
.Y(n_496)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_387),
.Y(n_437)
);

XOR2x2_ASAP7_75t_L g435 ( 
.A(n_389),
.B(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_393),
.Y(n_461)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

NAND3xp33_ASAP7_75t_SL g401 ( 
.A(n_402),
.B(n_403),
.C(n_504),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_404),
.A2(n_499),
.B(n_503),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_485),
.B(n_498),
.Y(n_404)
);

OAI21x1_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_444),
.B(n_484),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_432),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_407),
.B(n_432),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_415),
.C(n_424),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_408),
.B(n_480),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_413),
.Y(n_409)
);

INVx5_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_414),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_415),
.A2(n_416),
.B1(n_424),
.B2(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_421),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_417),
.B(n_421),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx4_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx6_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_424),
.Y(n_481)
);

AO22x1_ASAP7_75t_SL g424 ( 
.A1(n_425),
.A2(n_429),
.B1(n_430),
.B2(n_431),
.Y(n_424)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_425),
.Y(n_430)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_429),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_429),
.B(n_430),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_431),
.B(n_472),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_438),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_435),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_434),
.B(n_435),
.C(n_438),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

MAJx2_ASAP7_75t_L g493 ( 
.A(n_439),
.B(n_441),
.C(n_442),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_445),
.A2(n_478),
.B(n_483),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_446),
.A2(n_462),
.B(n_477),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_454),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_447),
.B(n_454),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_448),
.B(n_449),
.Y(n_447)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_449),
.Y(n_470)
);

INVx4_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx4_ASAP7_75t_SL g451 ( 
.A(n_452),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_455),
.A2(n_456),
.B1(n_457),
.B2(n_458),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_463),
.A2(n_471),
.B(n_476),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_469),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_464),
.B(n_469),
.Y(n_476)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_479),
.B(n_482),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_479),
.B(n_482),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_486),
.B(n_497),
.Y(n_485)
);

NOR2xp67_ASAP7_75t_SL g498 ( 
.A(n_486),
.B(n_497),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_487),
.A2(n_488),
.B1(n_494),
.B2(n_495),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_489),
.A2(n_490),
.B1(n_492),
.B2(n_493),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_493),
.C(n_494),
.Y(n_500)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

NOR2x1_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_501),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_500),
.B(n_501),
.Y(n_503)
);

NOR3xp33_ASAP7_75t_SL g508 ( 
.A(n_509),
.B(n_527),
.C(n_540),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_509),
.A2(n_546),
.B(n_549),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_510),
.B(n_525),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_510),
.B(n_525),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_517),
.C(n_522),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_511),
.B(n_530),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_514),
.C(n_516),
.Y(n_511)
);

INVxp33_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_513),
.B(n_535),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_514),
.B(n_516),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_517),
.A2(n_522),
.B1(n_523),
.B2(n_531),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_517),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_520),
.C(n_521),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_518),
.B(n_537),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_520),
.B(n_521),
.Y(n_537)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_528),
.A2(n_547),
.B(n_548),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_529),
.B(n_532),
.Y(n_528)
);

NOR2xp67_ASAP7_75t_SL g548 ( 
.A(n_529),
.B(n_532),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_536),
.C(n_538),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_533),
.A2(n_534),
.B1(n_536),
.B2(n_544),
.Y(n_543)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_536),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_538),
.B(n_543),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_541),
.B(n_542),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_541),
.B(n_542),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_R g551 ( 
.A(n_552),
.B(n_562),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_553),
.B(n_561),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_553),
.B(n_561),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_554),
.B(n_555),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_556),
.Y(n_560)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);


endmodule