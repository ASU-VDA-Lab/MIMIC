module fake_jpeg_29313_n_550 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_550);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_550;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_33),
.B(n_9),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_62),
.B(n_66),
.Y(n_150)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_65),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_33),
.B(n_10),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_67),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_28),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g152 ( 
.A(n_69),
.B(n_61),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_23),
.B(n_10),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_70),
.B(n_72),
.Y(n_122)
);

BUFx8_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_71),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_36),
.B(n_8),
.Y(n_72)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_73),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_36),
.B(n_8),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_76),
.B(n_85),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_77),
.Y(n_143)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_41),
.B(n_48),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_41),
.B(n_8),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_46),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_91),
.B(n_100),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_92),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_93),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_42),
.B(n_11),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

BUFx10_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_70),
.A2(n_42),
.B1(n_48),
.B2(n_47),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_108),
.A2(n_129),
.B1(n_141),
.B2(n_151),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_109),
.B(n_152),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_46),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_110),
.B(n_128),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_104),
.A2(n_51),
.B1(n_40),
.B2(n_49),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_117),
.A2(n_121),
.B1(n_127),
.B2(n_153),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_104),
.A2(n_51),
.B1(n_40),
.B2(n_49),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_56),
.A2(n_51),
.B1(n_82),
.B2(n_96),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_71),
.B(n_47),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_54),
.A2(n_50),
.B1(n_27),
.B2(n_45),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_71),
.A2(n_50),
.B(n_27),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_138),
.A2(n_139),
.B(n_164),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_83),
.A2(n_50),
.B1(n_27),
.B2(n_45),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_65),
.A2(n_34),
.B1(n_45),
.B2(n_44),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_67),
.A2(n_34),
.B1(n_44),
.B2(n_43),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_95),
.A2(n_102),
.B1(n_101),
.B2(n_58),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_68),
.A2(n_34),
.B1(n_44),
.B2(n_43),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_154),
.A2(n_60),
.B1(n_74),
.B2(n_87),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_55),
.A2(n_43),
.B1(n_38),
.B2(n_26),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_80),
.B(n_38),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_19),
.Y(n_179)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_169),
.Y(n_259)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_122),
.A2(n_19),
.B(n_38),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_170),
.Y(n_272)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_172),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_117),
.Y(n_173)
);

INVx6_ASAP7_75t_SL g279 ( 
.A(n_173),
.Y(n_279)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_174),
.Y(n_235)
);

BUFx4f_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

INVx11_ASAP7_75t_L g239 ( 
.A(n_176),
.Y(n_239)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_107),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_178),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_179),
.B(n_210),
.Y(n_264)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_130),
.Y(n_181)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_181),
.Y(n_244)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_130),
.Y(n_182)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_182),
.Y(n_254)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_135),
.Y(n_183)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_183),
.Y(n_240)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_135),
.Y(n_184)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_184),
.Y(n_257)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_119),
.Y(n_185)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_185),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_19),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_186),
.B(n_191),
.Y(n_251)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_132),
.A2(n_94),
.B1(n_93),
.B2(n_77),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_189),
.A2(n_212),
.B1(n_218),
.B2(n_230),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_123),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_190),
.B(n_192),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_26),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_125),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_134),
.Y(n_193)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_193),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_166),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_194),
.B(n_197),
.Y(n_255)
);

INVx4_ASAP7_75t_SL g195 ( 
.A(n_126),
.Y(n_195)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_195),
.Y(n_245)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_136),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_196),
.B(n_204),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_140),
.B(n_26),
.Y(n_197)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_142),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_199),
.Y(n_275)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_112),
.Y(n_200)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_200),
.Y(n_274)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_106),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_201),
.Y(n_269)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_202),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_115),
.B(n_124),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_203),
.B(n_226),
.Y(n_265)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

BUFx12_ASAP7_75t_L g205 ( 
.A(n_119),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_205),
.B(n_208),
.Y(n_258)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_145),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_206),
.Y(n_262)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_145),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_207),
.Y(n_278)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_126),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_209),
.A2(n_213),
.B1(n_215),
.B2(n_220),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_113),
.B(n_73),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_157),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_211),
.B(n_214),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_107),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_158),
.A2(n_92),
.B1(n_88),
.B2(n_118),
.Y(n_213)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_158),
.A2(n_77),
.B1(n_49),
.B2(n_40),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_216),
.B(n_217),
.Y(n_261)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_162),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_132),
.A2(n_37),
.B1(n_73),
.B2(n_91),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_163),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_219),
.B(n_221),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_118),
.A2(n_37),
.B1(n_91),
.B2(n_12),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_163),
.Y(n_221)
);

BUFx8_ASAP7_75t_L g222 ( 
.A(n_137),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_222),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_161),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_223),
.B(n_225),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_L g224 ( 
.A1(n_144),
.A2(n_7),
.B1(n_17),
.B2(n_16),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_224),
.A2(n_144),
.B1(n_156),
.B2(n_168),
.Y(n_231)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_147),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_146),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_105),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_227),
.B(n_228),
.Y(n_267)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_161),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_160),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_229),
.B(n_113),
.Y(n_232)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_105),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_231),
.A2(n_213),
.B1(n_220),
.B2(n_215),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_232),
.Y(n_324)
);

OR2x2_ASAP7_75t_SL g238 ( 
.A(n_170),
.B(n_121),
.Y(n_238)
);

OAI21xp33_ASAP7_75t_L g296 ( 
.A1(n_238),
.A2(n_148),
.B(n_222),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_180),
.B(n_114),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_243),
.B(n_249),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_171),
.B(n_114),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_198),
.B(n_116),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_252),
.B(n_256),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_173),
.A2(n_175),
.B1(n_188),
.B2(n_184),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_253),
.A2(n_279),
.B1(n_268),
.B2(n_272),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_175),
.B(n_116),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_224),
.B(n_168),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_266),
.B(n_273),
.Y(n_302)
);

FAx1_ASAP7_75t_SL g268 ( 
.A(n_210),
.B(n_127),
.CI(n_153),
.CON(n_268),
.SN(n_268)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_268),
.B(n_276),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_225),
.B(n_111),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_181),
.B(n_14),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_188),
.B(n_160),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_280),
.B(n_7),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_182),
.B(n_111),
.C(n_167),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_149),
.C(n_185),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_195),
.A2(n_167),
.B1(n_149),
.B2(n_137),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_282),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_283),
.A2(n_289),
.B1(n_295),
.B2(n_318),
.Y(n_336)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_273),
.Y(n_284)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_284),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_286),
.B(n_310),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_176),
.C(n_218),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_287),
.B(n_258),
.C(n_241),
.Y(n_334)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_247),
.Y(n_288)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_288),
.Y(n_347)
);

OAI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_272),
.A2(n_183),
.B1(n_223),
.B2(n_214),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_249),
.B(n_148),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_290),
.B(n_303),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_291),
.A2(n_299),
.B1(n_300),
.B2(n_326),
.Y(n_348)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_247),
.Y(n_292)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_292),
.Y(n_351)
);

INVx6_ASAP7_75t_L g293 ( 
.A(n_242),
.Y(n_293)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_293),
.Y(n_341)
);

OAI22xp33_ASAP7_75t_L g295 ( 
.A1(n_252),
.A2(n_189),
.B1(n_212),
.B2(n_178),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_296),
.A2(n_263),
.B(n_250),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_242),
.Y(n_297)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_297),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_243),
.A2(n_222),
.B(n_11),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_298),
.A2(n_308),
.B(n_319),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_264),
.A2(n_7),
.B1(n_18),
.B2(n_16),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_264),
.A2(n_6),
.B1(n_18),
.B2(n_15),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_236),
.B(n_205),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_301),
.B(n_305),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_0),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_262),
.Y(n_304)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_304),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_246),
.B(n_205),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_267),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_306),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_251),
.B(n_0),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_307),
.B(n_309),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_238),
.A2(n_5),
.B(n_15),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_268),
.B(n_256),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_260),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_311),
.B(n_312),
.Y(n_353)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_262),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_275),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_313),
.B(n_320),
.Y(n_344)
);

OAI21xp33_ASAP7_75t_L g314 ( 
.A1(n_255),
.A2(n_7),
.B(n_15),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_314),
.A2(n_241),
.B1(n_245),
.B2(n_254),
.Y(n_335)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_278),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_315),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_279),
.A2(n_4),
.B1(n_15),
.B2(n_14),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_317),
.A2(n_297),
.B1(n_293),
.B2(n_311),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_248),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_280),
.A2(n_3),
.B1(n_4),
.B2(n_13),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_261),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_270),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_321),
.B(n_235),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_248),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_322),
.A2(n_325),
.B1(n_328),
.B2(n_329),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_232),
.A2(n_3),
.B(n_4),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_323),
.A2(n_254),
.B(n_244),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_266),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_277),
.A2(n_13),
.B1(n_18),
.B2(n_259),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_281),
.A2(n_13),
.B1(n_269),
.B2(n_259),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_269),
.A2(n_233),
.B1(n_276),
.B2(n_271),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_302),
.A2(n_269),
.B1(n_233),
.B2(n_250),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_333),
.A2(n_364),
.B1(n_365),
.B2(n_367),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_334),
.B(n_360),
.C(n_362),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_335),
.B(n_350),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_327),
.A2(n_245),
.B1(n_263),
.B2(n_234),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_340),
.A2(n_342),
.B(n_358),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_346),
.A2(n_349),
.B(n_369),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_309),
.A2(n_244),
.B(n_234),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_302),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_352),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_329),
.Y(n_354)
);

CKINVDCx14_ASAP7_75t_R g376 ( 
.A(n_354),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_318),
.A2(n_257),
.B1(n_274),
.B2(n_242),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_357),
.A2(n_361),
.B1(n_292),
.B2(n_293),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_324),
.A2(n_257),
.B1(n_240),
.B2(n_274),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_284),
.B(n_235),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_359),
.B(n_325),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_309),
.B(n_237),
.C(n_278),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_322),
.A2(n_237),
.B1(n_240),
.B2(n_239),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_285),
.B(n_239),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_316),
.A2(n_285),
.B(n_291),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_363),
.A2(n_323),
.B(n_300),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_294),
.A2(n_290),
.B1(n_324),
.B2(n_287),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_294),
.A2(n_298),
.B1(n_326),
.B2(n_316),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_288),
.Y(n_366)
);

CKINVDCx14_ASAP7_75t_R g378 ( 
.A(n_366),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_306),
.A2(n_286),
.B1(n_319),
.B2(n_321),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_320),
.A2(n_310),
.B1(n_283),
.B2(n_303),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_370),
.A2(n_364),
.B1(n_348),
.B2(n_367),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_330),
.B(n_307),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_371),
.B(n_383),
.C(n_402),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_344),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_375),
.B(n_397),
.Y(n_409)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_347),
.Y(n_377)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_377),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_355),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_379),
.B(n_384),
.Y(n_417)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_347),
.Y(n_380)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_380),
.Y(n_419)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_351),
.Y(n_381)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_381),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_334),
.B(n_313),
.C(n_328),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_385),
.B(n_374),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_345),
.B(n_308),
.Y(n_386)
);

NAND3xp33_ASAP7_75t_L g413 ( 
.A(n_386),
.B(n_405),
.C(n_400),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_387),
.A2(n_391),
.B1(n_403),
.B2(n_366),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_349),
.A2(n_304),
.B(n_312),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_388),
.A2(n_390),
.B(n_392),
.Y(n_430)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_351),
.Y(n_389)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_389),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_331),
.A2(n_299),
.B(n_315),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_354),
.A2(n_297),
.B1(n_343),
.B2(n_352),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_331),
.A2(n_365),
.B(n_346),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_359),
.Y(n_393)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_393),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_395),
.A2(n_401),
.B1(n_360),
.B2(n_332),
.Y(n_418)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_350),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_396),
.Y(n_423)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_344),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_353),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_398),
.B(n_399),
.Y(n_415)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_353),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_332),
.B(n_339),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_400),
.B(n_404),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_348),
.A2(n_370),
.B1(n_333),
.B2(n_338),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_330),
.B(n_362),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_343),
.A2(n_336),
.B1(n_363),
.B2(n_338),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_356),
.Y(n_404)
);

OA21x2_ASAP7_75t_L g406 ( 
.A1(n_394),
.A2(n_339),
.B(n_336),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_406),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_378),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_407),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_408),
.B(n_372),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_378),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_411),
.B(n_429),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_394),
.A2(n_334),
.B(n_369),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_412),
.A2(n_430),
.B(n_408),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_413),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_414),
.A2(n_435),
.B1(n_437),
.B2(n_396),
.Y(n_443)
);

OAI21xp33_ASAP7_75t_L g416 ( 
.A1(n_386),
.A2(n_345),
.B(n_368),
.Y(n_416)
);

NAND3xp33_ASAP7_75t_L g452 ( 
.A(n_416),
.B(n_421),
.C(n_415),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_418),
.A2(n_431),
.B1(n_432),
.B2(n_384),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_405),
.B(n_362),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_420),
.B(n_424),
.Y(n_451)
);

HAxp5_ASAP7_75t_SL g421 ( 
.A(n_392),
.B(n_342),
.CON(n_421),
.SN(n_421)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_375),
.B(n_360),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_397),
.B(n_368),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_427),
.Y(n_463)
);

CKINVDCx14_ASAP7_75t_R g428 ( 
.A(n_388),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_428),
.B(n_382),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_377),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_376),
.A2(n_357),
.B1(n_361),
.B2(n_358),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_401),
.A2(n_376),
.B1(n_372),
.B2(n_395),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_380),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_433),
.B(n_399),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_403),
.A2(n_355),
.B1(n_337),
.B2(n_341),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_391),
.A2(n_337),
.B1(n_341),
.B2(n_356),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_438),
.A2(n_450),
.B1(n_464),
.B2(n_406),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_440),
.A2(n_452),
.B(n_448),
.Y(n_472)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_441),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_443),
.A2(n_454),
.B1(n_420),
.B2(n_409),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_444),
.B(n_435),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_426),
.B(n_373),
.C(n_383),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_445),
.B(n_456),
.C(n_424),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_407),
.B(n_398),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_446),
.B(n_448),
.Y(n_466)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_427),
.Y(n_447)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_447),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_411),
.B(n_413),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_415),
.B(n_393),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_449),
.B(n_453),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_432),
.A2(n_418),
.B1(n_431),
.B2(n_430),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_429),
.B(n_389),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_414),
.A2(n_390),
.B1(n_374),
.B2(n_382),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_455),
.A2(n_417),
.B(n_425),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_426),
.B(n_373),
.C(n_402),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_433),
.B(n_381),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_458),
.B(n_461),
.Y(n_465)
);

AOI322xp5_ASAP7_75t_L g460 ( 
.A1(n_412),
.A2(n_385),
.A3(n_387),
.B1(n_402),
.B2(n_404),
.C1(n_371),
.C2(n_335),
.Y(n_460)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_460),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_409),
.B(n_379),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_425),
.B(n_371),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_462),
.B(n_419),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_428),
.A2(n_340),
.B1(n_423),
.B2(n_436),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_468),
.B(n_474),
.C(n_475),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_470),
.A2(n_476),
.B1(n_459),
.B2(n_449),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_471),
.B(n_473),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_472),
.A2(n_477),
.B(n_481),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_445),
.B(n_417),
.C(n_423),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_456),
.B(n_436),
.C(n_437),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_454),
.A2(n_406),
.B1(n_410),
.B2(n_419),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_440),
.A2(n_406),
.B(n_410),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_478),
.B(n_479),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_457),
.B(n_422),
.Y(n_480)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_480),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_442),
.A2(n_455),
.B(n_464),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_444),
.B(n_422),
.C(n_434),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_483),
.B(n_457),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_462),
.B(n_434),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_485),
.B(n_486),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_451),
.B(n_450),
.Y(n_486)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_480),
.Y(n_489)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_489),
.Y(n_511)
);

XNOR2x1_ASAP7_75t_L g490 ( 
.A(n_483),
.B(n_460),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_490),
.B(n_496),
.Y(n_514)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_469),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_491),
.A2(n_495),
.B1(n_498),
.B2(n_503),
.Y(n_507)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_469),
.Y(n_495)
);

NOR3xp33_ASAP7_75t_L g497 ( 
.A(n_466),
.B(n_452),
.C(n_446),
.Y(n_497)
);

NAND3xp33_ASAP7_75t_L g512 ( 
.A(n_497),
.B(n_502),
.C(n_465),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_467),
.A2(n_438),
.B1(n_459),
.B2(n_449),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_466),
.B(n_441),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_499),
.B(n_501),
.Y(n_513)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_482),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_465),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_482),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_504),
.B(n_494),
.C(n_493),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_500),
.A2(n_481),
.B(n_477),
.Y(n_505)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_505),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_489),
.A2(n_476),
.B1(n_467),
.B2(n_472),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_506),
.A2(n_518),
.B1(n_504),
.B2(n_487),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_508),
.B(n_492),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_500),
.A2(n_470),
.B(n_484),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_509),
.B(n_512),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_488),
.B(n_468),
.C(n_475),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_510),
.B(n_516),
.C(n_517),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_491),
.A2(n_473),
.B(n_484),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_515),
.A2(n_439),
.B(n_503),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_488),
.B(n_474),
.C(n_490),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_494),
.B(n_486),
.C(n_471),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_495),
.A2(n_447),
.B1(n_463),
.B2(n_479),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_514),
.B(n_487),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_519),
.B(n_520),
.Y(n_533)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_521),
.Y(n_530)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_524),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_514),
.B(n_492),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_525),
.B(n_526),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_510),
.B(n_485),
.C(n_478),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_516),
.B(n_443),
.C(n_451),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_528),
.B(n_529),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_506),
.B(n_439),
.Y(n_529)
);

BUFx24_ASAP7_75t_SL g534 ( 
.A(n_520),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_534),
.A2(n_536),
.B1(n_527),
.B2(n_511),
.Y(n_540)
);

AOI31xp33_ASAP7_75t_L g536 ( 
.A1(n_527),
.A2(n_523),
.A3(n_522),
.B(n_513),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_531),
.B(n_523),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_537),
.B(n_538),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_533),
.B(n_530),
.C(n_535),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_532),
.B(n_508),
.Y(n_539)
);

OAI31xp33_ASAP7_75t_SL g542 ( 
.A1(n_539),
.A2(n_540),
.A3(n_526),
.B(n_513),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_542),
.A2(n_528),
.B(n_539),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_541),
.B(n_538),
.C(n_537),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_543),
.A2(n_544),
.B(n_515),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_545),
.B(n_511),
.C(n_509),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_546),
.B(n_507),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_547),
.B(n_453),
.C(n_458),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_548),
.B(n_518),
.Y(n_549)
);

O2A1O1Ixp33_ASAP7_75t_SL g550 ( 
.A1(n_549),
.A2(n_505),
.B(n_461),
.C(n_517),
.Y(n_550)
);


endmodule