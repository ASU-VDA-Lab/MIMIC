module fake_netlist_1_8259_n_20 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_20);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_20;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_7;
NAND2xp5_ASAP7_75t_SL g7 ( .A(n_2), .B(n_6), .Y(n_7) );
BUFx6f_ASAP7_75t_L g8 ( .A(n_5), .Y(n_8) );
CKINVDCx16_ASAP7_75t_R g9 ( .A(n_1), .Y(n_9) );
INVx3_ASAP7_75t_L g10 ( .A(n_3), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
CKINVDCx16_ASAP7_75t_R g13 ( .A(n_9), .Y(n_13) );
AOI21xp5_ASAP7_75t_L g14 ( .A1(n_7), .A2(n_0), .B(n_4), .Y(n_14) );
HB1xp67_ASAP7_75t_L g15 ( .A(n_12), .Y(n_15) );
BUFx2_ASAP7_75t_L g16 ( .A(n_13), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_15), .B(n_14), .Y(n_17) );
OAI31xp33_ASAP7_75t_L g18 ( .A1(n_17), .A2(n_15), .A3(n_16), .B(n_11), .Y(n_18) );
CKINVDCx20_ASAP7_75t_R g19 ( .A(n_18), .Y(n_19) );
CKINVDCx5p33_ASAP7_75t_R g20 ( .A(n_19), .Y(n_20) );
endmodule