module real_jpeg_32194_n_3 (n_1, n_0, n_2, n_3);

input n_1;
input n_0;
input n_2;

output n_3;

wire n_5;
wire n_8;
wire n_4;
wire n_6;
wire n_7;
wire n_10;
wire n_9;

BUFx2_ASAP7_75t_R g5 ( 
.A(n_0),
.Y(n_5)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx2_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_SL g3 ( 
.A1(n_4),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_3)
);

CKINVDCx14_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

OAI21xp5_ASAP7_75t_SL g4 ( 
.A1(n_5),
.A2(n_6),
.B(n_7),
.Y(n_4)
);

NAND2xp33_ASAP7_75t_SL g7 ( 
.A(n_5),
.B(n_6),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_9),
.Y(n_8)
);


endmodule