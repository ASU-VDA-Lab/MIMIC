module fake_jpeg_27692_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

CKINVDCx6p67_ASAP7_75t_R g64 ( 
.A(n_36),
.Y(n_64)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx2_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_20),
.Y(n_41)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_8),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_46),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx5_ASAP7_75t_SL g110 ( 
.A(n_49),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_19),
.B1(n_23),
.B2(n_17),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_50),
.A2(n_51),
.B1(n_58),
.B2(n_32),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_19),
.B1(n_23),
.B2(n_17),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_23),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_57),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_46),
.A2(n_25),
.B1(n_22),
.B2(n_21),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_53),
.A2(n_29),
.B1(n_26),
.B2(n_33),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_68),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_35),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_17),
.B1(n_35),
.B2(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_63),
.Y(n_80)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_65),
.Y(n_104)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_30),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_39),
.A2(n_35),
.B1(n_16),
.B2(n_33),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_69),
.A2(n_33),
.B1(n_42),
.B2(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_16),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_72),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_36),
.B(n_16),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_45),
.Y(n_88)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_76),
.A2(n_94),
.B1(n_91),
.B2(n_97),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_53),
.B(n_30),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_78),
.B(n_83),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_26),
.B1(n_29),
.B2(n_42),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_79),
.A2(n_90),
.B1(n_102),
.B2(n_64),
.Y(n_138)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_28),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_52),
.B(n_39),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_27),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_103),
.Y(n_114)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_88),
.B(n_31),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_65),
.A2(n_42),
.B1(n_67),
.B2(n_60),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_36),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_94),
.C(n_64),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_36),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_95),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_36),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_36),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_48),
.Y(n_96)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_55),
.B(n_28),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_100),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_28),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_36),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_106),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_60),
.A2(n_24),
.B1(n_32),
.B2(n_15),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_111),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_59),
.A2(n_32),
.B1(n_24),
.B2(n_27),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_18),
.Y(n_119)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_132),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_63),
.C(n_62),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_123),
.C(n_95),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_122),
.B(n_141),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_120),
.A2(n_109),
.B1(n_85),
.B2(n_88),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_94),
.A2(n_62),
.B(n_1),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_64),
.C(n_73),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_80),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_125),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_80),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_133),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_93),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_134),
.B(n_135),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_98),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_82),
.B(n_32),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_136),
.B(n_137),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_78),
.B(n_24),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_81),
.Y(n_143)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_143),
.Y(n_201)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_144),
.B(n_145),
.Y(n_198)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_151),
.Y(n_178)
);

BUFx12_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_147),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_31),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_140),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_171),
.Y(n_181)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_91),
.B1(n_76),
.B2(n_77),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_152),
.A2(n_156),
.B1(n_163),
.B2(n_175),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_86),
.C(n_77),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_153),
.B(n_157),
.C(n_124),
.Y(n_206)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_161),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_114),
.A2(n_86),
.B1(n_92),
.B2(n_110),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_132),
.C(n_116),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_159),
.A2(n_141),
.B1(n_112),
.B2(n_121),
.Y(n_185)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_115),
.B(n_108),
.Y(n_162)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_162),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_114),
.A2(n_110),
.B1(n_106),
.B2(n_74),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_108),
.Y(n_164)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_170),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_122),
.A2(n_96),
.B1(n_75),
.B2(n_111),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_167),
.A2(n_124),
.B1(n_131),
.B2(n_34),
.Y(n_191)
);

OAI32xp33_ASAP7_75t_L g169 ( 
.A1(n_129),
.A2(n_101),
.A3(n_107),
.B1(n_105),
.B2(n_104),
.Y(n_169)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_126),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_117),
.B(n_104),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_138),
.A2(n_96),
.B1(n_99),
.B2(n_11),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_172),
.A2(n_168),
.B1(n_146),
.B2(n_121),
.Y(n_188)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_120),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_174),
.Y(n_184)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_119),
.A2(n_99),
.B1(n_34),
.B2(n_18),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_113),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_177),
.B(n_183),
.Y(n_228)
);

OAI22x1_ASAP7_75t_SL g180 ( 
.A1(n_160),
.A2(n_119),
.B1(n_133),
.B2(n_125),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_180),
.A2(n_185),
.B1(n_188),
.B2(n_175),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_160),
.A2(n_113),
.B1(n_112),
.B2(n_135),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_182),
.A2(n_192),
.B1(n_207),
.B2(n_166),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_141),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_31),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_186),
.B(n_194),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_173),
.A2(n_131),
.B(n_27),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_190),
.A2(n_197),
.B(n_199),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_191),
.A2(n_170),
.B1(n_165),
.B2(n_154),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_161),
.A2(n_124),
.B1(n_34),
.B2(n_18),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_206),
.C(n_142),
.Y(n_208)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_169),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_195),
.B(n_196),
.Y(n_233)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_163),
.Y(n_196)
);

XNOR2x1_ASAP7_75t_L g197 ( 
.A(n_142),
.B(n_34),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_148),
.A2(n_0),
.B(n_1),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_148),
.A2(n_0),
.B(n_1),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_200),
.A2(n_2),
.B(n_3),
.Y(n_229)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_174),
.Y(n_204)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_204),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_144),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_209),
.C(n_215),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_177),
.C(n_183),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_226),
.B1(n_207),
.B2(n_196),
.Y(n_237)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_214),
.Y(n_249)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_153),
.C(n_145),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_187),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_216),
.B(n_222),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_217),
.A2(n_220),
.B1(n_194),
.B2(n_189),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_179),
.A2(n_159),
.B1(n_156),
.B2(n_151),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_221),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_179),
.A2(n_152),
.B1(n_10),
.B2(n_11),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_178),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_224),
.Y(n_236)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_176),
.A2(n_150),
.B1(n_147),
.B2(n_9),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_225),
.A2(n_234),
.B1(n_12),
.B2(n_13),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_195),
.A2(n_147),
.B1(n_3),
.B2(n_4),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_180),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_231),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_229),
.A2(n_230),
.B(n_4),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_184),
.A2(n_190),
.B(n_185),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_201),
.B(n_10),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_176),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_237),
.A2(n_239),
.B1(n_251),
.B2(n_253),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_232),
.A2(n_192),
.B1(n_198),
.B2(n_197),
.Y(n_239)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_241),
.B(n_246),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_189),
.C(n_204),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_243),
.C(n_218),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_205),
.C(n_203),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_200),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_247),
.Y(n_267)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_215),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_248),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_199),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_252),
.Y(n_271)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_186),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_227),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_211),
.B(n_220),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_SL g270 ( 
.A(n_255),
.B(n_229),
.C(n_234),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_224),
.C(n_211),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_259),
.B(n_272),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_261),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_230),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_247),
.C(n_243),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_269),
.C(n_275),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_245),
.B(n_233),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_274),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_268),
.A2(n_270),
.B(n_256),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_212),
.C(n_214),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_222),
.C(n_221),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_236),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_5),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_13),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_239),
.B(n_14),
.C(n_5),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_238),
.B(n_14),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_5),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_266),
.A2(n_256),
.B1(n_254),
.B2(n_253),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_277),
.A2(n_260),
.B1(n_265),
.B2(n_271),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_262),
.Y(n_278)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_278),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_279),
.A2(n_286),
.B(n_289),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_258),
.A2(n_255),
.B(n_244),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_280),
.A2(n_6),
.B(n_7),
.Y(n_301)
);

INVx13_ASAP7_75t_L g282 ( 
.A(n_276),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_282),
.B(n_287),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_237),
.Y(n_283)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_264),
.B(n_4),
.Y(n_288)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_288),
.Y(n_299)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_291),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_292),
.A2(n_290),
.B1(n_280),
.B2(n_7),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_263),
.C(n_267),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_296),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_295),
.A2(n_298),
.B1(n_286),
.B2(n_292),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_267),
.C(n_271),
.Y(n_296)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_301),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_7),
.C(n_281),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_291),
.Y(n_309)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_305),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_295),
.A2(n_278),
.B1(n_282),
.B2(n_277),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_306),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_SL g308 ( 
.A(n_294),
.B(n_284),
.C(n_281),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_309),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_299),
.B(n_290),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_312),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_301),
.C(n_302),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_297),
.B1(n_300),
.B2(n_293),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_318),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_312),
.B(n_296),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_307),
.C(n_316),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_319),
.A2(n_314),
.B(n_315),
.Y(n_323)
);

BUFx4f_ASAP7_75t_SL g320 ( 
.A(n_314),
.Y(n_320)
);

AND2x4_ASAP7_75t_SL g322 ( 
.A(n_320),
.B(n_305),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_322),
.A2(n_323),
.B(n_321),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_306),
.C(n_311),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_325),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_326),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_304),
.Y(n_328)
);


endmodule