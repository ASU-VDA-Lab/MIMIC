module fake_jpeg_3636_n_202 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_202);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_9),
.B(n_13),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_44),
.Y(n_53)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_19),
.Y(n_55)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_47),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_31),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_57),
.Y(n_80)
);

CKINVDCx12_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_55),
.B(n_65),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_26),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_26),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_0),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_66),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_36),
.A2(n_17),
.B1(n_27),
.B2(n_23),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_36),
.A2(n_17),
.B1(n_27),
.B2(n_23),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_42),
.B1(n_23),
.B2(n_18),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_40),
.B(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_20),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_25),
.B1(n_24),
.B2(n_22),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_39),
.B1(n_41),
.B2(n_48),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_41),
.A2(n_30),
.B1(n_23),
.B2(n_18),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_0),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_49),
.B(n_24),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_22),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_74),
.Y(n_86)
);

CKINVDCx12_ASAP7_75t_R g75 ( 
.A(n_47),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_87),
.Y(n_107)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_39),
.B(n_30),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_81),
.A2(n_85),
.B1(n_89),
.B2(n_102),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_42),
.B1(n_18),
.B2(n_30),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_53),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_46),
.C(n_1),
.Y(n_88)
);

FAx1_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_94),
.CI(n_73),
.CON(n_109),
.SN(n_109)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_1),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVxp67_ASAP7_75t_SL g112 ( 
.A(n_93),
.Y(n_112)
);

OR2x4_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_54),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_1),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_102),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_69),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_101),
.A2(n_56),
.B1(n_68),
.B2(n_61),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_2),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_110),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_94),
.A2(n_50),
.B1(n_68),
.B2(n_56),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_118),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_88),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_83),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_70),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_121),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_84),
.A2(n_61),
.B1(n_60),
.B2(n_73),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_116),
.A2(n_84),
.B1(n_98),
.B2(n_96),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_80),
.A2(n_50),
.B1(n_65),
.B2(n_55),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_2),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_120),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_91),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_6),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_127),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_107),
.B(n_100),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_79),
.B(n_77),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_128),
.A2(n_131),
.B(n_133),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_112),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_132),
.Y(n_151)
);

AOI32xp33_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_85),
.A3(n_89),
.B1(n_102),
.B2(n_12),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_109),
.A2(n_89),
.B(n_99),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_82),
.C(n_99),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_142),
.C(n_104),
.Y(n_150)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_99),
.Y(n_138)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_124),
.A2(n_95),
.B1(n_5),
.B2(n_8),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_106),
.B1(n_104),
.B2(n_113),
.Y(n_149)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_5),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_114),
.Y(n_153)
);

NOR2xp67_ASAP7_75t_SL g145 ( 
.A(n_135),
.B(n_119),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_127),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_120),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_157),
.C(n_159),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_154),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_150),
.B(n_129),
.Y(n_169)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_134),
.A2(n_109),
.B1(n_113),
.B2(n_108),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_122),
.B(n_123),
.Y(n_155)
);

AOI22x1_ASAP7_75t_SL g166 ( 
.A1(n_155),
.A2(n_136),
.B1(n_139),
.B2(n_132),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_142),
.Y(n_156)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_123),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_122),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_153),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_160),
.B(n_165),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_150),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_149),
.A2(n_134),
.B1(n_136),
.B2(n_126),
.Y(n_165)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_137),
.C(n_141),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_169),
.Y(n_179)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_170),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_143),
.C(n_130),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_144),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_180),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_174),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_159),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_157),
.C(n_167),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_148),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_162),
.C(n_171),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_184),
.B(n_186),
.Y(n_188)
);

FAx1_ASAP7_75t_SL g185 ( 
.A(n_172),
.B(n_164),
.CI(n_165),
.CON(n_185),
.SN(n_185)
);

NOR3xp33_ASAP7_75t_SL g189 ( 
.A(n_185),
.B(n_173),
.C(n_151),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_176),
.Y(n_187)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_187),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_190),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_186),
.A2(n_178),
.B(n_179),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_179),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_191),
.B(n_184),
.Y(n_195)
);

BUFx24_ASAP7_75t_SL g192 ( 
.A(n_188),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_192),
.B(n_195),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_194),
.A2(n_167),
.B(n_183),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_196),
.A2(n_156),
.B(n_193),
.Y(n_199)
);

MAJx2_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_183),
.C(n_185),
.Y(n_198)
);

AOI322xp5_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_199),
.A3(n_166),
.B1(n_158),
.B2(n_155),
.C1(n_152),
.C2(n_154),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_7),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_14),
.Y(n_202)
);


endmodule