module fake_jpeg_23095_n_256 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_19),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_18),
.C(n_27),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_28),
.B1(n_27),
.B2(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_7),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_50),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_48),
.B1(n_23),
.B2(n_32),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_28),
.B1(n_18),
.B2(n_27),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_21),
.B1(n_31),
.B2(n_23),
.Y(n_62)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_31),
.C(n_21),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_57),
.B(n_66),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_68),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_62),
.A2(n_73),
.B1(n_26),
.B2(n_16),
.Y(n_101)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_64),
.Y(n_87)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_49),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_75),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_54),
.B(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_22),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

CKINVDCx10_ASAP7_75t_R g107 ( 
.A(n_70),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_22),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_74),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_24),
.B1(n_30),
.B2(n_19),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_22),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_25),
.Y(n_77)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_78),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_25),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_43),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_84),
.B1(n_29),
.B2(n_26),
.Y(n_93)
);

CKINVDCx12_ASAP7_75t_R g83 ( 
.A(n_43),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_83),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_52),
.A2(n_23),
.B1(n_21),
.B2(n_30),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_72),
.A2(n_52),
.B(n_44),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_85),
.A2(n_88),
.B(n_106),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_0),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_93),
.B(n_8),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_48),
.B1(n_45),
.B2(n_29),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_99),
.B1(n_64),
.B2(n_63),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_78),
.B1(n_71),
.B2(n_2),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_48),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_105),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_45),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_0),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_57),
.B(n_24),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_108),
.B(n_9),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_65),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_100),
.Y(n_128)
);

A2O1A1O1Ixp25_ASAP7_75t_L g110 ( 
.A1(n_99),
.A2(n_60),
.B(n_82),
.C(n_84),
.D(n_56),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_132),
.C(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_107),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_115),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_66),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_117),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_85),
.A2(n_62),
.B1(n_45),
.B2(n_58),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_149)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_108),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_116),
.B(n_120),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_70),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_109),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_118),
.Y(n_135)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_97),
.A2(n_58),
.B1(n_64),
.B2(n_81),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_96),
.A2(n_61),
.B1(n_70),
.B2(n_71),
.Y(n_122)
);

AOI221xp5_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_16),
.B1(n_70),
.B2(n_22),
.C(n_3),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_124),
.Y(n_145)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_126),
.Y(n_139)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_128),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_91),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_129),
.A2(n_98),
.B(n_103),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_102),
.B1(n_92),
.B2(n_90),
.Y(n_150)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_133),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_78),
.C(n_71),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_93),
.C(n_94),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_88),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_159),
.C(n_9),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_107),
.B(n_91),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_137),
.A2(n_148),
.B(n_157),
.Y(n_179)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_140),
.B(n_146),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_100),
.B(n_94),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_143),
.A2(n_151),
.B(n_160),
.Y(n_169)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_107),
.B(n_88),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_150),
.A2(n_154),
.B1(n_92),
.B2(n_4),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_113),
.A2(n_88),
.B(n_106),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_106),
.Y(n_153)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_114),
.A2(n_131),
.B1(n_120),
.B2(n_130),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_121),
.A2(n_101),
.B1(n_90),
.B2(n_106),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_111),
.B1(n_102),
.B2(n_92),
.Y(n_171)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_158),
.B(n_161),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_103),
.C(n_98),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_118),
.A2(n_0),
.B(n_1),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_147),
.B(n_134),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_165),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_147),
.B(n_126),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_143),
.B(n_132),
.Y(n_166)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_139),
.B(n_129),
.Y(n_168)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_168),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_133),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_152),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_171),
.A2(n_154),
.B1(n_146),
.B2(n_142),
.Y(n_194)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_173),
.Y(n_196)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_175),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_102),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_176),
.A2(n_181),
.B1(n_155),
.B2(n_153),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_157),
.Y(n_177)
);

INVxp33_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_151),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_139),
.B(n_9),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_180),
.A2(n_145),
.B1(n_142),
.B2(n_144),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_1),
.Y(n_181)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_137),
.A2(n_11),
.B(n_5),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_182),
.A2(n_145),
.B1(n_138),
.B2(n_140),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_183),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_11),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_152),
.C(n_144),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_187),
.A2(n_190),
.B1(n_173),
.B2(n_172),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_200),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_174),
.A2(n_158),
.B1(n_149),
.B2(n_141),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_193),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_192),
.A2(n_194),
.B1(n_176),
.B2(n_179),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_195),
.B(n_168),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_152),
.C(n_159),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_178),
.C(n_164),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_159),
.Y(n_200)
);

XOR2x1_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_169),
.Y(n_202)
);

XNOR2x1_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_205),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_208),
.C(n_212),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_209),
.Y(n_221)
);

XOR2x2_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_179),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_196),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_207),
.B(n_160),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_166),
.C(n_167),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_201),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_198),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_211),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_167),
.C(n_162),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_194),
.A2(n_163),
.B1(n_149),
.B2(n_183),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_213),
.A2(n_216),
.B1(n_202),
.B2(n_214),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_148),
.C(n_169),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_193),
.C(n_200),
.Y(n_223)
);

FAx1_ASAP7_75t_SL g217 ( 
.A(n_208),
.B(n_181),
.CI(n_199),
.CON(n_217),
.SN(n_217)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_217),
.B(n_227),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_205),
.A2(n_165),
.B(n_188),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_219),
.A2(n_8),
.B(n_5),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_224),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_192),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_188),
.C(n_180),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_12),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_226),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_220),
.A2(n_212),
.B1(n_203),
.B2(n_206),
.Y(n_228)
);

OAI21x1_ASAP7_75t_SL g242 ( 
.A1(n_228),
.A2(n_230),
.B(n_222),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_234),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_12),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_235),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_224),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_12),
.Y(n_235)
);

INVxp67_ASAP7_75t_SL g237 ( 
.A(n_230),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_237),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_220),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_241),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_217),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_229),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_234),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_238),
.B(n_222),
.Y(n_245)
);

AOI322xp5_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_246),
.A3(n_248),
.B1(n_7),
.B2(n_8),
.C1(n_13),
.C2(n_14),
.Y(n_251)
);

OAI221xp5_ASAP7_75t_L g249 ( 
.A1(n_247),
.A2(n_241),
.B1(n_240),
.B2(n_218),
.C(n_229),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_249),
.A2(n_251),
.B(n_15),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_218),
.C(n_6),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_250),
.A2(n_13),
.B(n_15),
.Y(n_252)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_252),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_254),
.A2(n_253),
.B(n_1),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_1),
.Y(n_256)
);


endmodule