module fake_ibex_1934_n_891 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_891);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_891;

wire n_599;
wire n_822;
wire n_778;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_270;
wire n_170;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_281;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_769;
wire n_487;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_433;
wire n_262;
wire n_439;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_837;
wire n_797;
wire n_796;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_392;
wire n_206;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_444;
wire n_200;
wire n_506;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_520;
wire n_411;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_499;
wire n_227;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_379;
wire n_288;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_440;
wire n_268;
wire n_858;
wire n_385;
wire n_233;
wire n_414;
wire n_342;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g168 ( 
.A(n_11),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_36),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_25),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_149),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_112),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_62),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_37),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_47),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_66),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_16),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_81),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_54),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_35),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_131),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_122),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_35),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_65),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_79),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_163),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_152),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_119),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_28),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_41),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_109),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_77),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_103),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_55),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_92),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_124),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_141),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_120),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_86),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_100),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_127),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_58),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_96),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_110),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_144),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_60),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_7),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_2),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_73),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_84),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_158),
.Y(n_214)
);

BUFx2_ASAP7_75t_SL g215 ( 
.A(n_140),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_25),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_102),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_64),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_20),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_72),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_133),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_51),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_167),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g225 ( 
.A(n_0),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_76),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_74),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_61),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_59),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_31),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_139),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_69),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_142),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_12),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_91),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_150),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_26),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_106),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_128),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_147),
.B(n_115),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_107),
.B(n_45),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_134),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_83),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_8),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_166),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_154),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_37),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_143),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_87),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_78),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_159),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_121),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_88),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_63),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_5),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_36),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_126),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_44),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_7),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_21),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_4),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_118),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_148),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_20),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_95),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_53),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_98),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_68),
.Y(n_268)
);

XNOR2x1_ASAP7_75t_L g269 ( 
.A(n_113),
.B(n_43),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_123),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_9),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_104),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_105),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_132),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_49),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_156),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_39),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_16),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_34),
.B(n_138),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_93),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_75),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_89),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_111),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_108),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_57),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_239),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_179),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_260),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_288)
);

OA21x2_ASAP7_75t_L g289 ( 
.A1(n_179),
.A2(n_94),
.B(n_165),
.Y(n_289)
);

BUFx12f_ASAP7_75t_L g290 ( 
.A(n_267),
.Y(n_290)
);

BUFx8_ASAP7_75t_SL g291 ( 
.A(n_181),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_230),
.Y(n_292)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_242),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_192),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_250),
.B(n_1),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_192),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_255),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_211),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_187),
.A2(n_3),
.B1(n_6),
.B2(n_8),
.Y(n_299)
);

OA21x2_ASAP7_75t_L g300 ( 
.A1(n_254),
.A2(n_97),
.B(n_164),
.Y(n_300)
);

CKINVDCx6p67_ASAP7_75t_R g301 ( 
.A(n_267),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_255),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_278),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_211),
.Y(n_304)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_267),
.Y(n_305)
);

AND2x6_ASAP7_75t_L g306 ( 
.A(n_239),
.B(n_46),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_173),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_254),
.Y(n_308)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_283),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_175),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_280),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_178),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_280),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_243),
.Y(n_314)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_183),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_193),
.Y(n_317)
);

AND2x4_ASAP7_75t_L g318 ( 
.A(n_243),
.B(n_168),
.Y(n_318)
);

AND2x4_ASAP7_75t_L g319 ( 
.A(n_169),
.B(n_6),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_195),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_197),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_283),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_201),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_247),
.Y(n_324)
);

BUFx12f_ASAP7_75t_L g325 ( 
.A(n_225),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_278),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_247),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_225),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_247),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g330 ( 
.A(n_174),
.B(n_10),
.Y(n_330)
);

AND2x4_ASAP7_75t_L g331 ( 
.A(n_191),
.B(n_10),
.Y(n_331)
);

OAI22x1_ASAP7_75t_L g332 ( 
.A1(n_210),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_247),
.Y(n_333)
);

BUFx12f_ASAP7_75t_L g334 ( 
.A(n_225),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_202),
.Y(n_335)
);

OA21x2_ASAP7_75t_L g336 ( 
.A1(n_204),
.A2(n_99),
.B(n_160),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_170),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_285),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_208),
.Y(n_339)
);

AND2x4_ASAP7_75t_L g340 ( 
.A(n_220),
.B(n_237),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_212),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_213),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_244),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_269),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_214),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_216),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_219),
.Y(n_347)
);

BUFx8_ASAP7_75t_SL g348 ( 
.A(n_181),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_221),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_223),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_224),
.Y(n_351)
);

OA21x2_ASAP7_75t_L g352 ( 
.A1(n_226),
.A2(n_101),
.B(n_157),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_228),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_229),
.B(n_15),
.Y(n_354)
);

OAI22x1_ASAP7_75t_SL g355 ( 
.A1(n_234),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_231),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_269),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_232),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_256),
.Y(n_359)
);

INVxp33_ASAP7_75t_SL g360 ( 
.A(n_176),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_338),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_286),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_338),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_338),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_315),
.B(n_293),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_293),
.B(n_176),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_293),
.B(n_180),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_315),
.B(n_180),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_326),
.A2(n_303),
.B1(n_360),
.B2(n_301),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_338),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_305),
.B(n_182),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_338),
.Y(n_372)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_306),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_315),
.B(n_182),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_286),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_286),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_301),
.B(n_185),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_286),
.Y(n_378)
);

NAND2xp33_ASAP7_75t_L g379 ( 
.A(n_306),
.B(n_240),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_286),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_337),
.B(n_177),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_289),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_305),
.B(n_185),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_324),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_322),
.B(n_186),
.Y(n_385)
);

XNOR2x2_ASAP7_75t_SL g386 ( 
.A(n_357),
.B(n_234),
.Y(n_386)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_306),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g388 ( 
.A(n_305),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_322),
.B(n_186),
.Y(n_389)
);

NAND3xp33_ASAP7_75t_L g390 ( 
.A(n_295),
.B(n_217),
.C(n_190),
.Y(n_390)
);

NAND2xp33_ASAP7_75t_L g391 ( 
.A(n_306),
.B(n_241),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_331),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_331),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_360),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_327),
.Y(n_395)
);

NAND2xp33_ASAP7_75t_L g396 ( 
.A(n_306),
.B(n_222),
.Y(n_396)
);

BUFx10_ASAP7_75t_L g397 ( 
.A(n_328),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_345),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_327),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_345),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_289),
.Y(n_401)
);

AOI21x1_ASAP7_75t_L g402 ( 
.A1(n_336),
.A2(n_238),
.B(n_233),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_345),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_305),
.B(n_222),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_345),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_305),
.B(n_273),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_345),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_309),
.B(n_273),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_309),
.B(n_276),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_309),
.B(n_276),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_350),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_350),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_350),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_298),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_350),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_351),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_351),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_289),
.Y(n_418)
);

INVx2_ASAP7_75t_SL g419 ( 
.A(n_318),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_290),
.B(n_172),
.Y(n_420)
);

NOR2x1p5_ASAP7_75t_L g421 ( 
.A(n_325),
.B(n_264),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_318),
.B(n_259),
.Y(n_422)
);

AND2x2_ASAP7_75t_SL g423 ( 
.A(n_319),
.B(n_330),
.Y(n_423)
);

NAND2xp33_ASAP7_75t_SL g424 ( 
.A(n_332),
.B(n_171),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_340),
.B(n_277),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_325),
.B(n_188),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_351),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_329),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_334),
.B(n_189),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_329),
.Y(n_430)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_298),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_318),
.B(n_261),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_306),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_319),
.Y(n_434)
);

NAND3xp33_ASAP7_75t_L g435 ( 
.A(n_319),
.B(n_271),
.C(n_279),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_333),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_333),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_333),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_291),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_343),
.B(n_184),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_287),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_287),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_343),
.B(n_215),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_314),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_299),
.A2(n_171),
.B1(n_196),
.B2(n_253),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_314),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_294),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_294),
.Y(n_448)
);

NAND3xp33_ASAP7_75t_L g449 ( 
.A(n_330),
.B(n_246),
.C(n_245),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_334),
.B(n_194),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_296),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_296),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_348),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_308),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_365),
.B(n_339),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_443),
.B(n_339),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_433),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_373),
.B(n_330),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_443),
.B(n_318),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_414),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_366),
.B(n_367),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_368),
.B(n_307),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_374),
.B(n_307),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_406),
.B(n_310),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_419),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_414),
.Y(n_466)
);

NAND3xp33_ASAP7_75t_L g467 ( 
.A(n_379),
.B(n_344),
.C(n_354),
.Y(n_467)
);

AND2x6_ASAP7_75t_L g468 ( 
.A(n_433),
.B(n_248),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_406),
.B(n_410),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_394),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_377),
.B(n_359),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_377),
.B(n_359),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_385),
.B(n_312),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_389),
.B(n_316),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_422),
.B(n_316),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_373),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_432),
.B(n_317),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_440),
.B(n_320),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_431),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_423),
.A2(n_196),
.B1(n_253),
.B2(n_270),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_423),
.B(n_320),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_441),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_441),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_425),
.B(n_346),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_387),
.B(n_346),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_425),
.B(n_347),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_387),
.B(n_347),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_434),
.B(n_349),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_392),
.A2(n_358),
.B1(n_353),
.B2(n_321),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_397),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_442),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_393),
.B(n_382),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_435),
.A2(n_274),
.B1(n_270),
.B2(n_288),
.Y(n_493)
);

O2A1O1Ixp5_ASAP7_75t_L g494 ( 
.A1(n_371),
.A2(n_358),
.B(n_353),
.C(n_342),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_379),
.A2(n_391),
.B1(n_396),
.B2(n_442),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_369),
.A2(n_356),
.B1(n_341),
.B2(n_321),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_449),
.B(n_323),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_382),
.B(n_249),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_382),
.B(n_251),
.Y(n_499)
);

NOR2x1p5_ASAP7_75t_L g500 ( 
.A(n_453),
.B(n_355),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_447),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_448),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_382),
.B(n_258),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_381),
.B(n_356),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_397),
.B(n_335),
.Y(n_505)
);

INVx4_ASAP7_75t_L g506 ( 
.A(n_397),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_391),
.A2(n_342),
.B1(n_306),
.B2(n_355),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_401),
.B(n_262),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_447),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_451),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_454),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_388),
.B(n_304),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_451),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_381),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_421),
.B(n_304),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_454),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_452),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_444),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_401),
.B(n_263),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_390),
.B(n_292),
.Y(n_520)
);

BUFx6f_ASAP7_75t_SL g521 ( 
.A(n_439),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_446),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_445),
.B(n_439),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_446),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_383),
.B(n_297),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_405),
.Y(n_526)
);

NOR3xp33_ASAP7_75t_L g527 ( 
.A(n_424),
.B(n_302),
.C(n_275),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_401),
.B(n_198),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_361),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_404),
.B(n_302),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_408),
.B(n_199),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_407),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_361),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_409),
.B(n_200),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_418),
.B(n_402),
.Y(n_535)
);

NAND2x1p5_ASAP7_75t_L g536 ( 
.A(n_420),
.B(n_289),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_386),
.A2(n_332),
.B1(n_336),
.B2(n_352),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_407),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_535),
.A2(n_492),
.B(n_498),
.Y(n_539)
);

AND2x2_ASAP7_75t_SL g540 ( 
.A(n_480),
.B(n_300),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_514),
.B(n_426),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_470),
.B(n_429),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_535),
.A2(n_402),
.B(n_352),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_507),
.A2(n_450),
.B1(n_418),
.B2(n_203),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_498),
.A2(n_418),
.B(n_300),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_499),
.A2(n_418),
.B(n_300),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_524),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_504),
.B(n_308),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_490),
.Y(n_549)
);

A2O1A1Ixp33_ASAP7_75t_L g550 ( 
.A1(n_475),
.A2(n_313),
.B(n_311),
.C(n_398),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_499),
.A2(n_352),
.B(n_336),
.Y(n_551)
);

A2O1A1Ixp33_ASAP7_75t_L g552 ( 
.A1(n_475),
.A2(n_313),
.B(n_311),
.C(n_398),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_495),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_479),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_490),
.B(n_209),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_506),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_478),
.B(n_266),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_L g558 ( 
.A1(n_469),
.A2(n_352),
.B(n_336),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_506),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_495),
.A2(n_218),
.B1(n_227),
.B2(n_235),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_457),
.B(n_236),
.Y(n_561)
);

AOI33xp33_ASAP7_75t_L g562 ( 
.A1(n_515),
.A2(n_400),
.A3(n_363),
.B1(n_364),
.B2(n_370),
.B3(n_372),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_476),
.B(n_252),
.Y(n_563)
);

NOR2xp67_ASAP7_75t_L g564 ( 
.A(n_493),
.B(n_22),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_481),
.B(n_471),
.Y(n_565)
);

O2A1O1Ixp33_ASAP7_75t_L g566 ( 
.A1(n_459),
.A2(n_438),
.B(n_437),
.C(n_436),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_503),
.A2(n_372),
.B(n_370),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_472),
.B(n_257),
.Y(n_568)
);

OAI321xp33_ASAP7_75t_L g569 ( 
.A1(n_537),
.A2(n_378),
.A3(n_362),
.B1(n_375),
.B2(n_376),
.C(n_380),
.Y(n_569)
);

A2O1A1Ixp33_ASAP7_75t_L g570 ( 
.A1(n_520),
.A2(n_403),
.B(n_412),
.C(n_415),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_489),
.A2(n_467),
.B1(n_474),
.B2(n_473),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_484),
.B(n_265),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_456),
.B(n_268),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_464),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_486),
.B(n_272),
.Y(n_575)
);

NOR3xp33_ASAP7_75t_L g576 ( 
.A(n_527),
.B(n_281),
.C(n_282),
.Y(n_576)
);

OAI321xp33_ASAP7_75t_L g577 ( 
.A1(n_496),
.A2(n_380),
.A3(n_362),
.B1(n_375),
.B2(n_376),
.C(n_378),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_508),
.A2(n_519),
.B(n_458),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_477),
.B(n_284),
.Y(n_579)
);

OAI21xp33_ASAP7_75t_L g580 ( 
.A1(n_462),
.A2(n_438),
.B(n_437),
.Y(n_580)
);

OAI21xp33_ASAP7_75t_L g581 ( 
.A1(n_463),
.A2(n_436),
.B(n_430),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_505),
.B(n_23),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_461),
.B(n_24),
.Y(n_583)
);

A2O1A1Ixp33_ASAP7_75t_L g584 ( 
.A1(n_520),
.A2(n_411),
.B(n_413),
.C(n_427),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_488),
.B(n_27),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_518),
.B(n_27),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_518),
.B(n_28),
.Y(n_587)
);

A2O1A1Ixp33_ASAP7_75t_L g588 ( 
.A1(n_482),
.A2(n_417),
.B(n_416),
.C(n_428),
.Y(n_588)
);

AO21x1_ASAP7_75t_L g589 ( 
.A1(n_536),
.A2(n_399),
.B(n_395),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_509),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_476),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_522),
.B(n_29),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_513),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_465),
.A2(n_384),
.B1(n_30),
.B2(n_31),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_485),
.A2(n_114),
.B(n_155),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_483),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_531),
.B(n_33),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_491),
.B(n_33),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_502),
.Y(n_599)
);

AO21x1_ASAP7_75t_L g600 ( 
.A1(n_528),
.A2(n_34),
.B(n_38),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_485),
.A2(n_487),
.B(n_455),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_511),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_497),
.A2(n_48),
.B1(n_50),
.B2(n_52),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_534),
.B(n_56),
.Y(n_604)
);

BUFx4f_ASAP7_75t_L g605 ( 
.A(n_468),
.Y(n_605)
);

OA22x2_ASAP7_75t_L g606 ( 
.A1(n_500),
.A2(n_67),
.B1(n_70),
.B2(n_71),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_516),
.B(n_517),
.Y(n_607)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_468),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_501),
.B(n_510),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_512),
.A2(n_80),
.B(n_82),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_466),
.A2(n_85),
.B(n_90),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_521),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_460),
.Y(n_613)
);

NAND3xp33_ASAP7_75t_SL g614 ( 
.A(n_494),
.B(n_525),
.C(n_530),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_468),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_L g616 ( 
.A1(n_558),
.A2(n_533),
.B(n_529),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_559),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_565),
.B(n_538),
.Y(n_618)
);

AOI21xp33_ASAP7_75t_L g619 ( 
.A1(n_542),
.A2(n_532),
.B(n_526),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_541),
.B(n_117),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_599),
.B(n_557),
.Y(n_621)
);

AOI211x1_ASAP7_75t_L g622 ( 
.A1(n_600),
.A2(n_125),
.B(n_129),
.C(n_130),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_612),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_548),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_607),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_549),
.Y(n_626)
);

AND3x2_ASAP7_75t_L g627 ( 
.A(n_615),
.B(n_145),
.C(n_146),
.Y(n_627)
);

OAI21x1_ASAP7_75t_L g628 ( 
.A1(n_546),
.A2(n_543),
.B(n_589),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_572),
.B(n_151),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_605),
.A2(n_540),
.B1(n_586),
.B2(n_587),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_575),
.B(n_564),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_579),
.B(n_556),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_556),
.B(n_568),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_598),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_592),
.A2(n_544),
.B1(n_582),
.B2(n_585),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_576),
.B(n_573),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_601),
.A2(n_567),
.B(n_609),
.Y(n_637)
);

NAND3x1_ASAP7_75t_L g638 ( 
.A(n_606),
.B(n_603),
.C(n_562),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_596),
.Y(n_639)
);

A2O1A1Ixp33_ASAP7_75t_L g640 ( 
.A1(n_566),
.A2(n_552),
.B(n_550),
.C(n_604),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_L g641 ( 
.A1(n_570),
.A2(n_584),
.B(n_614),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_602),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_594),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_593),
.B(n_547),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_591),
.Y(n_645)
);

AO31x2_ASAP7_75t_L g646 ( 
.A1(n_588),
.A2(n_610),
.A3(n_611),
.B(n_595),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_590),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_577),
.A2(n_580),
.B(n_581),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_606),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_553),
.B(n_560),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_555),
.B(n_563),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_561),
.Y(n_652)
);

OAI21xp5_ASAP7_75t_L g653 ( 
.A1(n_577),
.A2(n_613),
.B(n_569),
.Y(n_653)
);

A2O1A1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_569),
.A2(n_583),
.B(n_597),
.C(n_475),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_574),
.B(n_514),
.Y(n_655)
);

INVx5_ASAP7_75t_L g656 ( 
.A(n_559),
.Y(n_656)
);

BUFx5_ASAP7_75t_L g657 ( 
.A(n_593),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_591),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_545),
.A2(n_535),
.B(n_546),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_559),
.B(n_574),
.Y(n_660)
);

INVx5_ASAP7_75t_L g661 ( 
.A(n_559),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_574),
.B(n_514),
.Y(n_662)
);

OR2x6_ASAP7_75t_L g663 ( 
.A(n_559),
.B(n_608),
.Y(n_663)
);

BUFx12f_ASAP7_75t_L g664 ( 
.A(n_559),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_554),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_559),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_574),
.B(n_514),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_559),
.Y(n_668)
);

AOI21xp33_ASAP7_75t_L g669 ( 
.A1(n_542),
.A2(n_470),
.B(n_394),
.Y(n_669)
);

OR2x6_ASAP7_75t_L g670 ( 
.A(n_559),
.B(n_608),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_574),
.B(n_514),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_574),
.B(n_514),
.Y(n_672)
);

BUFx4f_ASAP7_75t_SL g673 ( 
.A(n_559),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_558),
.A2(n_539),
.B(n_578),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_559),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_574),
.B(n_514),
.Y(n_676)
);

CKINVDCx6p67_ASAP7_75t_R g677 ( 
.A(n_612),
.Y(n_677)
);

A2O1A1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_583),
.A2(n_597),
.B(n_475),
.C(n_571),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_L g679 ( 
.A1(n_558),
.A2(n_539),
.B(n_578),
.Y(n_679)
);

A2O1A1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_583),
.A2(n_597),
.B(n_475),
.C(n_571),
.Y(n_680)
);

NAND2x1p5_ASAP7_75t_L g681 ( 
.A(n_559),
.B(n_549),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_554),
.Y(n_682)
);

CKINVDCx6p67_ASAP7_75t_R g683 ( 
.A(n_612),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_574),
.B(n_514),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_612),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_574),
.B(n_514),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_574),
.B(n_514),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_574),
.B(n_514),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_574),
.B(n_514),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_554),
.Y(n_690)
);

A2O1A1Ixp33_ASAP7_75t_L g691 ( 
.A1(n_583),
.A2(n_597),
.B(n_475),
.C(n_571),
.Y(n_691)
);

O2A1O1Ixp33_ASAP7_75t_L g692 ( 
.A1(n_571),
.A2(n_514),
.B(n_583),
.C(n_585),
.Y(n_692)
);

AO31x2_ASAP7_75t_L g693 ( 
.A1(n_589),
.A2(n_600),
.A3(n_551),
.B(n_552),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_554),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_667),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_656),
.B(n_661),
.Y(n_696)
);

OR2x6_ASAP7_75t_L g697 ( 
.A(n_664),
.B(n_663),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_682),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_686),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_665),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_649),
.A2(n_642),
.B1(n_639),
.B2(n_643),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_660),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_673),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_624),
.A2(n_630),
.B1(n_654),
.B2(n_638),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_617),
.Y(n_705)
);

OA21x2_ASAP7_75t_L g706 ( 
.A1(n_628),
.A2(n_679),
.B(n_674),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_692),
.A2(n_621),
.B1(n_635),
.B2(n_634),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_650),
.A2(n_631),
.B1(n_690),
.B2(n_694),
.Y(n_708)
);

OR2x6_ASAP7_75t_L g709 ( 
.A(n_663),
.B(n_670),
.Y(n_709)
);

OAI21xp5_ASAP7_75t_L g710 ( 
.A1(n_637),
.A2(n_641),
.B(n_616),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_636),
.A2(n_684),
.B1(n_662),
.B2(n_672),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_655),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_671),
.B(n_676),
.Y(n_713)
);

OAI21xp5_ASAP7_75t_L g714 ( 
.A1(n_616),
.A2(n_640),
.B(n_618),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_687),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_623),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_688),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_663),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_656),
.B(n_661),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_689),
.A2(n_620),
.B1(n_632),
.B2(n_633),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_661),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_668),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_670),
.B(n_666),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_675),
.B(n_626),
.Y(n_724)
);

INVx5_ASAP7_75t_L g725 ( 
.A(n_670),
.Y(n_725)
);

NAND3xp33_ASAP7_75t_L g726 ( 
.A(n_622),
.B(n_669),
.C(n_651),
.Y(n_726)
);

BUFx10_ASAP7_75t_L g727 ( 
.A(n_652),
.Y(n_727)
);

AOI221xp5_ASAP7_75t_L g728 ( 
.A1(n_685),
.A2(n_619),
.B1(n_647),
.B2(n_629),
.C(n_625),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_644),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_681),
.Y(n_730)
);

AOI222xp33_ASAP7_75t_L g731 ( 
.A1(n_626),
.A2(n_658),
.B1(n_645),
.B2(n_683),
.C1(n_677),
.C2(n_627),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_657),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_646),
.B(n_693),
.Y(n_733)
);

OAI21xp5_ASAP7_75t_L g734 ( 
.A1(n_678),
.A2(n_691),
.B(n_680),
.Y(n_734)
);

AOI221xp5_ASAP7_75t_L g735 ( 
.A1(n_639),
.A2(n_344),
.B1(n_514),
.B2(n_424),
.C(n_571),
.Y(n_735)
);

OAI21xp5_ASAP7_75t_L g736 ( 
.A1(n_678),
.A2(n_691),
.B(n_680),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_667),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_673),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_649),
.A2(n_537),
.B1(n_642),
.B2(n_639),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_667),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_SL g741 ( 
.A1(n_649),
.A2(n_606),
.B1(n_523),
.B2(n_234),
.Y(n_741)
);

INVx6_ASAP7_75t_L g742 ( 
.A(n_656),
.Y(n_742)
);

AO21x2_ASAP7_75t_L g743 ( 
.A1(n_648),
.A2(n_653),
.B(n_659),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_684),
.B(n_514),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_660),
.B(n_656),
.Y(n_745)
);

NAND2x1p5_ASAP7_75t_L g746 ( 
.A(n_656),
.B(n_661),
.Y(n_746)
);

NAND2x1_ASAP7_75t_L g747 ( 
.A(n_663),
.B(n_670),
.Y(n_747)
);

AOI21xp33_ASAP7_75t_L g748 ( 
.A1(n_692),
.A2(n_649),
.B(n_630),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_667),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_649),
.A2(n_680),
.B1(n_691),
.B2(n_678),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_649),
.A2(n_680),
.B1(n_691),
.B2(n_678),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_705),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_712),
.B(n_715),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_701),
.B(n_739),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_746),
.Y(n_755)
);

NAND2x1p5_ASAP7_75t_L g756 ( 
.A(n_725),
.B(n_747),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_700),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_746),
.Y(n_758)
);

NAND2x1p5_ASAP7_75t_L g759 ( 
.A(n_725),
.B(n_719),
.Y(n_759)
);

OR2x2_ASAP7_75t_L g760 ( 
.A(n_713),
.B(n_701),
.Y(n_760)
);

AND2x4_ASAP7_75t_SL g761 ( 
.A(n_709),
.B(n_745),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_750),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_719),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_717),
.B(n_744),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_751),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_751),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_739),
.B(n_698),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_706),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_695),
.B(n_699),
.Y(n_769)
);

INVxp33_ASAP7_75t_L g770 ( 
.A(n_696),
.Y(n_770)
);

CKINVDCx11_ASAP7_75t_R g771 ( 
.A(n_727),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_706),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_741),
.B(n_731),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_708),
.B(n_702),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_722),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_741),
.B(n_731),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_742),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_737),
.B(n_740),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_709),
.B(n_725),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_732),
.Y(n_780)
);

AO21x2_ASAP7_75t_L g781 ( 
.A1(n_734),
.A2(n_736),
.B(n_710),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_735),
.A2(n_707),
.B1(n_711),
.B2(n_708),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_725),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_736),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_735),
.A2(n_707),
.B1(n_748),
.B2(n_726),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_714),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_749),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_733),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_720),
.B(n_729),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_781),
.B(n_743),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_781),
.B(n_704),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_771),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_781),
.B(n_704),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_773),
.B(n_723),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_776),
.A2(n_720),
.B1(n_697),
.B2(n_728),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_756),
.B(n_723),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_788),
.Y(n_797)
);

CKINVDCx6p67_ASAP7_75t_R g798 ( 
.A(n_763),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_780),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_784),
.B(n_786),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_760),
.B(n_774),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_760),
.B(n_721),
.Y(n_802)
);

OR2x2_ASAP7_75t_L g803 ( 
.A(n_774),
.B(n_718),
.Y(n_803)
);

OR2x2_ASAP7_75t_L g804 ( 
.A(n_762),
.B(n_697),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_756),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_790),
.B(n_768),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_800),
.B(n_754),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_800),
.B(n_754),
.Y(n_808)
);

OAI21xp5_ASAP7_75t_SL g809 ( 
.A1(n_795),
.A2(n_756),
.B(n_761),
.Y(n_809)
);

OAI222xp33_ASAP7_75t_L g810 ( 
.A1(n_795),
.A2(n_804),
.B1(n_782),
.B2(n_799),
.C1(n_805),
.C2(n_802),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_801),
.B(n_765),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_791),
.B(n_772),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_801),
.B(n_766),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_791),
.B(n_772),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_791),
.B(n_767),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_797),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_799),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_816),
.Y(n_818)
);

AND2x2_ASAP7_75t_SL g819 ( 
.A(n_817),
.B(n_761),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_807),
.B(n_789),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_812),
.B(n_790),
.Y(n_821)
);

OR2x2_ASAP7_75t_L g822 ( 
.A(n_811),
.B(n_801),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_817),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_811),
.B(n_803),
.Y(n_824)
);

NAND2xp33_ASAP7_75t_R g825 ( 
.A(n_806),
.B(n_792),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_807),
.B(n_789),
.Y(n_826)
);

OR2x2_ASAP7_75t_L g827 ( 
.A(n_813),
.B(n_803),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_814),
.B(n_793),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_814),
.B(n_793),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_828),
.B(n_815),
.Y(n_830)
);

OAI21xp5_ASAP7_75t_SL g831 ( 
.A1(n_825),
.A2(n_809),
.B(n_810),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_828),
.B(n_808),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_829),
.B(n_815),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_818),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_819),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_822),
.Y(n_836)
);

CKINVDCx16_ASAP7_75t_R g837 ( 
.A(n_822),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_823),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_834),
.Y(n_839)
);

OR2x2_ASAP7_75t_L g840 ( 
.A(n_837),
.B(n_821),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_831),
.A2(n_809),
.B1(n_819),
.B2(n_798),
.Y(n_841)
);

NOR2xp67_ASAP7_75t_SL g842 ( 
.A(n_835),
.B(n_783),
.Y(n_842)
);

O2A1O1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_835),
.A2(n_810),
.B(n_752),
.C(n_697),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_838),
.A2(n_819),
.B(n_796),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_836),
.A2(n_794),
.B(n_761),
.C(n_805),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_832),
.A2(n_798),
.B1(n_805),
.B2(n_824),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_834),
.Y(n_847)
);

OAI22xp33_ASAP7_75t_L g848 ( 
.A1(n_830),
.A2(n_798),
.B1(n_827),
.B2(n_824),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_830),
.B(n_829),
.Y(n_849)
);

INVx1_ASAP7_75t_SL g850 ( 
.A(n_833),
.Y(n_850)
);

OAI22xp33_ASAP7_75t_L g851 ( 
.A1(n_841),
.A2(n_827),
.B1(n_826),
.B2(n_820),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_839),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_847),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_850),
.B(n_833),
.Y(n_854)
);

INVx1_ASAP7_75t_SL g855 ( 
.A(n_840),
.Y(n_855)
);

NAND2xp67_ASAP7_75t_SL g856 ( 
.A(n_851),
.B(n_842),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_855),
.B(n_849),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_853),
.B(n_848),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_858),
.A2(n_857),
.B(n_843),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_856),
.Y(n_860)
);

NOR3xp33_ASAP7_75t_L g861 ( 
.A(n_860),
.B(n_716),
.C(n_703),
.Y(n_861)
);

AND4x2_ASAP7_75t_L g862 ( 
.A(n_859),
.B(n_844),
.C(n_843),
.D(n_728),
.Y(n_862)
);

NOR2x1_ASAP7_75t_L g863 ( 
.A(n_862),
.B(n_852),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_861),
.B(n_852),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_863),
.B(n_854),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_864),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_866),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_865),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_866),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_869),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_869),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_867),
.B(n_846),
.Y(n_872)
);

AOI31xp33_ASAP7_75t_L g873 ( 
.A1(n_868),
.A2(n_738),
.A3(n_727),
.B(n_764),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_869),
.A2(n_845),
.B(n_794),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_871),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_870),
.B(n_769),
.Y(n_876)
);

INVx1_ASAP7_75t_SL g877 ( 
.A(n_872),
.Y(n_877)
);

OAI21xp5_ASAP7_75t_L g878 ( 
.A1(n_873),
.A2(n_770),
.B(n_777),
.Y(n_878)
);

OR4x1_ASAP7_75t_L g879 ( 
.A(n_874),
.B(n_730),
.C(n_777),
.D(n_757),
.Y(n_879)
);

OAI22x1_ASAP7_75t_L g880 ( 
.A1(n_871),
.A2(n_775),
.B1(n_778),
.B2(n_787),
.Y(n_880)
);

OAI21xp5_ASAP7_75t_SL g881 ( 
.A1(n_873),
.A2(n_759),
.B(n_779),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_877),
.A2(n_758),
.B(n_755),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_875),
.A2(n_804),
.B1(n_785),
.B2(n_742),
.Y(n_883)
);

AOI21x1_ASAP7_75t_L g884 ( 
.A1(n_876),
.A2(n_753),
.B(n_724),
.Y(n_884)
);

OAI21xp33_ASAP7_75t_L g885 ( 
.A1(n_878),
.A2(n_881),
.B(n_880),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_885),
.B(n_884),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_882),
.Y(n_887)
);

OAI221xp5_ASAP7_75t_L g888 ( 
.A1(n_883),
.A2(n_879),
.B1(n_742),
.B2(n_759),
.C(n_783),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_886),
.A2(n_779),
.B(n_759),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_889),
.B(n_887),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_890),
.A2(n_888),
.B(n_779),
.Y(n_891)
);


endmodule