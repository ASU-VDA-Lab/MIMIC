module fake_jpeg_22475_n_178 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

AOI21xp33_ASAP7_75t_L g26 ( 
.A1(n_5),
.A2(n_2),
.B(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_27),
.Y(n_50)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_16),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_SL g37 ( 
.A1(n_34),
.A2(n_26),
.B(n_25),
.Y(n_37)
);

NAND2x1p5_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_26),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_38),
.B(n_13),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_43),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_28),
.A2(n_21),
.B1(n_19),
.B2(n_18),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_21),
.B1(n_28),
.B2(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_29),
.B(n_20),
.Y(n_43)
);

CKINVDCx12_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_46),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_47),
.Y(n_54)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_33),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_45),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_55),
.B(n_57),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_28),
.B1(n_21),
.B2(n_18),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_44),
.B1(n_50),
.B2(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_62),
.Y(n_71)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_43),
.Y(n_70)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_65),
.Y(n_83)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_25),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_75),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_70),
.B(n_49),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_72),
.A2(n_73),
.B1(n_78),
.B2(n_50),
.Y(n_98)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_82),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_63),
.A2(n_34),
.B1(n_46),
.B2(n_52),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_63),
.A2(n_33),
.B1(n_30),
.B2(n_51),
.Y(n_79)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_57),
.A2(n_13),
.B1(n_48),
.B2(n_44),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_55),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_81),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_82),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_78),
.C(n_54),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_93),
.C(n_96),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_71),
.B(n_59),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_86),
.B(n_49),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_83),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_89),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_77),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_62),
.C(n_61),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_59),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_95),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_66),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_60),
.B1(n_74),
.B2(n_75),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_67),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_74),
.Y(n_107)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_107),
.Y(n_119)
);

NOR3xp33_ASAP7_75t_SL g105 ( 
.A(n_84),
.B(n_45),
.C(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_106),
.Y(n_125)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_68),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_111),
.A2(n_113),
.B1(n_98),
.B2(n_97),
.Y(n_122)
);

OAI22x1_ASAP7_75t_SL g113 ( 
.A1(n_95),
.A2(n_72),
.B1(n_73),
.B2(n_52),
.Y(n_113)
);

BUFx24_ASAP7_75t_SL g123 ( 
.A(n_114),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_93),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_118),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_96),
.C(n_85),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_101),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_100),
.B(n_102),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_122),
.A2(n_95),
.B1(n_111),
.B2(n_104),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_92),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_105),
.Y(n_133)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_127),
.Y(n_141)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_92),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_72),
.Y(n_140)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_135),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_137),
.B(n_125),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_121),
.B1(n_115),
.B2(n_112),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_140),
.C(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_118),
.B(n_108),
.Y(n_136)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_123),
.C(n_60),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_106),
.Y(n_138)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_116),
.B(n_103),
.Y(n_139)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_146),
.C(n_149),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_65),
.B(n_40),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_31),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_76),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_30),
.C(n_53),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_140),
.C(n_136),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_141),
.A2(n_65),
.B1(n_53),
.B2(n_15),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_14),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_152),
.B(n_151),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_155),
.C(n_159),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_134),
.C(n_24),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_158),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_147),
.B(n_143),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_23),
.C(n_15),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_166),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_162),
.A2(n_164),
.B(n_3),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_149),
.A3(n_23),
.B1(n_12),
.B2(n_11),
.C1(n_22),
.C2(n_25),
.Y(n_163)
);

OAI21x1_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_22),
.B(n_4),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_157),
.A2(n_12),
.B(n_4),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_31),
.C(n_27),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_167),
.B(n_160),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_169),
.B(n_3),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_165),
.A2(n_3),
.B(n_5),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_163),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_170),
.A2(n_5),
.B(n_6),
.Y(n_174)
);

AOI322xp5_ASAP7_75t_L g176 ( 
.A1(n_172),
.A2(n_173),
.A3(n_174),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_27),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_174),
.A2(n_171),
.B(n_27),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_176),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_31),
.Y(n_178)
);


endmodule