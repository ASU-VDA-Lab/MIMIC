module fake_jpeg_4725_n_177 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx6_ASAP7_75t_SL g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_34),
.Y(n_52)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_22),
.Y(n_34)
);

NOR3xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_1),
.C(n_2),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_37),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_36),
.Y(n_46)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_17),
.B1(n_27),
.B2(n_25),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_40),
.A2(n_32),
.B1(n_19),
.B2(n_23),
.Y(n_68)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_30),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_22),
.Y(n_64)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_33),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_27),
.B1(n_25),
.B2(n_17),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_26),
.B1(n_29),
.B2(n_21),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_68),
.B1(n_15),
.B2(n_20),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_24),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_58),
.Y(n_76)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_61),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_48),
.B1(n_37),
.B2(n_45),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_24),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_38),
.C(n_32),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_19),
.Y(n_85)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_71),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_38),
.B1(n_33),
.B2(n_32),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_66),
.A2(n_47),
.B1(n_50),
.B2(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_41),
.B(n_29),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_23),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_70),
.B(n_39),
.Y(n_88)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_24),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_23),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_38),
.B(n_24),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_38),
.B(n_47),
.C(n_20),
.Y(n_82)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_16),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_80),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_90),
.B(n_73),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_20),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_93),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_19),
.B1(n_15),
.B2(n_20),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_89),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_66),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_87),
.B(n_88),
.Y(n_100)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_1),
.B(n_2),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_39),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_60),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_59),
.B(n_8),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_12),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_1),
.Y(n_93)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_75),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_96),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_86),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_97),
.B(n_101),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_108),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_106),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_93),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_110),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_68),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_85),
.C(n_83),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_111),
.C(n_113),
.Y(n_116)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_79),
.A2(n_66),
.B(n_55),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_79),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_91),
.C(n_94),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_129),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_119),
.A2(n_128),
.B(n_98),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_94),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_123),
.Y(n_138)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

XOR2x1_ASAP7_75t_SL g124 ( 
.A(n_101),
.B(n_89),
.Y(n_124)
);

NAND4xp25_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_126),
.C(n_98),
.D(n_129),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_77),
.Y(n_128)
);

A2O1A1O1Ixp25_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_77),
.B(n_81),
.C(n_61),
.D(n_16),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_105),
.B1(n_110),
.B2(n_114),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_131),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_127),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_137),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_139),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_115),
.A2(n_103),
.B1(n_113),
.B2(n_99),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_136),
.B(n_140),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_125),
.A2(n_98),
.B1(n_99),
.B2(n_74),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_128),
.B1(n_16),
.B2(n_56),
.Y(n_153)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_143),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_148),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_138),
.Y(n_148)
);

AOI322xp5_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_128),
.A3(n_116),
.B1(n_118),
.B2(n_117),
.C1(n_120),
.C2(n_56),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_151),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_116),
.Y(n_151)
);

AOI31xp67_ASAP7_75t_L g160 ( 
.A1(n_153),
.A2(n_16),
.A3(n_69),
.B(n_6),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_145),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_158),
.Y(n_161)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_143),
.B(n_137),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_152),
.Y(n_165)
);

OAI31xp33_ASAP7_75t_L g166 ( 
.A1(n_160),
.A2(n_153),
.A3(n_5),
.B(n_6),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_147),
.Y(n_162)
);

OAI221xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_164),
.B1(n_9),
.B2(n_13),
.C(n_69),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_154),
.B(n_150),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_165),
.A2(n_134),
.B1(n_5),
.B2(n_4),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_166),
.A2(n_4),
.B1(n_9),
.B2(n_13),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_161),
.A2(n_159),
.B1(n_134),
.B2(n_151),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_169),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_170),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_168),
.A2(n_163),
.B(n_166),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_165),
.Y(n_175)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_173),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_174),
.A2(n_175),
.B(n_172),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_4),
.Y(n_177)
);


endmodule