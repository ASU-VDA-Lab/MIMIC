module fake_jpeg_31771_n_164 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_28),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_29),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_8),
.B(n_7),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_5),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_0),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_0),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_75),
.Y(n_88)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_90),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_46),
.B1(n_56),
.B2(n_60),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_80),
.A2(n_83),
.B1(n_73),
.B2(n_55),
.Y(n_92)
);

CKINVDCx12_ASAP7_75t_R g82 ( 
.A(n_72),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_82),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_75),
.A2(n_46),
.B1(n_60),
.B2(n_61),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_76),
.Y(n_85)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_100),
.Y(n_111)
);

NOR2x1_ASAP7_75t_R g96 ( 
.A(n_88),
.B(n_71),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_79),
.B(n_58),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_97),
.B(n_99),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_65),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_102),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_66),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_51),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_101),
.B(n_107),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_85),
.B(n_48),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_66),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_104),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_53),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_74),
.B1(n_50),
.B2(n_64),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_84),
.B(n_67),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_64),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_18),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_63),
.B1(n_47),
.B2(n_62),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_110),
.A2(n_119),
.B1(n_124),
.B2(n_12),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_115),
.B(n_120),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_52),
.B1(n_66),
.B2(n_44),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_38),
.B1(n_17),
.B2(n_20),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_117),
.A2(n_125),
.B1(n_92),
.B2(n_119),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_121),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_94),
.B(n_1),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_6),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_93),
.A2(n_34),
.B1(n_21),
.B2(n_23),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_25),
.B1(n_31),
.B2(n_30),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_127),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_112),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_130),
.B(n_132),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_135),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_13),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_140),
.C(n_133),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_14),
.B(n_15),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_117),
.A2(n_16),
.B1(n_26),
.B2(n_27),
.Y(n_137)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_32),
.B(n_122),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_109),
.C(n_123),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_134),
.C(n_136),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_142),
.A2(n_140),
.B1(n_141),
.B2(n_131),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_149),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_129),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_154),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_150),
.C(n_149),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_138),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_151),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_155),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_143),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_146),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_144),
.Y(n_163)
);

BUFx24_ASAP7_75t_SL g164 ( 
.A(n_163),
.Y(n_164)
);


endmodule