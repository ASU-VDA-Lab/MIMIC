module fake_aes_12008_n_909 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_909);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_909;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_903;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_228;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_167;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_171;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_529;
wire n_455;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_769;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_818;
wire n_844;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_711;
wire n_238;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_699;
wire n_338;
wire n_519;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_649;
wire n_526;
wire n_276;
wire n_527;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_420;
wire n_621;
wire n_666;
wire n_342;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_200;
wire n_208;
wire n_573;
wire n_898;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_899;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g110 ( .A(n_76), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_61), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_17), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_21), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_18), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_42), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_23), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_5), .Y(n_117) );
BUFx10_ASAP7_75t_L g118 ( .A(n_77), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_3), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_22), .Y(n_120) );
INVxp67_ASAP7_75t_L g121 ( .A(n_53), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_79), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_17), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_99), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_72), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_28), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_25), .Y(n_127) );
BUFx3_ASAP7_75t_L g128 ( .A(n_6), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_46), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_29), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_60), .Y(n_131) );
INVxp67_ASAP7_75t_L g132 ( .A(n_57), .Y(n_132) );
BUFx3_ASAP7_75t_L g133 ( .A(n_62), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_47), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_59), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_56), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_63), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_40), .Y(n_138) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_2), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_91), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_98), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_71), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_49), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_30), .Y(n_144) );
BUFx3_ASAP7_75t_L g145 ( .A(n_103), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_50), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_27), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_19), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_85), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_94), .Y(n_150) );
INVxp67_ASAP7_75t_SL g151 ( .A(n_11), .Y(n_151) );
NOR2xp67_ASAP7_75t_L g152 ( .A(n_78), .B(n_34), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_139), .B(n_0), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_118), .B(n_0), .Y(n_154) );
OAI22xp5_ASAP7_75t_SL g155 ( .A1(n_112), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_128), .Y(n_156) );
CKINVDCx6p67_ASAP7_75t_R g157 ( .A(n_118), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_125), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_125), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_128), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_118), .Y(n_161) );
INVx5_ASAP7_75t_L g162 ( .A(n_125), .Y(n_162) );
NOR2x1_ASAP7_75t_L g163 ( .A(n_119), .B(n_20), .Y(n_163) );
AND2x6_ASAP7_75t_L g164 ( .A(n_133), .B(n_24), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_125), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_111), .Y(n_166) );
AND2x6_ASAP7_75t_L g167 ( .A(n_133), .B(n_26), .Y(n_167) );
NAND2xp33_ASAP7_75t_L g168 ( .A(n_113), .B(n_109), .Y(n_168) );
AND2x2_ASAP7_75t_SL g169 ( .A(n_115), .B(n_31), .Y(n_169) );
BUFx8_ASAP7_75t_L g170 ( .A(n_110), .Y(n_170) );
NAND2xp33_ASAP7_75t_L g171 ( .A(n_113), .B(n_108), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_112), .Y(n_172) );
BUFx3_ASAP7_75t_L g173 ( .A(n_145), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_120), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_122), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_166), .B(n_110), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_156), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_161), .B(n_116), .Y(n_178) );
BUFx10_ASAP7_75t_L g179 ( .A(n_164), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_161), .B(n_116), .Y(n_180) );
NAND2xp33_ASAP7_75t_R g181 ( .A(n_172), .B(n_114), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_161), .B(n_127), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_173), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_169), .A2(n_114), .B1(n_117), .B2(n_148), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_166), .B(n_129), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_157), .B(n_117), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_162), .Y(n_187) );
AND2x6_ASAP7_75t_L g188 ( .A(n_153), .B(n_145), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_158), .Y(n_189) );
INVxp67_ASAP7_75t_L g190 ( .A(n_172), .Y(n_190) );
OAI22xp33_ASAP7_75t_L g191 ( .A1(n_157), .A2(n_151), .B1(n_123), .B2(n_141), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_174), .B(n_129), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_162), .Y(n_193) );
INVx6_ASAP7_75t_L g194 ( .A(n_170), .Y(n_194) );
BUFx4f_ASAP7_75t_L g195 ( .A(n_164), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_162), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_162), .Y(n_197) );
NOR2x1p5_ASAP7_75t_L g198 ( .A(n_153), .B(n_127), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_174), .B(n_121), .Y(n_199) );
INVx2_ASAP7_75t_SL g200 ( .A(n_170), .Y(n_200) );
INVxp67_ASAP7_75t_L g201 ( .A(n_173), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_156), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_170), .B(n_130), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_162), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_158), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_162), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_158), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_160), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_160), .Y(n_209) );
CKINVDCx6p67_ASAP7_75t_R g210 ( .A(n_169), .Y(n_210) );
INVx3_ASAP7_75t_L g211 ( .A(n_175), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_158), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_158), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_175), .B(n_130), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_159), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_159), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_159), .Y(n_217) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_154), .A2(n_124), .B(n_150), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_163), .B(n_132), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_159), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_200), .B(n_136), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_183), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_211), .B(n_201), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_178), .B(n_168), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_211), .Y(n_225) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_181), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_211), .B(n_136), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_177), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_177), .Y(n_229) );
NOR2xp67_ASAP7_75t_L g230 ( .A(n_200), .B(n_32), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_186), .B(n_138), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_199), .B(n_138), .Y(n_232) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_186), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_195), .B(n_141), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_202), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_202), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_214), .B(n_144), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_188), .B(n_144), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_188), .B(n_147), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_188), .B(n_147), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_180), .B(n_171), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_188), .B(n_149), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_208), .Y(n_243) );
NOR3xp33_ASAP7_75t_L g244 ( .A(n_191), .B(n_155), .C(n_126), .Y(n_244) );
BUFx3_ASAP7_75t_L g245 ( .A(n_194), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_194), .B(n_149), .Y(n_246) );
BUFx3_ASAP7_75t_L g247 ( .A(n_194), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g248 ( .A1(n_176), .A2(n_142), .B(n_134), .C(n_135), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_188), .B(n_164), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_188), .B(n_164), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_188), .B(n_164), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_182), .B(n_137), .Y(n_252) );
NAND2xp33_ASAP7_75t_L g253 ( .A(n_198), .B(n_164), .Y(n_253) );
NAND3xp33_ASAP7_75t_SL g254 ( .A(n_184), .B(n_143), .C(n_146), .Y(n_254) );
INVx2_ASAP7_75t_SL g255 ( .A(n_194), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_208), .Y(n_256) );
INVx4_ASAP7_75t_L g257 ( .A(n_179), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_209), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_219), .B(n_164), .Y(n_259) );
INVx2_ASAP7_75t_SL g260 ( .A(n_179), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_209), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_183), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_195), .B(n_131), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_183), .Y(n_264) );
OAI22xp33_ASAP7_75t_L g265 ( .A1(n_210), .A2(n_184), .B1(n_190), .B2(n_192), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_195), .B(n_131), .Y(n_266) );
BUFx3_ASAP7_75t_L g267 ( .A(n_179), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_176), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_210), .A2(n_167), .B1(n_146), .B2(n_140), .Y(n_269) );
AOI22xp33_ASAP7_75t_SL g270 ( .A1(n_218), .A2(n_167), .B1(n_140), .B2(n_125), .Y(n_270) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_198), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_185), .B(n_167), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_185), .B(n_167), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_189), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_192), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_179), .B(n_167), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_203), .B(n_167), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_218), .B(n_167), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_218), .B(n_152), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_272), .A2(n_206), .B(n_193), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_245), .B(n_187), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_233), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_268), .B(n_187), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_268), .Y(n_284) );
NAND2xp33_ASAP7_75t_L g285 ( .A(n_275), .B(n_193), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_275), .A2(n_206), .B1(n_196), .B2(n_197), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_231), .B(n_196), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_231), .B(n_197), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_229), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_229), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_273), .A2(n_204), .B(n_216), .Y(n_291) );
NAND2x1_ASAP7_75t_L g292 ( .A(n_235), .B(n_204), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_246), .B(n_1), .Y(n_293) );
NOR3xp33_ASAP7_75t_L g294 ( .A(n_265), .B(n_217), .C(n_216), .Y(n_294) );
OAI21xp5_ASAP7_75t_L g295 ( .A1(n_278), .A2(n_207), .B(n_212), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_246), .B(n_4), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_235), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_259), .A2(n_207), .B(n_212), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_254), .A2(n_159), .B1(n_165), .B2(n_217), .Y(n_299) );
OAI21xp33_ASAP7_75t_L g300 ( .A1(n_232), .A2(n_217), .B(n_165), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_236), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_225), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_225), .Y(n_303) );
NOR2xp67_ASAP7_75t_L g304 ( .A(n_271), .B(n_4), .Y(n_304) );
BUFx2_ASAP7_75t_L g305 ( .A(n_226), .Y(n_305) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_245), .Y(n_306) );
A2O1A1Ixp33_ASAP7_75t_L g307 ( .A1(n_236), .A2(n_165), .B(n_189), .C(n_220), .Y(n_307) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_245), .B(n_165), .Y(n_308) );
BUFx2_ASAP7_75t_L g309 ( .A(n_227), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_244), .A2(n_165), .B1(n_189), .B2(n_220), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_225), .Y(n_311) );
OR2x6_ASAP7_75t_SL g312 ( .A(n_238), .B(n_5), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_228), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_228), .B(n_6), .Y(n_314) );
OAI21xp5_ASAP7_75t_L g315 ( .A1(n_243), .A2(n_215), .B(n_213), .Y(n_315) );
AO32x1_ASAP7_75t_L g316 ( .A1(n_262), .A2(n_220), .A3(n_215), .B1(n_213), .B2(n_205), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_223), .B(n_7), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_269), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_318) );
AO21x1_ASAP7_75t_L g319 ( .A1(n_279), .A2(n_8), .B(n_9), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_247), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g321 ( .A1(n_243), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_321) );
NOR3xp33_ASAP7_75t_L g322 ( .A(n_248), .B(n_10), .C(n_12), .Y(n_322) );
OAI22xp5_ASAP7_75t_SL g323 ( .A1(n_270), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_323) );
AO21x1_ASAP7_75t_L g324 ( .A1(n_253), .A2(n_13), .B(n_14), .Y(n_324) );
BUFx6f_ASAP7_75t_SL g325 ( .A(n_247), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_256), .A2(n_15), .B1(n_16), .B2(n_18), .Y(n_326) );
O2A1O1Ixp33_ASAP7_75t_L g327 ( .A1(n_256), .A2(n_16), .B(n_33), .C(n_35), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_258), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_285), .A2(n_277), .B(n_250), .Y(n_329) );
O2A1O1Ixp33_ASAP7_75t_SL g330 ( .A1(n_327), .A2(n_249), .B(n_251), .C(n_258), .Y(n_330) );
INVx1_ASAP7_75t_SL g331 ( .A(n_282), .Y(n_331) );
INVxp67_ASAP7_75t_SL g332 ( .A(n_284), .Y(n_332) );
AO31x2_ASAP7_75t_L g333 ( .A1(n_324), .A2(n_261), .A3(n_228), .B(n_264), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_325), .Y(n_334) );
OAI21xp33_ASAP7_75t_L g335 ( .A1(n_293), .A2(n_241), .B(n_224), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_309), .B(n_237), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_291), .A2(n_263), .B(n_266), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_313), .B(n_261), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_289), .B(n_252), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_287), .Y(n_340) );
INVxp67_ASAP7_75t_SL g341 ( .A(n_283), .Y(n_341) );
NOR2xp67_ASAP7_75t_SL g342 ( .A(n_320), .B(n_247), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_290), .B(n_261), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_288), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_305), .B(n_221), .Y(n_345) );
OAI21xp5_ASAP7_75t_L g346 ( .A1(n_291), .A2(n_276), .B(n_262), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_295), .A2(n_276), .B(n_262), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_314), .Y(n_348) );
AOI21xp5_ASAP7_75t_L g349 ( .A1(n_280), .A2(n_264), .B(n_234), .Y(n_349) );
AO31x2_ASAP7_75t_L g350 ( .A1(n_319), .A2(n_264), .A3(n_240), .B(n_239), .Y(n_350) );
BUFx3_ASAP7_75t_L g351 ( .A(n_320), .Y(n_351) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_320), .Y(n_352) );
OAI21x1_ASAP7_75t_L g353 ( .A1(n_298), .A2(n_230), .B(n_222), .Y(n_353) );
OAI21x1_ASAP7_75t_L g354 ( .A1(n_298), .A2(n_315), .B(n_280), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_312), .B(n_242), .Y(n_355) );
AOI21x1_ASAP7_75t_L g356 ( .A1(n_296), .A2(n_230), .B(n_274), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_325), .Y(n_357) );
OAI21x1_ASAP7_75t_L g358 ( .A1(n_327), .A2(n_222), .B(n_274), .Y(n_358) );
A2O1A1Ixp33_ASAP7_75t_L g359 ( .A1(n_297), .A2(n_222), .B(n_255), .C(n_267), .Y(n_359) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_341), .A2(n_316), .B(n_307), .Y(n_360) );
OA21x2_ASAP7_75t_L g361 ( .A1(n_358), .A2(n_300), .B(n_310), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_343), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_354), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_354), .Y(n_364) );
AO31x2_ASAP7_75t_L g365 ( .A1(n_359), .A2(n_301), .A3(n_328), .B(n_318), .Y(n_365) );
AO21x2_ASAP7_75t_L g366 ( .A1(n_358), .A2(n_322), .B(n_294), .Y(n_366) );
OA21x2_ASAP7_75t_L g367 ( .A1(n_353), .A2(n_310), .B(n_294), .Y(n_367) );
AOI21x1_ASAP7_75t_L g368 ( .A1(n_356), .A2(n_292), .B(n_316), .Y(n_368) );
NOR2xp67_ASAP7_75t_SL g369 ( .A(n_352), .B(n_320), .Y(n_369) );
AND2x4_ASAP7_75t_L g370 ( .A(n_351), .B(n_332), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_338), .Y(n_371) );
OAI21x1_ASAP7_75t_L g372 ( .A1(n_353), .A2(n_316), .B(n_317), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_343), .Y(n_373) );
AO21x2_ASAP7_75t_L g374 ( .A1(n_330), .A2(n_322), .B(n_326), .Y(n_374) );
INVx2_ASAP7_75t_SL g375 ( .A(n_351), .Y(n_375) );
AO31x2_ASAP7_75t_L g376 ( .A1(n_359), .A2(n_321), .A3(n_286), .B(n_311), .Y(n_376) );
OAI21x1_ASAP7_75t_L g377 ( .A1(n_349), .A2(n_299), .B(n_308), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_340), .Y(n_378) );
OA21x2_ASAP7_75t_L g379 ( .A1(n_347), .A2(n_303), .B(n_302), .Y(n_379) );
OAI21x1_ASAP7_75t_L g380 ( .A1(n_329), .A2(n_346), .B(n_337), .Y(n_380) );
BUFx2_ASAP7_75t_L g381 ( .A(n_352), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_338), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_352), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_334), .Y(n_384) );
OA21x2_ASAP7_75t_L g385 ( .A1(n_335), .A2(n_304), .B(n_281), .Y(n_385) );
OAI21x1_ASAP7_75t_L g386 ( .A1(n_348), .A2(n_222), .B(n_306), .Y(n_386) );
OAI21x1_ASAP7_75t_L g387 ( .A1(n_339), .A2(n_306), .B(n_274), .Y(n_387) );
OAI21xp5_ASAP7_75t_L g388 ( .A1(n_344), .A2(n_255), .B(n_260), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_378), .B(n_350), .Y(n_389) );
INVx2_ASAP7_75t_SL g390 ( .A(n_370), .Y(n_390) );
INVx3_ASAP7_75t_L g391 ( .A(n_383), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_362), .Y(n_392) );
HB1xp67_ASAP7_75t_SL g393 ( .A(n_370), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_363), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_362), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_363), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_363), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_387), .Y(n_398) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_387), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_378), .B(n_350), .Y(n_400) );
OAI21x1_ASAP7_75t_L g401 ( .A1(n_372), .A2(n_333), .B(n_355), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_364), .Y(n_402) );
INVx3_ASAP7_75t_L g403 ( .A(n_383), .Y(n_403) );
OA21x2_ASAP7_75t_L g404 ( .A1(n_372), .A2(n_333), .B(n_330), .Y(n_404) );
BUFx3_ASAP7_75t_L g405 ( .A(n_381), .Y(n_405) );
INVx3_ASAP7_75t_L g406 ( .A(n_383), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_364), .Y(n_407) );
BUFx2_ASAP7_75t_L g408 ( .A(n_387), .Y(n_408) );
OAI21x1_ASAP7_75t_L g409 ( .A1(n_372), .A2(n_333), .B(n_350), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_381), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_373), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_374), .B(n_350), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_381), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_373), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_376), .B(n_331), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_386), .Y(n_416) );
BUFx3_ASAP7_75t_L g417 ( .A(n_370), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_386), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_376), .B(n_333), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_364), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_376), .B(n_352), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_371), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_386), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_371), .Y(n_424) );
BUFx3_ASAP7_75t_L g425 ( .A(n_370), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_370), .Y(n_426) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_368), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_379), .Y(n_428) );
OA21x2_ASAP7_75t_L g429 ( .A1(n_380), .A2(n_336), .B(n_323), .Y(n_429) );
INVxp67_ASAP7_75t_SL g430 ( .A(n_379), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_376), .B(n_357), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_415), .B(n_376), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_431), .B(n_376), .Y(n_433) );
AND2x4_ASAP7_75t_L g434 ( .A(n_417), .B(n_425), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_431), .B(n_376), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_394), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_392), .Y(n_437) );
INVx5_ASAP7_75t_L g438 ( .A(n_393), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_394), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_431), .A2(n_429), .B1(n_415), .B2(n_400), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_392), .Y(n_441) );
INVxp33_ASAP7_75t_L g442 ( .A(n_393), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_389), .B(n_376), .Y(n_443) );
INVx2_ASAP7_75t_SL g444 ( .A(n_417), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_394), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_394), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_415), .B(n_365), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_426), .B(n_365), .Y(n_448) );
OAI221xp5_ASAP7_75t_L g449 ( .A1(n_429), .A2(n_345), .B1(n_334), .B2(n_384), .C(n_388), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_389), .B(n_366), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_429), .A2(n_374), .B1(n_366), .B2(n_367), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_389), .B(n_374), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_417), .B(n_384), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_417), .B(n_375), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_426), .B(n_365), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_400), .B(n_374), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_395), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_407), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_407), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_407), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_425), .B(n_371), .Y(n_461) );
BUFx3_ASAP7_75t_L g462 ( .A(n_405), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_400), .B(n_374), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_407), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_425), .B(n_365), .Y(n_465) );
AND2x4_ASAP7_75t_L g466 ( .A(n_425), .B(n_390), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_396), .Y(n_467) );
BUFx3_ASAP7_75t_L g468 ( .A(n_405), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_395), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_390), .B(n_365), .Y(n_470) );
INVxp67_ASAP7_75t_L g471 ( .A(n_410), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_421), .B(n_366), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_410), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_411), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_411), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_414), .Y(n_476) );
INVxp67_ASAP7_75t_L g477 ( .A(n_413), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_396), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_390), .B(n_365), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_414), .B(n_365), .Y(n_480) );
BUFx2_ASAP7_75t_L g481 ( .A(n_430), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_413), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_401), .B(n_365), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_421), .B(n_382), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_396), .Y(n_485) );
AND2x4_ASAP7_75t_L g486 ( .A(n_421), .B(n_382), .Y(n_486) );
NAND3xp33_ASAP7_75t_L g487 ( .A(n_412), .B(n_385), .C(n_360), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_419), .B(n_366), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_397), .Y(n_489) );
BUFx3_ASAP7_75t_L g490 ( .A(n_405), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_428), .Y(n_491) );
INVx8_ASAP7_75t_L g492 ( .A(n_391), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_428), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_397), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_397), .Y(n_495) );
INVx1_ASAP7_75t_SL g496 ( .A(n_405), .Y(n_496) );
BUFx3_ASAP7_75t_L g497 ( .A(n_391), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_419), .B(n_366), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_419), .B(n_382), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_429), .B(n_375), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_401), .B(n_367), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_391), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_429), .B(n_375), .Y(n_503) );
BUFx2_ASAP7_75t_L g504 ( .A(n_438), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_437), .Y(n_505) );
INVx2_ASAP7_75t_SL g506 ( .A(n_438), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_441), .B(n_429), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_473), .B(n_430), .Y(n_508) );
BUFx3_ASAP7_75t_L g509 ( .A(n_438), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_436), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_481), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_457), .Y(n_512) );
AND2x4_ASAP7_75t_SL g513 ( .A(n_434), .B(n_391), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_436), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_472), .B(n_401), .Y(n_515) );
INVx3_ASAP7_75t_L g516 ( .A(n_438), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_434), .B(n_391), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_472), .B(n_408), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_439), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_469), .B(n_412), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_471), .B(n_408), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_439), .Y(n_522) );
INVxp67_ASAP7_75t_SL g523 ( .A(n_481), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_474), .B(n_422), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_475), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_476), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_445), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_445), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_482), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_484), .B(n_408), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_450), .B(n_398), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_450), .B(n_398), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_477), .B(n_402), .Y(n_533) );
INVx1_ASAP7_75t_SL g534 ( .A(n_496), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_446), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_491), .Y(n_536) );
BUFx3_ASAP7_75t_L g537 ( .A(n_438), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_498), .B(n_399), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_498), .B(n_499), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_499), .B(n_399), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_493), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_462), .B(n_402), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_443), .B(n_416), .Y(n_543) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_497), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_443), .B(n_422), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_462), .B(n_402), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_467), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_446), .Y(n_548) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_458), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_458), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_433), .B(n_422), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_434), .B(n_403), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_466), .B(n_403), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_484), .B(n_416), .Y(n_554) );
INVx3_ASAP7_75t_L g555 ( .A(n_497), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_467), .Y(n_556) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_459), .Y(n_557) );
INVx3_ASAP7_75t_L g558 ( .A(n_492), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_478), .Y(n_559) );
INVxp67_ASAP7_75t_SL g560 ( .A(n_502), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_433), .B(n_424), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_478), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_435), .B(n_418), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_435), .B(n_418), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_485), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_466), .B(n_403), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_485), .Y(n_567) );
AND2x4_ASAP7_75t_SL g568 ( .A(n_466), .B(n_403), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_484), .B(n_423), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_488), .B(n_424), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_489), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_489), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_494), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_468), .B(n_420), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_468), .B(n_420), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_494), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_459), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_490), .B(n_420), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_460), .Y(n_579) );
BUFx2_ASAP7_75t_L g580 ( .A(n_490), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_444), .B(n_424), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_440), .B(n_403), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_486), .B(n_423), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_449), .B(n_453), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_495), .Y(n_585) );
BUFx2_ASAP7_75t_L g586 ( .A(n_492), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_495), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_486), .B(n_409), .Y(n_588) );
AND2x4_ASAP7_75t_L g589 ( .A(n_486), .B(n_409), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_452), .B(n_406), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_460), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_464), .Y(n_592) );
INVx2_ASAP7_75t_SL g593 ( .A(n_492), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_456), .B(n_406), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_444), .B(n_406), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_465), .B(n_409), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_464), .Y(n_597) );
INVxp67_ASAP7_75t_SL g598 ( .A(n_442), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_465), .Y(n_599) );
AND2x4_ASAP7_75t_L g600 ( .A(n_461), .B(n_406), .Y(n_600) );
BUFx3_ASAP7_75t_L g601 ( .A(n_492), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_501), .B(n_404), .Y(n_602) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_461), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_539), .B(n_448), .Y(n_604) );
AND2x4_ASAP7_75t_L g605 ( .A(n_580), .B(n_461), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_599), .B(n_480), .Y(n_606) );
AND2x4_ASAP7_75t_L g607 ( .A(n_523), .B(n_448), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_529), .Y(n_608) );
BUFx2_ASAP7_75t_L g609 ( .A(n_586), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_539), .B(n_442), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_543), .B(n_563), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_543), .B(n_480), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_563), .B(n_454), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_564), .B(n_455), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_564), .B(n_455), .Y(n_615) );
AND2x4_ASAP7_75t_L g616 ( .A(n_589), .B(n_470), .Y(n_616) );
OAI32xp33_ASAP7_75t_L g617 ( .A1(n_511), .A2(n_447), .A3(n_432), .B1(n_483), .B2(n_470), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_538), .B(n_479), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_505), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_512), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_525), .Y(n_621) );
AND2x4_ASAP7_75t_SL g622 ( .A(n_558), .B(n_406), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_536), .B(n_463), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_510), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_526), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_538), .B(n_479), .Y(n_626) );
NAND2x1_ASAP7_75t_SL g627 ( .A(n_516), .B(n_501), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_518), .B(n_500), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_518), .B(n_503), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_531), .B(n_447), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_541), .Y(n_631) );
INVx1_ASAP7_75t_SL g632 ( .A(n_534), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_549), .Y(n_633) );
BUFx2_ASAP7_75t_L g634 ( .A(n_601), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_508), .Y(n_635) );
NAND2x1p5_ASAP7_75t_L g636 ( .A(n_601), .B(n_369), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_531), .B(n_432), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_532), .B(n_483), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_524), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_515), .B(n_451), .Y(n_640) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_511), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_532), .B(n_404), .Y(n_642) );
OAI21xp33_ASAP7_75t_L g643 ( .A1(n_584), .A2(n_487), .B(n_427), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_517), .B(n_404), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_533), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_552), .B(n_553), .Y(n_646) );
OR2x2_ASAP7_75t_L g647 ( .A(n_551), .B(n_404), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_566), .B(n_404), .Y(n_648) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_549), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_557), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_561), .B(n_404), .Y(n_651) );
INVxp67_ASAP7_75t_L g652 ( .A(n_557), .Y(n_652) );
INVx3_ASAP7_75t_L g653 ( .A(n_516), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_515), .B(n_427), .Y(n_654) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_542), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_520), .B(n_427), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_507), .B(n_427), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_540), .B(n_427), .Y(n_658) );
INVxp67_ASAP7_75t_L g659 ( .A(n_560), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_570), .B(n_427), .Y(n_660) );
AND2x4_ASAP7_75t_L g661 ( .A(n_589), .B(n_427), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_521), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_540), .B(n_427), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_590), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_594), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_510), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_569), .B(n_367), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_596), .B(n_367), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_547), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_514), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_596), .B(n_367), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_556), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_559), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_569), .B(n_379), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_545), .B(n_602), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_546), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_562), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_602), .B(n_591), .Y(n_678) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_574), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_592), .B(n_380), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_583), .B(n_379), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_583), .B(n_379), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_565), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_567), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_571), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_588), .B(n_380), .Y(n_686) );
NOR2x1_ASAP7_75t_L g687 ( .A(n_558), .B(n_360), .Y(n_687) );
OR2x2_ASAP7_75t_L g688 ( .A(n_575), .B(n_385), .Y(n_688) );
OR2x2_ASAP7_75t_L g689 ( .A(n_578), .B(n_385), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_514), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_519), .Y(n_691) );
AND2x2_ASAP7_75t_L g692 ( .A(n_588), .B(n_385), .Y(n_692) );
NAND2x1p5_ASAP7_75t_L g693 ( .A(n_558), .B(n_369), .Y(n_693) );
NOR2x1_ASAP7_75t_L g694 ( .A(n_516), .B(n_509), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_597), .B(n_361), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_519), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_572), .B(n_361), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_530), .B(n_385), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_530), .B(n_361), .Y(n_699) );
AND2x4_ASAP7_75t_L g700 ( .A(n_589), .B(n_368), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_530), .B(n_361), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_573), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_603), .B(n_361), .Y(n_703) );
INVx2_ASAP7_75t_SL g704 ( .A(n_593), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_576), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_603), .B(n_368), .Y(n_706) );
AOI211xp5_ASAP7_75t_SL g707 ( .A1(n_584), .A2(n_369), .B(n_37), .C(n_38), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_611), .B(n_598), .Y(n_708) );
AOI21xp33_ASAP7_75t_SL g709 ( .A1(n_704), .A2(n_593), .B(n_506), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_619), .Y(n_710) );
NAND2x1_ASAP7_75t_L g711 ( .A(n_694), .B(n_504), .Y(n_711) );
NOR2xp67_ASAP7_75t_L g712 ( .A(n_653), .B(n_506), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_646), .B(n_554), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_649), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_664), .B(n_585), .Y(n_715) );
OR2x2_ASAP7_75t_L g716 ( .A(n_675), .B(n_582), .Y(n_716) );
NOR2x1p5_ASAP7_75t_SL g717 ( .A(n_688), .B(n_522), .Y(n_717) );
BUFx2_ASAP7_75t_L g718 ( .A(n_627), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_620), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_610), .B(n_638), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_613), .B(n_554), .Y(n_721) );
AND2x4_ASAP7_75t_L g722 ( .A(n_616), .B(n_554), .Y(n_722) );
INVx1_ASAP7_75t_SL g723 ( .A(n_609), .Y(n_723) );
BUFx3_ASAP7_75t_L g724 ( .A(n_634), .Y(n_724) );
NAND2xp5_ASAP7_75t_SL g725 ( .A(n_653), .B(n_509), .Y(n_725) );
AND2x4_ASAP7_75t_L g726 ( .A(n_616), .B(n_555), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_621), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_615), .B(n_600), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_635), .B(n_587), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_649), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_665), .B(n_522), .Y(n_731) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_655), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_662), .B(n_527), .Y(n_733) );
INVx1_ASAP7_75t_SL g734 ( .A(n_655), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_625), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_637), .B(n_600), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_679), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_639), .B(n_527), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_640), .B(n_528), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_679), .Y(n_740) );
CKINVDCx16_ASAP7_75t_R g741 ( .A(n_632), .Y(n_741) );
INVx3_ASAP7_75t_L g742 ( .A(n_700), .Y(n_742) );
NOR3xp33_ASAP7_75t_L g743 ( .A(n_643), .B(n_555), .C(n_595), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_608), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_631), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_618), .B(n_600), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_640), .B(n_535), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_623), .B(n_535), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_678), .Y(n_749) );
OR2x6_ASAP7_75t_L g750 ( .A(n_693), .B(n_537), .Y(n_750) );
OR2x2_ASAP7_75t_L g751 ( .A(n_675), .B(n_581), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_678), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_645), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_669), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_672), .Y(n_755) );
INVx1_ASAP7_75t_SL g756 ( .A(n_641), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_673), .Y(n_757) );
OR2x2_ASAP7_75t_L g758 ( .A(n_604), .B(n_579), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_612), .B(n_579), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_626), .B(n_513), .Y(n_760) );
INVx2_ASAP7_75t_SL g761 ( .A(n_622), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_612), .B(n_544), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_677), .Y(n_763) );
OR2x2_ASAP7_75t_L g764 ( .A(n_614), .B(n_577), .Y(n_764) );
OR2x2_ASAP7_75t_L g765 ( .A(n_630), .B(n_577), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_683), .Y(n_766) );
INVx2_ASAP7_75t_SL g767 ( .A(n_622), .Y(n_767) );
OR2x2_ASAP7_75t_L g768 ( .A(n_676), .B(n_550), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_628), .B(n_513), .Y(n_769) );
NAND2xp5_ASAP7_75t_SL g770 ( .A(n_659), .B(n_537), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_684), .Y(n_771) );
A2O1A1Ixp33_ASAP7_75t_L g772 ( .A1(n_707), .A2(n_568), .B(n_555), .C(n_544), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_623), .B(n_550), .Y(n_773) );
OAI21xp33_ASAP7_75t_L g774 ( .A1(n_617), .A2(n_568), .B(n_548), .Y(n_774) );
OR2x2_ASAP7_75t_L g775 ( .A(n_606), .B(n_548), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_629), .B(n_544), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_685), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_606), .B(n_528), .Y(n_778) );
INVxp67_ASAP7_75t_L g779 ( .A(n_641), .Y(n_779) );
NAND2x1p5_ASAP7_75t_L g780 ( .A(n_605), .B(n_544), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_659), .B(n_650), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_702), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_605), .B(n_644), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_642), .B(n_377), .Y(n_784) );
INVx2_ASAP7_75t_L g785 ( .A(n_633), .Y(n_785) );
INVx2_ASAP7_75t_SL g786 ( .A(n_636), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_652), .B(n_377), .Y(n_787) );
NAND2x2_ASAP7_75t_L g788 ( .A(n_654), .B(n_36), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_705), .B(n_377), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_652), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_781), .Y(n_791) );
OAI22xp33_ASAP7_75t_L g792 ( .A1(n_788), .A2(n_707), .B1(n_693), .B2(n_636), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_741), .A2(n_607), .B1(n_654), .B2(n_671), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_732), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_774), .A2(n_686), .B1(n_700), .B2(n_661), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_749), .B(n_660), .Y(n_796) );
OR2x2_ASAP7_75t_L g797 ( .A(n_734), .B(n_647), .Y(n_797) );
O2A1O1Ixp33_ASAP7_75t_L g798 ( .A1(n_772), .A2(n_687), .B(n_660), .C(n_656), .Y(n_798) );
AOI22x1_ASAP7_75t_L g799 ( .A1(n_718), .A2(n_607), .B1(n_661), .B2(n_689), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_752), .B(n_656), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_790), .Y(n_801) );
OR2x2_ASAP7_75t_L g802 ( .A(n_734), .B(n_651), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_723), .B(n_648), .Y(n_803) );
OAI211xp5_ASAP7_75t_SL g804 ( .A1(n_774), .A2(n_657), .B(n_668), .C(n_671), .Y(n_804) );
OAI221xp5_ASAP7_75t_L g805 ( .A1(n_723), .A2(n_657), .B1(n_668), .B2(n_698), .C(n_680), .Y(n_805) );
AOI222xp33_ASAP7_75t_L g806 ( .A1(n_753), .A2(n_692), .B1(n_703), .B2(n_706), .C1(n_681), .C2(n_674), .Y(n_806) );
A2O1A1Ixp33_ASAP7_75t_L g807 ( .A1(n_709), .A2(n_682), .B(n_663), .C(n_658), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_783), .B(n_667), .Y(n_808) );
XOR2x2_ASAP7_75t_L g809 ( .A(n_724), .B(n_720), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_715), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_716), .B(n_690), .Y(n_811) );
OR2x2_ASAP7_75t_L g812 ( .A(n_765), .B(n_691), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_715), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_737), .B(n_690), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_739), .B(n_691), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_751), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_759), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_759), .Y(n_818) );
INVx2_ASAP7_75t_L g819 ( .A(n_756), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_710), .Y(n_820) );
INVxp67_ASAP7_75t_SL g821 ( .A(n_779), .Y(n_821) );
OAI21xp5_ASAP7_75t_L g822 ( .A1(n_709), .A2(n_680), .B(n_624), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_740), .B(n_624), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_719), .Y(n_824) );
AND2x2_ASAP7_75t_L g825 ( .A(n_721), .B(n_701), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_727), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_756), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_747), .B(n_696), .Y(n_828) );
AOI22xp5_ASAP7_75t_L g829 ( .A1(n_762), .A2(n_699), .B1(n_670), .B2(n_696), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_735), .Y(n_830) );
INVxp67_ASAP7_75t_L g831 ( .A(n_744), .Y(n_831) );
O2A1O1Ixp33_ASAP7_75t_SL g832 ( .A1(n_711), .A2(n_670), .B(n_666), .C(n_695), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_714), .Y(n_833) );
OAI221xp5_ASAP7_75t_L g834 ( .A1(n_743), .A2(n_666), .B1(n_695), .B2(n_697), .C(n_388), .Y(n_834) );
AND2x4_ASAP7_75t_L g835 ( .A(n_712), .B(n_697), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_786), .A2(n_342), .B1(n_205), .B2(n_43), .Y(n_836) );
INVx2_ASAP7_75t_L g837 ( .A(n_730), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_745), .Y(n_838) );
INVxp67_ASAP7_75t_SL g839 ( .A(n_712), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_722), .A2(n_205), .B1(n_41), .B2(n_44), .Y(n_840) );
OAI22xp5_ASAP7_75t_L g841 ( .A1(n_793), .A2(n_750), .B1(n_722), .B2(n_726), .Y(n_841) );
A2O1A1Ixp33_ASAP7_75t_L g842 ( .A1(n_839), .A2(n_717), .B(n_761), .C(n_767), .Y(n_842) );
AOI22xp5_ASAP7_75t_L g843 ( .A1(n_793), .A2(n_726), .B1(n_742), .B2(n_776), .Y(n_843) );
AOI21xp5_ASAP7_75t_L g844 ( .A1(n_832), .A2(n_770), .B(n_725), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_810), .B(n_708), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_813), .B(n_773), .Y(n_846) );
OAI21xp5_ASAP7_75t_SL g847 ( .A1(n_792), .A2(n_780), .B(n_742), .Y(n_847) );
AOI332xp33_ASAP7_75t_L g848 ( .A1(n_791), .A2(n_795), .A3(n_816), .B1(n_794), .B2(n_818), .B3(n_817), .C1(n_801), .C2(n_830), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_804), .A2(n_750), .B1(n_784), .B2(n_769), .Y(n_849) );
OAI321xp33_ASAP7_75t_L g850 ( .A1(n_834), .A2(n_750), .A3(n_733), .B1(n_773), .B2(n_738), .C(n_787), .Y(n_850) );
OAI21xp5_ASAP7_75t_L g851 ( .A1(n_798), .A2(n_729), .B(n_713), .Y(n_851) );
AOI21xp33_ASAP7_75t_L g852 ( .A1(n_821), .A2(n_763), .B(n_754), .Y(n_852) );
A2O1A1Ixp33_ASAP7_75t_L g853 ( .A1(n_807), .A2(n_760), .B(n_736), .C(n_728), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_811), .Y(n_854) );
AOI211xp5_ASAP7_75t_L g855 ( .A1(n_805), .A2(n_766), .B(n_755), .C(n_782), .Y(n_855) );
NOR2xp33_ASAP7_75t_L g856 ( .A(n_831), .B(n_771), .Y(n_856) );
INVx3_ASAP7_75t_L g857 ( .A(n_835), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_806), .B(n_777), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_796), .Y(n_859) );
OAI21xp5_ASAP7_75t_L g860 ( .A1(n_822), .A2(n_757), .B(n_748), .Y(n_860) );
AND2x2_ASAP7_75t_L g861 ( .A(n_825), .B(n_746), .Y(n_861) );
A2O1A1Ixp33_ASAP7_75t_L g862 ( .A1(n_822), .A2(n_758), .B(n_764), .C(n_775), .Y(n_862) );
AND4x1_ASAP7_75t_L g863 ( .A(n_806), .B(n_778), .C(n_731), .D(n_789), .Y(n_863) );
NOR2xp33_ASAP7_75t_L g864 ( .A(n_820), .B(n_768), .Y(n_864) );
NOR2xp33_ASAP7_75t_L g865 ( .A(n_824), .B(n_785), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_799), .A2(n_789), .B1(n_205), .B2(n_48), .Y(n_866) );
AOI221xp5_ASAP7_75t_L g867 ( .A1(n_826), .A2(n_205), .B1(n_45), .B2(n_51), .C(n_52), .Y(n_867) );
AOI221x1_ASAP7_75t_L g868 ( .A1(n_819), .A2(n_39), .B1(n_54), .B2(n_55), .C(n_58), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g869 ( .A(n_858), .B(n_838), .Y(n_869) );
AOI221xp5_ASAP7_75t_L g870 ( .A1(n_850), .A2(n_800), .B1(n_796), .B2(n_803), .C(n_835), .Y(n_870) );
O2A1O1Ixp33_ASAP7_75t_L g871 ( .A1(n_847), .A2(n_827), .B(n_800), .C(n_802), .Y(n_871) );
NAND4xp25_ASAP7_75t_L g872 ( .A(n_866), .B(n_840), .C(n_836), .D(n_829), .Y(n_872) );
OAI221xp5_ASAP7_75t_L g873 ( .A1(n_849), .A2(n_809), .B1(n_797), .B2(n_815), .C(n_828), .Y(n_873) );
OAI21xp33_ASAP7_75t_L g874 ( .A1(n_863), .A2(n_815), .B(n_823), .Y(n_874) );
OAI221xp5_ASAP7_75t_SL g875 ( .A1(n_843), .A2(n_812), .B1(n_814), .B2(n_808), .C(n_837), .Y(n_875) );
NOR2xp67_ASAP7_75t_L g876 ( .A(n_841), .B(n_844), .Y(n_876) );
OAI21xp5_ASAP7_75t_SL g877 ( .A1(n_842), .A2(n_833), .B(n_65), .Y(n_877) );
AOI221xp5_ASAP7_75t_L g878 ( .A1(n_855), .A2(n_64), .B1(n_66), .B2(n_67), .C(n_68), .Y(n_878) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_856), .B(n_852), .Y(n_879) );
OAI221xp5_ASAP7_75t_L g880 ( .A1(n_857), .A2(n_69), .B1(n_70), .B2(n_73), .C(n_74), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_854), .Y(n_881) );
AOI221xp5_ASAP7_75t_L g882 ( .A1(n_862), .A2(n_75), .B1(n_80), .B2(n_81), .C(n_82), .Y(n_882) );
OAI221xp5_ASAP7_75t_L g883 ( .A1(n_857), .A2(n_83), .B1(n_84), .B2(n_86), .C(n_87), .Y(n_883) );
AOI222xp33_ASAP7_75t_L g884 ( .A1(n_876), .A2(n_860), .B1(n_851), .B2(n_859), .C1(n_848), .C2(n_865), .Y(n_884) );
AOI22xp5_ASAP7_75t_L g885 ( .A1(n_879), .A2(n_864), .B1(n_853), .B2(n_845), .Y(n_885) );
NAND3xp33_ASAP7_75t_L g886 ( .A(n_871), .B(n_867), .C(n_868), .Y(n_886) );
AOI21xp5_ASAP7_75t_L g887 ( .A1(n_877), .A2(n_846), .B(n_867), .Y(n_887) );
AND4x1_ASAP7_75t_L g888 ( .A(n_878), .B(n_861), .C(n_89), .D(n_90), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_881), .Y(n_889) );
NOR2xp33_ASAP7_75t_SL g890 ( .A(n_880), .B(n_257), .Y(n_890) );
NOR4xp25_ASAP7_75t_L g891 ( .A(n_873), .B(n_88), .C(n_92), .D(n_93), .Y(n_891) );
NAND3xp33_ASAP7_75t_L g892 ( .A(n_884), .B(n_869), .C(n_882), .Y(n_892) );
NOR4xp75_ASAP7_75t_L g893 ( .A(n_891), .B(n_874), .C(n_883), .D(n_875), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_889), .Y(n_894) );
NOR2x1_ASAP7_75t_L g895 ( .A(n_886), .B(n_872), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_894), .Y(n_896) );
AND3x4_ASAP7_75t_L g897 ( .A(n_895), .B(n_888), .C(n_887), .Y(n_897) );
BUFx2_ASAP7_75t_L g898 ( .A(n_892), .Y(n_898) );
XNOR2x1_ASAP7_75t_L g899 ( .A(n_897), .B(n_893), .Y(n_899) );
INVx2_ASAP7_75t_L g900 ( .A(n_896), .Y(n_900) );
AOI311xp33_ASAP7_75t_L g901 ( .A1(n_899), .A2(n_898), .A3(n_870), .B(n_885), .C(n_890), .Y(n_901) );
XOR2xp5_ASAP7_75t_L g902 ( .A(n_900), .B(n_95), .Y(n_902) );
CKINVDCx20_ASAP7_75t_R g903 ( .A(n_902), .Y(n_903) );
OAI22xp5_ASAP7_75t_L g904 ( .A1(n_901), .A2(n_257), .B1(n_267), .B2(n_260), .Y(n_904) );
OAI22xp33_ASAP7_75t_L g905 ( .A1(n_903), .A2(n_257), .B1(n_267), .B2(n_100), .Y(n_905) );
OR2x6_ASAP7_75t_L g906 ( .A(n_905), .B(n_904), .Y(n_906) );
AOI222xp33_ASAP7_75t_L g907 ( .A1(n_906), .A2(n_96), .B1(n_97), .B2(n_101), .C1(n_102), .C2(n_104), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_907), .B(n_105), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_908), .A2(n_257), .B1(n_106), .B2(n_107), .Y(n_909) );
endmodule