module fake_jpeg_1594_n_466 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_466);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_466;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_47),
.B(n_53),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_48),
.Y(n_152)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g119 ( 
.A(n_51),
.Y(n_119)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_52),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_16),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx11_ASAP7_75t_SL g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_55),
.Y(n_126)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_56),
.B(n_59),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_57),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_26),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_60),
.B(n_61),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_26),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_21),
.B(n_12),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_64),
.B(n_85),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_66),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_69),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_38),
.A2(n_12),
.B(n_11),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g135 ( 
.A(n_72),
.B(n_89),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_46),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_73),
.B(n_78),
.Y(n_139)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_74),
.B(n_87),
.Y(n_148)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_18),
.B(n_12),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_79),
.Y(n_155)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_14),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_81),
.Y(n_118)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_14),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_17),
.Y(n_84)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_21),
.B(n_10),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_14),
.Y(n_86)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_35),
.B(n_10),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_88),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

BUFx10_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g154 ( 
.A1(n_90),
.A2(n_23),
.B(n_24),
.Y(n_154)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_17),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_91),
.B(n_92),
.Y(n_151)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_93),
.B(n_94),
.Y(n_150)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_95),
.B(n_96),
.Y(n_156)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_20),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_97),
.B(n_98),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_26),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_37),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_18),
.B1(n_27),
.B2(n_32),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_101),
.A2(n_137),
.B1(n_144),
.B2(n_15),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_29),
.B1(n_37),
.B2(n_32),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_103),
.B(n_115),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_86),
.A2(n_30),
.B1(n_28),
.B2(n_31),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_108),
.A2(n_109),
.B1(n_120),
.B2(n_136),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_76),
.A2(n_30),
.B1(n_28),
.B2(n_31),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_63),
.A2(n_37),
.B1(n_29),
.B2(n_32),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_110),
.A2(n_117),
.B1(n_134),
.B2(n_93),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_82),
.A2(n_99),
.B1(n_97),
.B2(n_89),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_113),
.A2(n_151),
.B1(n_118),
.B2(n_103),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_77),
.A2(n_37),
.B1(n_29),
.B2(n_32),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_49),
.A2(n_30),
.B1(n_28),
.B2(n_44),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_55),
.B(n_52),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_145),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_83),
.B(n_22),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_141),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_91),
.A2(n_29),
.B1(n_27),
.B2(n_43),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_62),
.A2(n_44),
.B1(n_41),
.B2(n_36),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_84),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_51),
.B(n_41),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_50),
.A2(n_39),
.B1(n_40),
.B2(n_36),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_75),
.B(n_24),
.Y(n_145)
);

NAND2x1_ASAP7_75t_SL g172 ( 
.A(n_154),
.B(n_90),
.Y(n_172)
);

BUFx12_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_130),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_158),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_153),
.A2(n_133),
.B1(n_134),
.B2(n_139),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_160),
.A2(n_192),
.B1(n_159),
.B2(n_171),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_161),
.A2(n_177),
.B1(n_194),
.B2(n_107),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_135),
.A2(n_51),
.B(n_90),
.C(n_15),
.Y(n_162)
);

AOI21xp33_ASAP7_75t_L g208 ( 
.A1(n_162),
.A2(n_187),
.B(n_195),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_122),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_163),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_156),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_168),
.Y(n_209)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_58),
.B(n_48),
.C(n_67),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_166),
.A2(n_121),
.B(n_111),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_169),
.Y(n_217)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_116),
.Y(n_170)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_15),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_171),
.B(n_178),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_172),
.B(n_188),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_79),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_176),
.Y(n_214)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_116),
.Y(n_174)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_174),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_125),
.B(n_71),
.C(n_65),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_175),
.B(n_124),
.C(n_111),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_123),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_L g177 ( 
.A1(n_137),
.A2(n_70),
.B1(n_69),
.B2(n_68),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_115),
.B(n_0),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_129),
.B(n_66),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_186),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_0),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_181),
.B(n_189),
.Y(n_210)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_122),
.Y(n_183)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_185),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_105),
.Y(n_186)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_118),
.A2(n_88),
.B(n_23),
.C(n_94),
.Y(n_187)
);

AND2x2_ASAP7_75t_SL g188 ( 
.A(n_118),
.B(n_106),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_106),
.B(n_0),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_190),
.Y(n_228)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_140),
.B(n_66),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_197),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_142),
.A2(n_57),
.B1(n_23),
.B2(n_10),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_142),
.A2(n_57),
.B1(n_10),
.B2(n_9),
.Y(n_196)
);

OAI22x1_ASAP7_75t_L g233 ( 
.A1(n_196),
.A2(n_126),
.B1(n_100),
.B2(n_152),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_112),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_200),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_140),
.B(n_8),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_199),
.B(n_0),
.Y(n_223)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_146),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_112),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_114),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_124),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_202),
.B(n_172),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_165),
.A2(n_144),
.B1(n_132),
.B2(n_143),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_205),
.A2(n_218),
.B1(n_233),
.B2(n_166),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_207),
.A2(n_212),
.B1(n_230),
.B2(n_198),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_161),
.A2(n_165),
.B1(n_194),
.B2(n_162),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_165),
.A2(n_132),
.B1(n_143),
.B2(n_104),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_231),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_223),
.B(n_199),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_158),
.A2(n_107),
.B1(n_149),
.B2(n_128),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_188),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_234),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_169),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_163),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_236),
.B(n_249),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_212),
.A2(n_192),
.B1(n_179),
.B2(n_172),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_237),
.A2(n_262),
.B1(n_263),
.B2(n_226),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_221),
.Y(n_238)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_238),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_178),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_240),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_223),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_241),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_242),
.Y(n_288)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_214),
.B(n_176),
.Y(n_245)
);

INVxp33_ASAP7_75t_L g289 ( 
.A(n_245),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_184),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_246),
.B(n_251),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_228),
.Y(n_278)
);

AND2x2_ASAP7_75t_SL g248 ( 
.A(n_226),
.B(n_190),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_248),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_217),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_250),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_214),
.B(n_189),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_206),
.B(n_167),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_252),
.A2(n_255),
.B(n_261),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_181),
.Y(n_253)
);

A2O1A1O1Ixp25_ASAP7_75t_L g290 ( 
.A1(n_253),
.A2(n_254),
.B(n_227),
.C(n_188),
.D(n_193),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_202),
.B(n_188),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_164),
.Y(n_255)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_211),
.Y(n_258)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_231),
.A2(n_166),
.B(n_187),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_259),
.A2(n_213),
.B(n_229),
.Y(n_277)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_220),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_260),
.A2(n_241),
.B1(n_183),
.B2(n_235),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_209),
.B(n_173),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_226),
.C(n_222),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_268),
.C(n_278),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_266),
.B(n_273),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_206),
.Y(n_268)
);

AO22x1_ASAP7_75t_L g273 ( 
.A1(n_237),
.A2(n_205),
.B1(n_218),
.B2(n_208),
.Y(n_273)
);

FAx1_ASAP7_75t_SL g275 ( 
.A(n_248),
.B(n_213),
.CI(n_228),
.CON(n_275),
.SN(n_275)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_275),
.B(n_254),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_277),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_256),
.A2(n_229),
.B(n_219),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_281),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_256),
.A2(n_219),
.B(n_167),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_248),
.B(n_209),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_286),
.C(n_248),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_284),
.A2(n_291),
.B1(n_257),
.B2(n_264),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_237),
.A2(n_263),
.B1(n_253),
.B2(n_262),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_285),
.A2(n_243),
.B1(n_250),
.B2(n_260),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_248),
.B(n_227),
.C(n_175),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_256),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_242),
.A2(n_207),
.B1(n_227),
.B2(n_216),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_292),
.Y(n_320)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_293),
.Y(n_331)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_267),
.Y(n_295)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_295),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_273),
.A2(n_262),
.B1(n_256),
.B2(n_259),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_296),
.A2(n_298),
.B1(n_308),
.B2(n_314),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_297),
.B(n_233),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_273),
.A2(n_262),
.B1(n_259),
.B2(n_261),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_299),
.A2(n_269),
.B(n_277),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_300),
.B(n_303),
.C(n_318),
.Y(n_323)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_267),
.Y(n_301)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_301),
.Y(n_339)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_274),
.Y(n_302)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_302),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_254),
.C(n_251),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_274),
.Y(n_305)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_305),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_282),
.Y(n_306)
);

INVx4_ASAP7_75t_SL g340 ( 
.A(n_306),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_245),
.B1(n_242),
.B2(n_240),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_271),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_275),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_287),
.B(n_252),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_311),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_255),
.Y(n_312)
);

INVxp33_ASAP7_75t_SL g325 ( 
.A(n_312),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_313),
.A2(n_315),
.B1(n_317),
.B2(n_264),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_288),
.A2(n_246),
.B1(n_249),
.B2(n_239),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_285),
.A2(n_257),
.B1(n_244),
.B2(n_236),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_271),
.B(n_204),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_316),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_268),
.B(n_278),
.C(n_283),
.Y(n_318)
);

NOR2xp67_ASAP7_75t_SL g321 ( 
.A(n_300),
.B(n_281),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_321),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_312),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_322),
.B(n_258),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_314),
.Y(n_324)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_324),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_326),
.A2(n_327),
.B1(n_329),
.B2(n_336),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_309),
.A2(n_288),
.B1(n_266),
.B2(n_280),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_294),
.B(n_286),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_333),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_294),
.B(n_303),
.Y(n_333)
);

A2O1A1Ixp33_ASAP7_75t_L g334 ( 
.A1(n_307),
.A2(n_287),
.B(n_269),
.C(n_270),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_334),
.B(n_216),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_313),
.A2(n_270),
.B1(n_275),
.B2(n_276),
.Y(n_336)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_337),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_317),
.A2(n_276),
.B1(n_290),
.B2(n_279),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_341),
.A2(n_342),
.B1(n_238),
.B2(n_258),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_308),
.A2(n_279),
.B1(n_233),
.B2(n_241),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_318),
.B(n_180),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_343),
.B(n_293),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_345),
.B(n_241),
.Y(n_364)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_340),
.Y(n_348)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_348),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_324),
.A2(n_307),
.B1(n_315),
.B2(n_298),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_349),
.A2(n_363),
.B1(n_366),
.B2(n_225),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_338),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_350),
.B(n_361),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_330),
.B(n_304),
.C(n_296),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_356),
.C(n_357),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_326),
.A2(n_307),
.B1(n_304),
.B2(n_310),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_352),
.Y(n_375)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_340),
.Y(n_355)
);

BUFx4f_ASAP7_75t_SL g391 ( 
.A(n_355),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_333),
.B(n_306),
.C(n_310),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_323),
.B(n_311),
.C(n_295),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_337),
.A2(n_299),
.B(n_301),
.Y(n_358)
);

NOR2xp67_ASAP7_75t_SL g387 ( 
.A(n_358),
.B(n_225),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_359),
.B(n_353),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_327),
.A2(n_292),
.B(n_302),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_360),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_336),
.A2(n_305),
.B(n_203),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_364),
.B(n_368),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_365),
.A2(n_369),
.B1(n_332),
.B2(n_344),
.Y(n_379)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_332),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_367),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_323),
.B(n_343),
.Y(n_368)
);

OA22x2_ASAP7_75t_L g369 ( 
.A1(n_341),
.A2(n_238),
.B1(n_215),
.B2(n_203),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_325),
.B(n_238),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_370),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_372),
.B(n_234),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_353),
.B(n_334),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_377),
.B(n_381),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_379),
.A2(n_360),
.B1(n_349),
.B2(n_347),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_368),
.B(n_329),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_357),
.B(n_328),
.C(n_345),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_383),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_359),
.B(n_320),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_346),
.B(n_319),
.C(n_339),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_384),
.B(n_388),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_356),
.B(n_342),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_385),
.B(n_369),
.Y(n_400)
);

AO22x1_ASAP7_75t_L g386 ( 
.A1(n_354),
.A2(n_335),
.B1(n_331),
.B2(n_215),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_386),
.A2(n_183),
.B1(n_234),
.B2(n_200),
.Y(n_405)
);

OAI21x1_ASAP7_75t_SL g395 ( 
.A1(n_387),
.A2(n_363),
.B(n_358),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_351),
.B(n_197),
.C(n_211),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_389),
.B(n_364),
.C(n_370),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_392),
.B(n_400),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_380),
.A2(n_347),
.B1(n_362),
.B2(n_352),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_394),
.A2(n_405),
.B1(n_373),
.B2(n_146),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_395),
.A2(n_399),
.B(n_104),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_396),
.B(n_403),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_374),
.B(n_346),
.C(n_361),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_397),
.B(n_398),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_391),
.B(n_354),
.Y(n_398)
);

OAI22x1_ASAP7_75t_L g399 ( 
.A1(n_375),
.A2(n_369),
.B1(n_191),
.B2(n_182),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_376),
.A2(n_369),
.B1(n_185),
.B2(n_174),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_402),
.B(n_404),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_374),
.B(n_170),
.C(n_200),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_389),
.B(n_102),
.C(n_201),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_406),
.B(n_409),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_390),
.B(n_100),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_408),
.B(n_410),
.Y(n_425)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_386),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_378),
.B(n_102),
.C(n_152),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_393),
.A2(n_376),
.B(n_379),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_411),
.A2(n_119),
.B(n_157),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_397),
.B(n_385),
.C(n_382),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_413),
.B(n_416),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_403),
.B(n_378),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_415),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_396),
.B(n_371),
.C(n_391),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_401),
.B(n_391),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_417),
.B(n_421),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_420),
.A2(n_426),
.B1(n_127),
.B2(n_114),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_404),
.B(n_407),
.C(n_394),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_373),
.Y(n_423)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_423),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_410),
.B(n_149),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_424),
.B(n_138),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_428),
.B(n_434),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_413),
.B(n_399),
.C(n_138),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_429),
.B(n_431),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_415),
.B(n_119),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_430),
.B(n_436),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_416),
.B(n_128),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_412),
.A2(n_155),
.B(n_119),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_414),
.B(n_155),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_435),
.B(n_437),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_414),
.B(n_127),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_439),
.B(n_157),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_427),
.B(n_421),
.C(n_419),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_441),
.B(n_443),
.Y(n_452)
);

A2O1A1O1Ixp25_ASAP7_75t_L g442 ( 
.A1(n_438),
.A2(n_422),
.B(n_419),
.C(n_425),
.D(n_418),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_442),
.A2(n_449),
.B(n_440),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_433),
.B(n_420),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_432),
.B(n_424),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_445),
.B(n_446),
.Y(n_453)
);

NOR2xp67_ASAP7_75t_L g447 ( 
.A(n_432),
.B(n_157),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_447),
.A2(n_8),
.B(n_2),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_447),
.Y(n_450)
);

NOR3xp33_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_456),
.C(n_1),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_451),
.A2(n_454),
.B(n_455),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_444),
.B(n_429),
.C(n_436),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_448),
.A2(n_430),
.B(n_8),
.Y(n_455)
);

OAI311xp33_ASAP7_75t_L g458 ( 
.A1(n_452),
.A2(n_453),
.A3(n_2),
.B1(n_4),
.C1(n_5),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_458),
.A2(n_460),
.B(n_5),
.Y(n_463)
);

NOR3xp33_ASAP7_75t_L g461 ( 
.A(n_459),
.B(n_1),
.C(n_4),
.Y(n_461)
);

OAI21xp33_ASAP7_75t_L g460 ( 
.A1(n_452),
.A2(n_1),
.B(n_4),
.Y(n_460)
);

NAND2xp33_ASAP7_75t_SL g464 ( 
.A(n_461),
.B(n_462),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_457),
.A2(n_5),
.B1(n_6),
.B2(n_451),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_464),
.B(n_463),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_465),
.B(n_6),
.Y(n_466)
);


endmodule