module fake_ariane_852_n_442 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_44, n_30, n_82, n_31, n_42, n_57, n_70, n_10, n_117, n_85, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_112, n_45, n_11, n_126, n_122, n_52, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_442);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_117;
input n_85;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_112;
input n_45;
input n_11;
input n_126;
input n_122;
input n_52;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_442;

wire n_295;
wire n_356;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_332;
wire n_294;
wire n_197;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_373;
wire n_299;
wire n_133;
wire n_205;
wire n_341;
wire n_421;
wire n_245;
wire n_319;
wire n_416;
wire n_283;
wire n_187;
wire n_367;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_424;
wire n_387;
wire n_406;
wire n_139;
wire n_130;
wire n_349;
wire n_391;
wire n_346;
wire n_214;
wire n_348;
wire n_410;
wire n_379;
wire n_138;
wire n_162;
wire n_264;
wire n_137;
wire n_198;
wire n_232;
wire n_441;
wire n_385;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_399;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_167;
wire n_422;
wire n_153;
wire n_269;
wire n_158;
wire n_259;
wire n_143;
wire n_152;
wire n_405;
wire n_169;
wire n_173;
wire n_242;
wire n_309;
wire n_320;
wire n_331;
wire n_401;
wire n_267;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_200;
wire n_166;
wire n_253;
wire n_218;
wire n_271;
wire n_247;
wire n_240;
wire n_369;
wire n_128;
wire n_224;
wire n_420;
wire n_439;
wire n_222;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_330;
wire n_400;
wire n_129;
wire n_282;
wire n_328;
wire n_368;
wire n_277;
wire n_248;
wire n_301;
wire n_432;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_427;
wire n_303;
wire n_168;
wire n_206;
wire n_352;
wire n_238;
wire n_365;
wire n_429;
wire n_136;
wire n_334;
wire n_192;
wire n_300;
wire n_163;
wire n_141;
wire n_390;
wire n_438;
wire n_314;
wire n_440;
wire n_273;
wire n_305;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_413;
wire n_392;
wire n_376;
wire n_221;
wire n_321;
wire n_361;
wire n_149;
wire n_383;
wire n_237;
wire n_175;
wire n_181;
wire n_260;
wire n_362;
wire n_310;
wire n_236;
wire n_281;
wire n_209;
wire n_262;
wire n_225;
wire n_235;
wire n_297;
wire n_290;
wire n_371;
wire n_199;
wire n_217;
wire n_178;
wire n_308;
wire n_417;
wire n_201;
wire n_343;
wire n_414;
wire n_287;
wire n_302;
wire n_380;
wire n_284;
wire n_249;
wire n_212;
wire n_355;
wire n_278;
wire n_255;
wire n_257;
wire n_148;
wire n_135;
wire n_409;
wire n_171;
wire n_384;
wire n_182;
wire n_316;
wire n_196;
wire n_407;
wire n_254;
wire n_219;
wire n_231;
wire n_366;
wire n_234;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_298;
wire n_415;
wire n_216;
wire n_418;
wire n_223;
wire n_403;
wire n_389;
wire n_288;
wire n_179;
wire n_395;
wire n_195;
wire n_213;
wire n_304;
wire n_306;
wire n_313;
wire n_430;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_337;
wire n_437;
wire n_274;
wire n_296;
wire n_265;
wire n_208;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_132;
wire n_147;
wire n_204;
wire n_342;
wire n_246;
wire n_428;
wire n_159;
wire n_358;
wire n_131;
wire n_263;
wire n_434;
wire n_360;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_268;
wire n_266;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_411;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_191;
wire n_382;
wire n_211;
wire n_408;
wire n_322;
wire n_251;
wire n_397;
wire n_351;
wire n_393;
wire n_359;
wire n_155;

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_18),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_15),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_7),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_42),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_20),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_6),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_41),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_32),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_46),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_21),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_38),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_35),
.B(n_82),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_89),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_81),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_2),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g150 ( 
.A(n_49),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_27),
.Y(n_152)
);

INVxp67_ASAP7_75t_SL g153 ( 
.A(n_98),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_99),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_94),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_61),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_59),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_113),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_16),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_43),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_74),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_114),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_57),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_125),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_95),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_86),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_34),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_84),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_10),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_112),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_24),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_51),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_36),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_104),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_129),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_130),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_132),
.B(n_0),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_157),
.Y(n_185)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_150),
.B(n_0),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_133),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_137),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_138),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_139),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_140),
.Y(n_194)
);

OAI21x1_ASAP7_75t_L g195 ( 
.A1(n_171),
.A2(n_68),
.B(n_126),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_142),
.Y(n_196)
);

AND2x4_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_143),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_148),
.B(n_8),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_145),
.Y(n_200)
);

OAI21x1_ASAP7_75t_L g201 ( 
.A1(n_151),
.A2(n_69),
.B(n_123),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

O2A1O1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_183),
.B(n_191),
.C(n_199),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_155),
.Y(n_205)
);

NOR2xp67_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_152),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_158),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_198),
.B(n_163),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_185),
.B(n_166),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_156),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_197),
.A2(n_153),
.B(n_162),
.C(n_152),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_159),
.Y(n_214)
);

NAND2x1p5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_163),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_184),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_161),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_153),
.Y(n_219)
);

AND2x4_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_162),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_184),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_187),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_187),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_187),
.B(n_128),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_192),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_164),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_175),
.B1(n_173),
.B2(n_172),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_165),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_192),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_192),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_167),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_203),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_230),
.Y(n_233)
);

OR2x6_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_220),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_141),
.Y(n_235)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_230),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_205),
.B(n_147),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

A2O1A1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_204),
.A2(n_201),
.B(n_170),
.C(n_169),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

AND2x4_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_168),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_160),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_210),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_215),
.B(n_146),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_210),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_209),
.B(n_1),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_219),
.B(n_1),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

AND2x4_ASAP7_75t_L g255 ( 
.A(n_211),
.B(n_2),
.Y(n_255)
);

BUFx8_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_214),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_213),
.B(n_225),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_217),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_3),
.Y(n_260)
);

NAND2x1p5_ASAP7_75t_L g261 ( 
.A(n_224),
.B(n_3),
.Y(n_261)
);

AOI221xp5_ASAP7_75t_L g262 ( 
.A1(n_227),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.C(n_11),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_R g263 ( 
.A(n_228),
.B(n_12),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_231),
.A2(n_73),
.B(n_122),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_231),
.A2(n_4),
.B(n_5),
.C(n_13),
.Y(n_265)
);

NAND2x1_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_14),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_203),
.Y(n_267)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_230),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_220),
.B(n_17),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_215),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_205),
.B(n_19),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_230),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_203),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_22),
.Y(n_274)
);

AOI21xp33_ASAP7_75t_SL g275 ( 
.A1(n_234),
.A2(n_23),
.B(n_25),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_234),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_246),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_232),
.Y(n_278)
);

A2O1A1Ixp33_ASAP7_75t_SL g279 ( 
.A1(n_264),
.A2(n_127),
.B(n_28),
.C(n_29),
.Y(n_279)
);

OAI21xp33_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_26),
.B(n_30),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

INVx8_ASAP7_75t_L g282 ( 
.A(n_243),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_245),
.B(n_31),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_242),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_235),
.Y(n_285)
);

AND2x4_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_33),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_37),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_R g288 ( 
.A(n_256),
.B(n_39),
.Y(n_288)
);

INVx3_ASAP7_75t_SL g289 ( 
.A(n_255),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_244),
.B(n_40),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_118),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_258),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_249),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_242),
.Y(n_294)
);

INVxp67_ASAP7_75t_SL g295 ( 
.A(n_272),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_271),
.A2(n_44),
.B(n_45),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_238),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_254),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_270),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_252),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_300)
);

NAND2x1p5_ASAP7_75t_L g301 ( 
.A(n_236),
.B(n_52),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_237),
.A2(n_53),
.B(n_54),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_241),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_255),
.B(n_55),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_266),
.A2(n_58),
.B(n_60),
.Y(n_305)
);

A2O1A1Ixp33_ASAP7_75t_L g306 ( 
.A1(n_262),
.A2(n_240),
.B(n_265),
.C(n_248),
.Y(n_306)
);

BUFx4f_ASAP7_75t_SL g307 ( 
.A(n_239),
.Y(n_307)
);

NOR2x1_ASAP7_75t_SL g308 ( 
.A(n_236),
.B(n_62),
.Y(n_308)
);

AND2x4_ASAP7_75t_L g309 ( 
.A(n_247),
.B(n_63),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_233),
.Y(n_310)
);

INVx5_ASAP7_75t_L g311 ( 
.A(n_236),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_250),
.A2(n_64),
.B(n_65),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_261),
.B(n_117),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_263),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_285),
.B(n_268),
.Y(n_315)
);

OA21x2_ASAP7_75t_L g316 ( 
.A1(n_306),
.A2(n_268),
.B(n_67),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_278),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_281),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_282),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_297),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_276),
.B(n_268),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_66),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_282),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_293),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_286),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_303),
.Y(n_326)
);

OAI21x1_ASAP7_75t_L g327 ( 
.A1(n_305),
.A2(n_70),
.B(n_71),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_289),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_310),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_298),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_295),
.Y(n_331)
);

OAI21x1_ASAP7_75t_L g332 ( 
.A1(n_290),
.A2(n_75),
.B(n_76),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_294),
.Y(n_333)
);

OAI21x1_ASAP7_75t_L g334 ( 
.A1(n_291),
.A2(n_77),
.B(n_78),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_292),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_309),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_309),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_287),
.A2(n_79),
.B(n_80),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_274),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_294),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_277),
.B(n_83),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_284),
.B(n_85),
.Y(n_342)
);

OAI211xp5_ASAP7_75t_L g343 ( 
.A1(n_288),
.A2(n_88),
.B(n_90),
.C(n_92),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_308),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_283),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_311),
.B(n_93),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_317),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_324),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_325),
.B(n_314),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_319),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_335),
.B(n_304),
.Y(n_351)
);

BUFx2_ASAP7_75t_SL g352 ( 
.A(n_323),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_325),
.B(n_313),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_318),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_320),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_324),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_330),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_323),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_321),
.B(n_311),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_329),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_333),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_326),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_331),
.Y(n_363)
);

OR2x2_ASAP7_75t_L g364 ( 
.A(n_328),
.B(n_311),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_336),
.B(n_275),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_360),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_347),
.Y(n_367)
);

BUFx8_ASAP7_75t_L g368 ( 
.A(n_349),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_361),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_354),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_355),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_350),
.A2(n_337),
.B1(n_339),
.B2(n_315),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_350),
.Y(n_373)
);

AOI222xp33_ASAP7_75t_L g374 ( 
.A1(n_362),
.A2(n_335),
.B1(n_345),
.B2(n_338),
.C1(n_341),
.C2(n_322),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_357),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_353),
.B(n_340),
.Y(n_376)
);

INVx3_ASAP7_75t_R g377 ( 
.A(n_364),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_358),
.B(n_333),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_363),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_361),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_373),
.Y(n_381)
);

AND2x2_ASAP7_75t_SL g382 ( 
.A(n_378),
.B(n_380),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_367),
.Y(n_383)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_370),
.B(n_358),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_376),
.B(n_351),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_371),
.B(n_333),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_368),
.B(n_307),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_366),
.B(n_352),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_375),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_379),
.B(n_348),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_369),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_369),
.B(n_359),
.Y(n_392)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_368),
.Y(n_393)
);

NAND2x1_ASAP7_75t_L g394 ( 
.A(n_372),
.B(n_344),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_374),
.B(n_351),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_374),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_377),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_356),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_384),
.B(n_356),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_365),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_386),
.B(n_346),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_315),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_392),
.Y(n_403)
);

NAND2x1p5_ASAP7_75t_L g404 ( 
.A(n_393),
.B(n_346),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_383),
.B(n_342),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_395),
.B(n_344),
.Y(n_406)
);

NOR2x1_ASAP7_75t_L g407 ( 
.A(n_393),
.B(n_343),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_392),
.B(n_338),
.Y(n_408)
);

AOI221xp5_ASAP7_75t_L g409 ( 
.A1(n_396),
.A2(n_280),
.B1(n_302),
.B2(n_343),
.C(n_300),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_391),
.B(n_316),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_389),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_387),
.B(n_301),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_388),
.B(n_316),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_397),
.B(n_296),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_390),
.B(n_312),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_403),
.B(n_394),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_411),
.Y(n_417)
);

NAND3xp33_ASAP7_75t_L g418 ( 
.A(n_414),
.B(n_279),
.C(n_332),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_402),
.B(n_334),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_398),
.Y(n_420)
);

OAI31xp33_ASAP7_75t_L g421 ( 
.A1(n_400),
.A2(n_96),
.A3(n_97),
.B(n_100),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_406),
.B(n_101),
.Y(n_422)
);

NOR2x1_ASAP7_75t_L g423 ( 
.A(n_407),
.B(n_327),
.Y(n_423)
);

AOI21xp33_ASAP7_75t_SL g424 ( 
.A1(n_404),
.A2(n_102),
.B(n_103),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_417),
.Y(n_425)
);

NAND4xp25_ASAP7_75t_L g426 ( 
.A(n_419),
.B(n_418),
.C(n_412),
.D(n_421),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_420),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_422),
.B(n_403),
.Y(n_428)
);

NOR4xp25_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_405),
.C(n_415),
.D(n_401),
.Y(n_429)
);

AOI211xp5_ASAP7_75t_L g430 ( 
.A1(n_429),
.A2(n_424),
.B(n_408),
.C(n_409),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_427),
.B(n_399),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_426),
.A2(n_408),
.B1(n_413),
.B2(n_423),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_425),
.B(n_428),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_433),
.Y(n_434)
);

NOR3x2_ASAP7_75t_L g435 ( 
.A(n_430),
.B(n_410),
.C(n_106),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_434),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_435),
.Y(n_437)
);

AOI211xp5_ASAP7_75t_L g438 ( 
.A1(n_437),
.A2(n_432),
.B(n_436),
.C(n_431),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_438),
.B(n_105),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_439),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_440),
.Y(n_441)
);

AOI221xp5_ASAP7_75t_L g442 ( 
.A1(n_441),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.C(n_111),
.Y(n_442)
);


endmodule