module fake_jpeg_3218_n_461 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_461);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_461;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_10),
.B(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_25),
.B(n_15),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_48),
.B(n_56),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_25),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_51),
.B(n_57),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_53),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_54),
.Y(n_136)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_29),
.B(n_12),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_37),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_29),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_58),
.B(n_62),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_59),
.Y(n_142)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_18),
.B(n_0),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_63),
.Y(n_148)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_64),
.Y(n_149)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_26),
.B(n_0),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_65),
.B(n_93),
.Y(n_130)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_66),
.Y(n_150)
);

BUFx8_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_11),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_68),
.B(n_27),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_18),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_71),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_39),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_79),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_42),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

BUFx4f_ASAP7_75t_SL g84 ( 
.A(n_17),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_38),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_21),
.Y(n_90)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_19),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_95),
.Y(n_133)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_98),
.B(n_120),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_67),
.A2(n_38),
.B1(n_44),
.B2(n_42),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_103),
.A2(n_104),
.B1(n_128),
.B2(n_145),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_67),
.A2(n_87),
.B1(n_88),
.B2(n_86),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_111),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_55),
.A2(n_27),
.B1(n_45),
.B2(n_40),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_113),
.A2(n_31),
.B1(n_35),
.B2(n_33),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_94),
.B(n_44),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_36),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_127),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_36),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_80),
.A2(n_38),
.B1(n_46),
.B2(n_32),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_46),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_140),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_59),
.A2(n_63),
.B1(n_52),
.B2(n_53),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_135),
.A2(n_146),
.B1(n_11),
.B2(n_2),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_84),
.B(n_46),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_139),
.B(n_43),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_82),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_85),
.A2(n_24),
.B1(n_32),
.B2(n_19),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_49),
.A2(n_24),
.B1(n_32),
.B2(n_40),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_65),
.B(n_45),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_35),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_130),
.A2(n_65),
.B1(n_54),
.B2(n_74),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_151),
.A2(n_155),
.B1(n_171),
.B2(n_189),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_130),
.A2(n_61),
.B1(n_64),
.B2(n_69),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_152),
.A2(n_99),
.B(n_112),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_154),
.B(n_173),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_72),
.B1(n_91),
.B2(n_89),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_83),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_158),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_108),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_159),
.B(n_163),
.Y(n_236)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_161),
.Y(n_210)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_118),
.Y(n_162)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_162),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_150),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_164),
.Y(n_229)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_165),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_137),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_166),
.B(n_170),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_167),
.A2(n_193),
.B1(n_196),
.B2(n_197),
.Y(n_207)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

INVx2_ASAP7_75t_R g169 ( 
.A(n_123),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_169),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_114),
.B(n_75),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_103),
.A2(n_78),
.B1(n_76),
.B2(n_85),
.Y(n_171)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_172),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_109),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_175),
.B(n_186),
.Y(n_235)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_176),
.Y(n_240)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_116),
.B(n_43),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_178),
.B(n_183),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_102),
.A2(n_33),
.B(n_31),
.C(n_34),
.Y(n_179)
);

OA21x2_ASAP7_75t_L g214 ( 
.A1(n_179),
.A2(n_149),
.B(n_100),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_106),
.B(n_66),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_181),
.Y(n_231)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_132),
.Y(n_182)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_113),
.B(n_34),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_97),
.Y(n_184)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_184),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_101),
.Y(n_185)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_185),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_105),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_143),
.B(n_66),
.C(n_90),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_119),
.C(n_126),
.Y(n_206)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_104),
.A2(n_145),
.B1(n_148),
.B2(n_142),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_96),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_96),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_144),
.B(n_1),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_198),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_110),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_144),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_142),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_123),
.B(n_2),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_126),
.Y(n_199)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_112),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_200),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_201),
.Y(n_230)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_134),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_117),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_183),
.A2(n_121),
.B1(n_136),
.B2(n_131),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_203),
.A2(n_224),
.B1(n_231),
.B2(n_227),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_206),
.B(n_185),
.Y(n_279)
);

OAI21xp33_ASAP7_75t_L g271 ( 
.A1(n_214),
.A2(n_232),
.B(n_241),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_167),
.A2(n_105),
.B1(n_148),
.B2(n_131),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_178),
.A2(n_136),
.B1(n_99),
.B2(n_115),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_226),
.A2(n_241),
.B1(n_246),
.B2(n_171),
.Y(n_250)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_166),
.B(n_110),
.C(n_100),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_181),
.C(n_199),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_152),
.A2(n_115),
.B1(n_117),
.B2(n_6),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_242),
.B(n_180),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_153),
.B(n_4),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_244),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_194),
.B(n_4),
.Y(n_244)
);

OAI32xp33_ASAP7_75t_L g245 ( 
.A1(n_161),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_7),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_191),
.A2(n_151),
.B1(n_157),
.B2(n_189),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_216),
.Y(n_247)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_247),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_236),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_248),
.B(n_265),
.Y(n_313)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_216),
.Y(n_249)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_249),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_250),
.A2(n_253),
.B1(n_255),
.B2(n_256),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_213),
.A2(n_191),
.B1(n_155),
.B2(n_156),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_251),
.A2(n_258),
.B1(n_274),
.B2(n_284),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_213),
.A2(n_191),
.B1(n_197),
.B2(n_170),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_174),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_254),
.B(n_262),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_246),
.A2(n_223),
.B1(n_207),
.B2(n_221),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_223),
.A2(n_191),
.B1(n_158),
.B2(n_179),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_242),
.Y(n_257)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_257),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_221),
.A2(n_158),
.B1(n_187),
.B2(n_172),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_234),
.Y(n_259)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_259),
.Y(n_304)
);

XNOR2x1_ASAP7_75t_L g316 ( 
.A(n_260),
.B(n_279),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_181),
.C(n_165),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_261),
.B(n_283),
.C(n_222),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_188),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_214),
.A2(n_169),
.B(n_199),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_263),
.A2(n_211),
.B(n_222),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_280),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_176),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_164),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_266),
.B(n_270),
.Y(n_315)
);

OAI21xp33_ASAP7_75t_SL g292 ( 
.A1(n_267),
.A2(n_271),
.B(n_278),
.Y(n_292)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_217),
.Y(n_268)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_268),
.Y(n_309)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_217),
.Y(n_269)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_269),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_214),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_204),
.B(n_162),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_272),
.B(n_277),
.Y(n_320)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_229),
.Y(n_273)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_273),
.Y(n_312)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_229),
.Y(n_275)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_275),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_230),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_276),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_225),
.B(n_177),
.Y(n_277)
);

OA21x2_ASAP7_75t_L g278 ( 
.A1(n_226),
.A2(n_192),
.B(n_200),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_201),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_228),
.B(n_160),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_263),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_206),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_282),
.A2(n_209),
.B1(n_212),
.B2(n_205),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_228),
.B(n_7),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_210),
.A2(n_9),
.B1(n_10),
.B2(n_219),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_210),
.A2(n_9),
.B1(n_232),
.B2(n_245),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_285),
.A2(n_234),
.B1(n_208),
.B2(n_230),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_287),
.B(n_249),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_225),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_289),
.B(n_295),
.C(n_296),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_301),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_294),
.A2(n_317),
.B(n_299),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_261),
.B(n_212),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_260),
.B(n_215),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_255),
.B(n_233),
.Y(n_297)
);

MAJx2_ASAP7_75t_L g335 ( 
.A(n_297),
.B(n_268),
.C(n_275),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_253),
.A2(n_208),
.B1(n_233),
.B2(n_215),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_299),
.A2(n_250),
.B1(n_278),
.B2(n_247),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_300),
.B(n_259),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_238),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_302),
.B(n_306),
.C(n_319),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_257),
.B(n_238),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_273),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_258),
.B(n_240),
.C(n_211),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_276),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_276),
.Y(n_324)
);

BUFx5_ASAP7_75t_L g311 ( 
.A(n_269),
.Y(n_311)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_311),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_256),
.A2(n_218),
.B(n_240),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_283),
.B(n_218),
.Y(n_319)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_322),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_305),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_323),
.B(n_341),
.Y(n_376)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_324),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_313),
.B(n_252),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_325),
.B(n_327),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_286),
.B(n_252),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_328),
.A2(n_333),
.B1(n_298),
.B2(n_314),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_280),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_329),
.B(n_344),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_291),
.B(n_318),
.Y(n_330)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_330),
.Y(n_352)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_303),
.Y(n_331)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_331),
.Y(n_355)
);

OAI22x1_ASAP7_75t_SL g332 ( 
.A1(n_290),
.A2(n_251),
.B1(n_285),
.B2(n_267),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_332),
.A2(n_293),
.B1(n_296),
.B2(n_319),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_288),
.A2(n_278),
.B1(n_282),
.B2(n_284),
.Y(n_333)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_334),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_335),
.B(n_295),
.Y(n_365)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_307),
.Y(n_338)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_338),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_339),
.B(n_326),
.C(n_336),
.Y(n_374)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_309),
.Y(n_340)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_340),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_301),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_291),
.B(n_259),
.Y(n_342)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_342),
.Y(n_366)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_312),
.Y(n_343)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_343),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_315),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_300),
.B(n_318),
.Y(n_345)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_345),
.Y(n_371)
);

AO22x2_ASAP7_75t_L g346 ( 
.A1(n_294),
.A2(n_297),
.B1(n_287),
.B2(n_292),
.Y(n_346)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_346),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_302),
.B(n_306),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_347),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_317),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_348),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_349),
.A2(n_350),
.B(n_334),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_290),
.A2(n_316),
.B(n_289),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_360),
.A2(n_367),
.B1(n_368),
.B2(n_369),
.Y(n_394)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_362),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_365),
.B(n_342),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_332),
.A2(n_304),
.B1(n_310),
.B2(n_316),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_321),
.A2(n_304),
.B1(n_311),
.B2(n_341),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_321),
.A2(n_348),
.B1(n_333),
.B2(n_328),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_372),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_326),
.B(n_350),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_373),
.B(n_346),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_374),
.B(n_373),
.C(n_339),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_349),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_375),
.B(n_346),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_377),
.B(n_379),
.C(n_380),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_374),
.B(n_336),
.C(n_347),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_371),
.B(n_335),
.C(n_344),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_376),
.Y(n_381)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_381),
.Y(n_399)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_376),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_382),
.B(n_391),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_375),
.A2(n_323),
.B(n_330),
.Y(n_383)
);

XOR2x1_ASAP7_75t_L g406 ( 
.A(n_383),
.B(n_381),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_354),
.B(n_325),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_384),
.B(n_386),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_353),
.B(n_331),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_387),
.A2(n_346),
.B(n_391),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_388),
.B(n_392),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_363),
.B(n_322),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_389),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_361),
.B(n_340),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_390),
.A2(n_351),
.B1(n_352),
.B2(n_366),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_363),
.B(n_343),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_356),
.B(n_338),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_393),
.B(n_358),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_355),
.B(n_337),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_395),
.B(n_396),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_368),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_351),
.B(n_337),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_357),
.Y(n_410)
);

AO21x1_ASAP7_75t_L g398 ( 
.A1(n_387),
.A2(n_364),
.B(n_359),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_398),
.B(n_382),
.Y(n_415)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_400),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_385),
.A2(n_359),
.B(n_372),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_403),
.B(n_385),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_396),
.A2(n_369),
.B1(n_360),
.B2(n_367),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_405),
.A2(n_411),
.B1(n_413),
.B2(n_394),
.Y(n_422)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_406),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_407),
.A2(n_408),
.B1(n_389),
.B2(n_397),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_390),
.A2(n_352),
.B1(n_359),
.B2(n_366),
.Y(n_408)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_410),
.Y(n_428)
);

AO221x1_ASAP7_75t_L g411 ( 
.A1(n_383),
.A2(n_364),
.B1(n_346),
.B2(n_370),
.C(n_365),
.Y(n_411)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_415),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_412),
.B(n_380),
.Y(n_416)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_416),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_417),
.B(n_421),
.Y(n_438)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_419),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_412),
.B(n_378),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_420),
.B(n_424),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_409),
.B(n_392),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_422),
.A2(n_414),
.B1(n_399),
.B2(n_413),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_409),
.B(n_377),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_423),
.B(n_406),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_401),
.B(n_379),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_401),
.B(n_388),
.C(n_394),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_425),
.B(n_427),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_405),
.B(n_378),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_429),
.B(n_411),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_424),
.B(n_414),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_434),
.B(n_439),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_435),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_426),
.A2(n_403),
.B(n_398),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_437),
.A2(n_415),
.B(n_435),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_422),
.A2(n_399),
.B1(n_404),
.B2(n_402),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_433),
.A2(n_398),
.B(n_402),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_440),
.A2(n_437),
.B(n_430),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_441),
.B(n_438),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_431),
.B(n_418),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_442),
.B(n_443),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_432),
.A2(n_425),
.B(n_417),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_436),
.B(n_428),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_444),
.B(n_447),
.Y(n_451)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_448),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_445),
.B(n_438),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_450),
.B(n_429),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_452),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_454),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_455),
.B(n_449),
.C(n_451),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_457),
.B(n_453),
.C(n_448),
.Y(n_458)
);

BUFx24_ASAP7_75t_SL g459 ( 
.A(n_458),
.Y(n_459)
);

AOI322xp5_ASAP7_75t_L g460 ( 
.A1(n_459),
.A2(n_456),
.A3(n_444),
.B1(n_446),
.B2(n_404),
.C1(n_439),
.C2(n_395),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_460),
.A2(n_423),
.B(n_421),
.Y(n_461)
);


endmodule