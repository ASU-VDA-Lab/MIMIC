module fake_jpeg_5314_n_327 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_10),
.B(n_8),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_43),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_21),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_41),
.B(n_44),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_20),
.Y(n_42)
);

HAxp5_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_33),
.CON(n_55),
.SN(n_55)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_46),
.Y(n_94)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_48),
.Y(n_79)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_18),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_18),
.Y(n_78)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_52),
.Y(n_89)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_27),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_58),
.Y(n_71)
);

NOR3xp33_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_19),
.C(n_22),
.Y(n_90)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_27),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_61),
.Y(n_80)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_83),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_73),
.B(n_78),
.Y(n_107)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_75),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_19),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_29),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_43),
.B1(n_37),
.B2(n_17),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_81),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_104)
);

CKINVDCx12_ASAP7_75t_R g83 ( 
.A(n_50),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_90),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_55),
.A2(n_37),
.B1(n_17),
.B2(n_32),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_67),
.A2(n_37),
.B1(n_17),
.B2(n_32),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_57),
.A2(n_43),
.B1(n_34),
.B2(n_36),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_63),
.A2(n_24),
.B1(n_22),
.B2(n_29),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_24),
.Y(n_113)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_98),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_97),
.B(n_94),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

AO22x1_ASAP7_75t_SL g100 ( 
.A1(n_86),
.A2(n_57),
.B1(n_60),
.B2(n_34),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_100),
.A2(n_119),
.B1(n_82),
.B2(n_52),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_61),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_101),
.B(n_111),
.Y(n_133)
);

BUFx4f_ASAP7_75t_SL g103 ( 
.A(n_91),
.Y(n_103)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_106),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_130)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_89),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_78),
.B(n_73),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_115),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_80),
.Y(n_117)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_88),
.A2(n_34),
.B1(n_36),
.B2(n_51),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_121),
.Y(n_125)
);

NAND2xp33_ASAP7_75t_SL g122 ( 
.A(n_85),
.B(n_20),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_80),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_71),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_122),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_128),
.B(n_135),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_85),
.Y(n_129)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_99),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_132),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_102),
.B(n_71),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_117),
.B1(n_106),
.B2(n_105),
.Y(n_168)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_141),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_SL g160 ( 
.A1(n_140),
.A2(n_20),
.B(n_36),
.Y(n_160)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_142),
.A2(n_143),
.B1(n_145),
.B2(n_147),
.Y(n_156)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_151),
.B(n_164),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_145),
.A2(n_104),
.B1(n_100),
.B2(n_119),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_152),
.A2(n_16),
.B1(n_28),
.B2(n_30),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_144),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_165),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_155),
.C(n_163),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_100),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_53),
.B1(n_92),
.B2(n_108),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_157),
.A2(n_168),
.B1(n_170),
.B2(n_137),
.Y(n_193)
);

XNOR2x2_ASAP7_75t_SL g158 ( 
.A(n_140),
.B(n_49),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_160),
.B(n_20),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_138),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_159),
.B(n_161),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_132),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_162),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_120),
.C(n_59),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_130),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_166),
.B(n_127),
.Y(n_187)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_169),
.Y(n_191)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_124),
.A2(n_114),
.B1(n_74),
.B2(n_116),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_125),
.A2(n_116),
.B1(n_110),
.B2(n_70),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_172),
.A2(n_175),
.B1(n_127),
.B2(n_123),
.Y(n_188)
);

NAND3xp33_ASAP7_75t_L g173 ( 
.A(n_125),
.B(n_66),
.C(n_39),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_SL g195 ( 
.A(n_173),
.B(n_148),
.C(n_39),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_134),
.B1(n_139),
.B2(n_142),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_146),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_143),
.B(n_134),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_177),
.A2(n_156),
.B(n_167),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_151),
.Y(n_178)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_178),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_148),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_201),
.C(n_60),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_199),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_66),
.Y(n_182)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_189),
.Y(n_213)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_188),
.Y(n_223)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_192),
.Y(n_215)
);

AND2x6_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_148),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_193),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_137),
.B1(n_109),
.B2(n_141),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_194),
.A2(n_149),
.B1(n_153),
.B2(n_176),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_196),
.Y(n_217)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_197),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_175),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_174),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_153),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_200),
.A2(n_70),
.B1(n_112),
.B2(n_146),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_66),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_131),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_131),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_150),
.B(n_164),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_20),
.Y(n_212)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_186),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_209),
.A2(n_227),
.B(n_228),
.Y(n_247)
);

AOI21xp33_ASAP7_75t_L g210 ( 
.A1(n_192),
.A2(n_66),
.B(n_75),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_210),
.A2(n_200),
.B(n_195),
.C(n_199),
.Y(n_239)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_224),
.Y(n_229)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_178),
.A2(n_25),
.B(n_33),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_214),
.A2(n_21),
.B(n_30),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_33),
.Y(n_218)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_186),
.C(n_201),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_33),
.Y(n_221)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_221),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_222),
.Y(n_249)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_225),
.A2(n_196),
.B1(n_189),
.B2(n_184),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_180),
.A2(n_30),
.B1(n_28),
.B2(n_16),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_190),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_185),
.B(n_33),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_1),
.Y(n_228)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_224),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_243),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_233),
.C(n_235),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_236),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_179),
.C(n_198),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_181),
.C(n_177),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_188),
.Y(n_236)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_238),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_239),
.A2(n_205),
.B(n_217),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_240),
.A2(n_250),
.B1(n_226),
.B2(n_206),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_25),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_246),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_223),
.A2(n_204),
.B1(n_211),
.B2(n_220),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_242),
.A2(n_245),
.B(n_209),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_213),
.B(n_208),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_146),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_223),
.A2(n_30),
.B1(n_28),
.B2(n_16),
.Y(n_250)
);

INVxp33_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_234),
.A2(n_204),
.B1(n_205),
.B2(n_216),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_252),
.A2(n_261),
.B1(n_262),
.B2(n_242),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_239),
.B(n_244),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_254),
.A2(n_258),
.B(n_263),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_256),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_249),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_212),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_268),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_208),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_248),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_237),
.A2(n_220),
.B1(n_227),
.B2(n_218),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_247),
.A2(n_221),
.B1(n_228),
.B2(n_28),
.Y(n_262)
);

NOR2xp67_ASAP7_75t_SL g263 ( 
.A(n_231),
.B(n_235),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_16),
.C(n_74),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_246),
.C(n_250),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_232),
.B(n_9),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_269),
.A2(n_270),
.B(n_279),
.Y(n_290)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_257),
.C(n_264),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_241),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_281),
.Y(n_296)
);

NAND2xp33_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_7),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_275),
.A2(n_11),
.B(n_4),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_267),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_278)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_278),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_255),
.A2(n_10),
.B(n_14),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_2),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_283),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_10),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_268),
.B(n_11),
.Y(n_283)
);

NOR2x1_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_251),
.Y(n_284)
);

XOR2x1_ASAP7_75t_SL g305 ( 
.A(n_284),
.B(n_12),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_265),
.Y(n_285)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_289),
.C(n_292),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_264),
.C(n_265),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_291),
.A2(n_270),
.B1(n_276),
.B2(n_282),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_11),
.C(n_4),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_7),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_295),
.Y(n_297)
);

BUFx24_ASAP7_75t_SL g295 ( 
.A(n_273),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_298),
.B(n_302),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_290),
.A2(n_277),
.B(n_272),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_299),
.A2(n_303),
.B(n_304),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_287),
.B(n_12),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_3),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_284),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_6),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_12),
.C(n_4),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_296),
.C(n_291),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_308),
.B(n_311),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_300),
.A2(n_288),
.B(n_3),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_309),
.A2(n_310),
.B(n_314),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_301),
.B(n_5),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_297),
.B(n_6),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_313),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_6),
.C(n_13),
.Y(n_314)
);

NAND3xp33_ASAP7_75t_SL g316 ( 
.A(n_312),
.B(n_304),
.C(n_14),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_316),
.A2(n_318),
.B(n_13),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_13),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_307),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_321),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_322),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_323),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_319),
.B1(n_317),
.B2(n_15),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_15),
.B(n_291),
.Y(n_327)
);


endmodule