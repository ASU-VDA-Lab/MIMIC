module fake_jpeg_26571_n_116 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_116);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_116;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx11_ASAP7_75t_SL g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_21),
.Y(n_28)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx3_ASAP7_75t_SL g22 ( 
.A(n_11),
.Y(n_22)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_23),
.A2(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_0),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_26),
.B1(n_31),
.B2(n_22),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_22),
.A2(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_21),
.A2(n_13),
.B1(n_12),
.B2(n_10),
.Y(n_31)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_23),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_40),
.B(n_23),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_22),
.B1(n_29),
.B2(n_39),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_28),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_12),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_47),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_50),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_33),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_26),
.B(n_22),
.C(n_29),
.Y(n_55)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_21),
.B1(n_22),
.B2(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_20),
.Y(n_61)
);

NOR2x1_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_42),
.B(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_61),
.B(n_45),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_29),
.B1(n_21),
.B2(n_34),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_13),
.Y(n_57)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_20),
.C(n_23),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_59),
.C(n_44),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_10),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_45),
.B1(n_29),
.B2(n_47),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_27),
.B1(n_18),
.B2(n_20),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_56),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_63),
.B(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_24),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_20),
.B(n_51),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_44),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_67),
.B(n_59),
.Y(n_72)
);

OA21x2_ASAP7_75t_SL g83 ( 
.A1(n_72),
.A2(n_76),
.B(n_4),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_66),
.A2(n_60),
.B1(n_55),
.B2(n_58),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_64),
.C(n_70),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_77),
.C(n_62),
.Y(n_82)
);

OAI322xp33_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_6),
.A3(n_8),
.B1(n_2),
.B2(n_4),
.C1(n_5),
.C2(n_7),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_0),
.B(n_1),
.Y(n_79)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

MAJx2_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_89),
.C(n_79),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_7),
.B(n_8),
.Y(n_96)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_84),
.B(n_87),
.Y(n_95)
);

XNOR2x1_ASAP7_75t_SL g86 ( 
.A(n_75),
.B(n_66),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_86),
.B(n_5),
.Y(n_94)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

OAI21x1_ASAP7_75t_SL g88 ( 
.A1(n_81),
.A2(n_51),
.B(n_4),
.Y(n_88)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_20),
.C(n_27),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_94),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_86),
.A2(n_5),
.B(n_6),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_92),
.A2(n_1),
.B(n_24),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_87),
.A2(n_27),
.B1(n_18),
.B2(n_7),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_1),
.B(n_24),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_96),
.B(n_97),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_99),
.B(n_100),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_95),
.A2(n_82),
.B1(n_85),
.B2(n_89),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_95),
.A2(n_90),
.B1(n_27),
.B2(n_18),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_102),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_103),
.A2(n_19),
.B(n_32),
.Y(n_106)
);

NOR2xp67_ASAP7_75t_SL g105 ( 
.A(n_100),
.B(n_1),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_105),
.A2(n_107),
.B(n_101),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_32),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_110),
.C(n_98),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_109),
.A2(n_32),
.B(n_19),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_98),
.C(n_32),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_111),
.A2(n_112),
.B(n_19),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_19),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_19),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_115),
.B(n_18),
.Y(n_116)
);


endmodule