module real_aes_10093_n_8 (n_4, n_0, n_3, n_5, n_2, n_7, n_6, n_1, n_8);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_6;
input n_1;
output n_8;
wire n_17;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_25;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_9;
wire n_23;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_10;
NAND2xp5_ASAP7_75t_SL g11 ( .A(n_0), .B(n_12), .Y(n_11) );
INVx1_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
OAI22xp5_ASAP7_75t_L g17 ( .A1(n_2), .A2(n_18), .B1(n_20), .B2(n_22), .Y(n_17) );
INVx1_ASAP7_75t_L g22 ( .A(n_2), .Y(n_22) );
HB1xp67_ASAP7_75t_L g26 ( .A(n_3), .Y(n_26) );
AND2x2_ASAP7_75t_L g14 ( .A(n_4), .B(n_15), .Y(n_14) );
INVx1_ASAP7_75t_L g25 ( .A(n_4), .Y(n_25) );
INVx1_ASAP7_75t_L g16 ( .A(n_5), .Y(n_16) );
BUFx10_ASAP7_75t_L g19 ( .A(n_6), .Y(n_19) );
INVx1_ASAP7_75t_L g10 ( .A(n_7), .Y(n_10) );
AOI21xp5_ASAP7_75t_L g8 ( .A1(n_9), .A2(n_17), .B(n_23), .Y(n_8) );
NOR2x1_ASAP7_75t_L g9 ( .A(n_10), .B(n_11), .Y(n_9) );
INVx1_ASAP7_75t_L g12 ( .A(n_13), .Y(n_12) );
NAND2xp5_ASAP7_75t_SL g13 ( .A(n_14), .B(n_16), .Y(n_13) );
NAND3xp33_ASAP7_75t_SL g24 ( .A(n_15), .B(n_25), .C(n_26), .Y(n_24) );
BUFx12f_ASAP7_75t_L g18 ( .A(n_19), .Y(n_18) );
INVx2_ASAP7_75t_SL g21 ( .A(n_19), .Y(n_21) );
BUFx2_ASAP7_75t_L g20 ( .A(n_21), .Y(n_20) );
CKINVDCx20_ASAP7_75t_R g23 ( .A(n_24), .Y(n_23) );
endmodule