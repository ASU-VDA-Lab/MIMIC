module real_jpeg_25636_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_292;
wire n_221;
wire n_249;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_200;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_258;
wire n_195;
wire n_205;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_213;
wire n_138;
wire n_257;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_269;
wire n_253;
wire n_96;
wire n_273;
wire n_89;

INVx3_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_1),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_1),
.A2(n_59),
.B1(n_60),
.B2(n_69),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_1),
.A2(n_40),
.B1(n_41),
.B2(n_69),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_69),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_2),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_2),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_2),
.A2(n_59),
.B1(n_60),
.B2(n_86),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_2),
.A2(n_40),
.B1(n_41),
.B2(n_86),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_86),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_3),
.B(n_72),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_3),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_3),
.B(n_80),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_3),
.B(n_41),
.C(n_56),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_3),
.A2(n_59),
.B1(n_60),
.B2(n_183),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_3),
.B(n_152),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_183),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_3),
.B(n_28),
.C(n_46),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_3),
.A2(n_30),
.B(n_245),
.Y(n_270)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g77 ( 
.A(n_6),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_7),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_7),
.A2(n_43),
.B1(n_59),
.B2(n_60),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_43),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_9),
.A2(n_29),
.B1(n_40),
.B2(n_41),
.Y(n_95)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_11),
.A2(n_72),
.B1(n_85),
.B2(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_11),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_11),
.A2(n_59),
.B1(n_60),
.B2(n_133),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_11),
.A2(n_40),
.B1(n_41),
.B2(n_133),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_133),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_12),
.A2(n_40),
.B1(n_41),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_12),
.A2(n_51),
.B1(n_59),
.B2(n_60),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_51),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_13),
.A2(n_59),
.B1(n_60),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_13),
.A2(n_64),
.B1(n_85),
.B2(n_110),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_64),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_64),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_15),
.A2(n_33),
.B1(n_40),
.B2(n_41),
.Y(n_96)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_16),
.Y(n_102)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_16),
.Y(n_162)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_16),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_16),
.A2(n_158),
.B1(n_257),
.B2(n_259),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_136),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_134),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_114),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_20),
.B(n_114),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_87),
.B2(n_113),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_53),
.C(n_66),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_23),
.A2(n_24),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_25),
.A2(n_36),
.B1(n_37),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_25),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_26),
.A2(n_30),
.B1(n_31),
.B2(n_122),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_27),
.A2(n_28),
.B1(n_46),
.B2(n_48),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_27),
.B(n_269),
.Y(n_268)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_30),
.A2(n_32),
.B(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_30),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_30),
.A2(n_160),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_30),
.B(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_30),
.A2(n_244),
.B(n_245),
.Y(n_243)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_31),
.Y(n_213)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_44),
.B1(n_50),
.B2(n_52),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_39),
.A2(n_49),
.B1(n_93),
.B2(n_125),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_41),
.B1(n_46),
.B2(n_48),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_41),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_41),
.B(n_253),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_44),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_44),
.A2(n_50),
.B1(n_52),
.B2(n_95),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_44),
.B(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_44),
.A2(n_52),
.B1(n_217),
.B2(n_219),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_49),
.Y(n_44)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_49),
.A2(n_93),
.B1(n_94),
.B2(n_96),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_49),
.A2(n_125),
.B(n_176),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_49),
.A2(n_176),
.B(n_218),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_49),
.B(n_183),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_52),
.B(n_177),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_53),
.B(n_66),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_63),
.B2(n_65),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_54),
.A2(n_55),
.B1(n_65),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_54),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_54),
.A2(n_149),
.B(n_151),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_L g221 ( 
.A1(n_54),
.A2(n_151),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_55),
.A2(n_63),
.B(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_55),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_55),
.A2(n_128),
.B(n_188),
.Y(n_187)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_60),
.B1(n_77),
.B2(n_78),
.Y(n_80)
);

AOI32xp33_ASAP7_75t_L g154 ( 
.A1(n_59),
.A2(n_70),
.A3(n_78),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_SL g156 ( 
.A(n_60),
.B(n_77),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_60),
.B(n_208),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_74),
.B(n_81),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_68),
.A2(n_75),
.B1(n_80),
.B2(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_71),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_73),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_75),
.A2(n_82),
.B(n_179),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_79),
.A2(n_109),
.B(n_111),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_79),
.A2(n_111),
.B(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_98),
.B2(n_99),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_92),
.B(n_97),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_92),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_93),
.A2(n_232),
.B(n_233),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_93),
.A2(n_233),
.B(n_251),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_105),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_101),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_101),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_101),
.A2(n_103),
.B1(n_104),
.B2(n_106),
.Y(n_118)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_102),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_102),
.B(n_183),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.C(n_119),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_118),
.Y(n_164)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_126),
.C(n_131),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_121),
.B(n_124),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_158),
.B1(n_159),
.B2(n_161),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_127),
.B1(n_131),
.B2(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_129),
.B(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_130),
.A2(n_150),
.B1(n_152),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_132),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_165),
.B(n_293),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_163),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_138),
.B(n_163),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.C(n_145),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_139),
.A2(n_140),
.B1(n_143),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_143),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_145),
.B(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.C(n_153),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_148),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_153),
.B(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_157),
.Y(n_185)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_162),
.A2(n_258),
.B(n_266),
.Y(n_265)
);

O2A1O1Ixp33_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_200),
.B(n_287),
.C(n_292),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_194),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_194),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_185),
.C(n_186),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_168),
.A2(n_169),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_178),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_174),
.C(n_178),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_173),
.Y(n_188)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_183),
.B(n_184),
.Y(n_179)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_185),
.B(n_186),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.C(n_191),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_227),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_191),
.Y(n_227)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_195),
.B(n_198),
.C(n_199),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_281),
.B(n_286),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_234),
.B(n_280),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_223),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_205),
.B(n_223),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_216),
.C(n_220),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_206),
.B(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_209),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B(n_214),
.Y(n_209)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_216),
.A2(n_220),
.B1(n_221),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_216),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_219),
.Y(n_232)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_228),
.B2(n_229),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_224),
.B(n_230),
.C(n_231),
.Y(n_285)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_274),
.B(n_279),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_254),
.B(n_273),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_248),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_248),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_243),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_239),
.B(n_242),
.C(n_243),
.Y(n_278)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_252),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_249),
.A2(n_250),
.B1(n_252),
.B2(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_262),
.B(n_272),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_260),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_260),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_267),
.B(n_271),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_265),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_270),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_278),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_278),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_285),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_285),
.Y(n_286)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_289),
.Y(n_292)
);


endmodule