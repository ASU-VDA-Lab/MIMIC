module fake_jpeg_12868_n_118 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_118);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_25),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_6),
.B(n_18),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_2),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_54),
.B(n_57),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_17),
.B1(n_37),
.B2(n_36),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_59),
.B1(n_52),
.B2(n_50),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_0),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_49),
.B(n_46),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_61),
.B(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_49),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_63),
.B(n_66),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_47),
.B1(n_50),
.B2(n_48),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_56),
.B1(n_46),
.B2(n_19),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_67),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_39),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_71),
.B(n_72),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_51),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_73),
.A2(n_23),
.B1(n_34),
.B2(n_33),
.Y(n_86)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_85),
.B1(n_87),
.B2(n_13),
.Y(n_101)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_14),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_82),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_15),
.C(n_35),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_1),
.B(n_3),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_89),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_74),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_79),
.B(n_88),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_62),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_86),
.A2(n_8),
.B(n_9),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_21),
.B1(n_30),
.B2(n_27),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_38),
.C(n_26),
.Y(n_88)
);

XNOR2x2_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_24),
.Y(n_91)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_98),
.C(n_84),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_86),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_92),
.A2(n_101),
.B1(n_104),
.B2(n_102),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_99),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_10),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_94),
.B(n_97),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_13),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_81),
.A2(n_11),
.B(n_12),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_90),
.B(n_11),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_100),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_107),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_108),
.A2(n_92),
.B1(n_98),
.B2(n_96),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_95),
.C(n_104),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_110),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_107),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_110),
.C(n_113),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_113),
.B1(n_111),
.B2(n_109),
.Y(n_116)
);

BUFx24_ASAP7_75t_SL g117 ( 
.A(n_116),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_106),
.B1(n_103),
.B2(n_101),
.Y(n_118)
);


endmodule