module real_jpeg_16961_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_518),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_0),
.B(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_1),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_1),
.B(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_1),
.A2(n_14),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

AND2x2_ASAP7_75t_SL g314 ( 
.A(n_1),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_1),
.B(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_1),
.B(n_467),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_1),
.B(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_2),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_3),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_3),
.Y(n_286)
);

BUFx5_ASAP7_75t_L g424 ( 
.A(n_3),
.Y(n_424)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_3),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_4),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_4),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_4),
.B(n_74),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_4),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_4),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_4),
.B(n_122),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_4),
.B(n_192),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_4),
.B(n_246),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_5),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_5),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_5),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_5),
.B(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_5),
.B(n_137),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_5),
.B(n_142),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_5),
.B(n_145),
.Y(n_144)
);

NAND2x1p5_ASAP7_75t_L g154 ( 
.A(n_5),
.B(n_105),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_6),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_6),
.B(n_205),
.Y(n_204)
);

AND2x2_ASAP7_75t_SL g276 ( 
.A(n_6),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_6),
.B(n_105),
.Y(n_287)
);

AND2x2_ASAP7_75t_SL g317 ( 
.A(n_6),
.B(n_114),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_6),
.B(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_6),
.B(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_6),
.B(n_312),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_7),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_7),
.B(n_354),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_7),
.B(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_7),
.B(n_445),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_7),
.B(n_479),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_7),
.B(n_500),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_7),
.B(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_8),
.B(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_8),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_8),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_8),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_8),
.B(n_311),
.Y(n_310)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_9),
.Y(n_142)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_9),
.Y(n_247)
);

BUFx5_ASAP7_75t_L g312 ( 
.A(n_9),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_10),
.Y(n_93)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_10),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_10),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_10),
.Y(n_383)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_11),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_12),
.Y(n_79)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_12),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g228 ( 
.A(n_12),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_13),
.B(n_45),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_13),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_13),
.B(n_348),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_13),
.B(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_13),
.B(n_440),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_13),
.B(n_30),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_13),
.B(n_490),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_13),
.B(n_492),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_14),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_14),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_14),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_14),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_14),
.B(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_14),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_14),
.B(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_14),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_15),
.Y(n_106)
);

BUFx4f_ASAP7_75t_L g102 ( 
.A(n_16),
.Y(n_102)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_16),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_16),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g275 ( 
.A(n_16),
.Y(n_275)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_17),
.Y(n_145)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_17),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_168),
.Y(n_19)
);

NAND2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_167),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_146),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_23),
.B(n_146),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_80),
.C(n_107),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_24),
.B(n_80),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_54),
.B2(n_55),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_41),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_27),
.B(n_41),
.C(n_54),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_33),
.C(n_38),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_28),
.A2(n_29),
.B1(n_38),
.B2(n_52),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_28),
.A2(n_29),
.B1(n_98),
.B2(n_99),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_28),
.A2(n_29),
.B1(n_314),
.B2(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_29),
.B(n_98),
.C(n_103),
.Y(n_97)
);

MAJx2_ASAP7_75t_L g313 ( 
.A(n_29),
.B(n_314),
.C(n_317),
.Y(n_313)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_33),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_34),
.B(n_104),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_37),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_38),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_38),
.B(n_121),
.C(n_289),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_38),
.A2(n_52),
.B1(n_120),
.B2(n_121),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_46),
.Y(n_41)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_42),
.Y(n_162)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_45),
.Y(n_189)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_47),
.A2(n_53),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_47),
.B(n_52),
.C(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_47),
.A2(n_53),
.B1(n_225),
.B2(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_53),
.B(n_127),
.C(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_71),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_56),
.B(n_72),
.C(n_76),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_63),
.C(n_67),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_57),
.A2(n_58),
.B1(n_67),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_60),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_61),
.Y(n_267)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_62),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_63),
.A2(n_129),
.B1(n_130),
.B2(n_132),
.Y(n_128)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g198 ( 
.A(n_67),
.B(n_199),
.C(n_202),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_67),
.B(n_202),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_69),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_70),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_71)
);

MAJx2_ASAP7_75t_L g197 ( 
.A(n_72),
.B(n_198),
.C(n_204),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_72),
.A2(n_73),
.B1(n_204),
.B2(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_73),
.B(n_134),
.C(n_143),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_73),
.B(n_144),
.Y(n_208)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_78),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_79),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_83),
.C(n_97),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_81),
.B(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_83),
.B(n_97),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_90),
.C(n_94),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_84),
.A2(n_85),
.B1(n_90),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_90),
.A2(n_127),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_93),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_94),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_98),
.A2(n_99),
.B1(n_140),
.B2(n_141),
.Y(n_185)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_136),
.C(n_140),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_99),
.B(n_245),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_99),
.B(n_261),
.Y(n_418)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_103),
.B(n_110),
.Y(n_109)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_106),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_107),
.B(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_128),
.C(n_133),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_108),
.B(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.C(n_125),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_109),
.B(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_111),
.B(n_125),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_117),
.C(n_120),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_112),
.A2(n_113),
.B1(n_117),
.B2(n_118),
.Y(n_196)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_L g446 ( 
.A(n_119),
.Y(n_446)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_121),
.B(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_124),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_128),
.B(n_133),
.Y(n_178)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AO22x1_ASAP7_75t_SL g207 ( 
.A1(n_134),
.A2(n_135),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_187),
.C(n_190),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_140),
.A2(n_141),
.B1(n_190),
.B2(n_191),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_140),
.B(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_141),
.B(n_426),
.Y(n_470)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_142),
.Y(n_493)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_165),
.B2(n_166),
.Y(n_148)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_155),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_153),
.B(n_238),
.C(n_248),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_153),
.A2(n_154),
.B1(n_248),
.B2(n_249),
.Y(n_296)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_161),
.B1(n_163),
.B2(n_164),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_156),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_159),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_251),
.B(n_515),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_210),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_173),
.A2(n_516),
.B(n_517),
.Y(n_515)
);

NOR2xp67_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_174),
.B(n_176),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.C(n_181),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_179),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_212),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_197),
.C(n_207),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_182),
.A2(n_183),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.C(n_195),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_184),
.B(n_337),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_186),
.B(n_195),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_187),
.B(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_188),
.B(n_358),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_188),
.B(n_382),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_190),
.A2(n_191),
.B1(n_309),
.B2(n_310),
.Y(n_376)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_191),
.B(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_197),
.B(n_207),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_234),
.Y(n_233)
);

XNOR2x2_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_204),
.Y(n_235)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_208),
.Y(n_209)
);

OR2x6_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_211),
.B(n_213),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.C(n_219),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_214),
.B(n_217),
.Y(n_404)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_215),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_219),
.B(n_404),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_232),
.C(n_236),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_220),
.A2(n_221),
.B1(n_333),
.B2(n_335),
.Y(n_332)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.C(n_229),
.Y(n_221)
);

XNOR2x1_ASAP7_75t_L g300 ( 
.A(n_222),
.B(n_301),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_224),
.A2(n_229),
.B1(n_230),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_224),
.Y(n_302)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_225),
.Y(n_322)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_233),
.A2(n_236),
.B1(n_237),
.B2(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_233),
.Y(n_334)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_238),
.A2(n_239),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_244),
.C(n_245),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_240),
.A2(n_245),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_243),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_245),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_246),
.Y(n_365)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

NAND2x1_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_406),
.Y(n_251)
);

A2O1A1O1Ixp25_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_340),
.B(n_399),
.C(n_400),
.D(n_405),
.Y(n_252)
);

NAND4xp25_ASAP7_75t_L g406 ( 
.A(n_253),
.B(n_400),
.C(n_407),
.D(n_409),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_326),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_254),
.B(n_326),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_299),
.C(n_303),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_255),
.A2(n_256),
.B1(n_300),
.B2(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_283),
.Y(n_256)
);

INVxp33_ASAP7_75t_SL g328 ( 
.A(n_257),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_262),
.C(n_268),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_258),
.B(n_391),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_262),
.A2(n_263),
.B1(n_268),
.B2(n_269),
.Y(n_391)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_263),
.A2(n_357),
.B(n_362),
.Y(n_356)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_276),
.C(n_280),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_270),
.B(n_280),
.Y(n_306)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_275),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_275),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_306),
.Y(n_305)
);

INVx8_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_294),
.B1(n_297),
.B2(n_298),
.Y(n_283)
);

INVxp67_ASAP7_75t_SL g297 ( 
.A(n_284),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_284),
.Y(n_329)
);

A2O1A1Ixp33_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_287),
.B(n_288),
.C(n_291),
.Y(n_284)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_285),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_285),
.A2(n_287),
.B1(n_292),
.B2(n_293),
.Y(n_325)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_287),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_325),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_289),
.B(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_294),
.Y(n_298)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_298),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_300),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_303),
.B(n_396),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_318),
.C(n_323),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_304),
.B(n_388),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_307),
.C(n_313),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_305),
.B(n_370),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_307),
.A2(n_308),
.B1(n_313),
.B2(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

BUFx12f_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_313),
.Y(n_371)
);

CKINVDCx14_ASAP7_75t_R g375 ( 
.A(n_314),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g373 ( 
.A(n_317),
.B(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_319),
.B(n_324),
.Y(n_388)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_331),
.Y(n_326)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_327),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.C(n_330),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_332),
.A2(n_336),
.B1(n_338),
.B2(n_339),
.Y(n_331)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_332),
.Y(n_338)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_333),
.Y(n_335)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_336),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_336),
.B(n_338),
.C(n_402),
.Y(n_401)
);

OAI21x1_ASAP7_75t_SL g340 ( 
.A1(n_341),
.A2(n_393),
.B(n_398),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_386),
.Y(n_341)
);

NOR2x1_ASAP7_75t_L g408 ( 
.A(n_342),
.B(n_386),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_368),
.C(n_372),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_343),
.B(n_430),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_355),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_344),
.B(n_356),
.C(n_366),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.C(n_352),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_345),
.B(n_416),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_346),
.A2(n_347),
.B1(n_352),
.B2(n_353),
.Y(n_416)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_366),
.Y(n_355)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_368),
.A2(n_369),
.B1(n_372),
.B2(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_372),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_376),
.C(n_377),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_373),
.B(n_414),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_376),
.B(n_377),
.Y(n_414)
);

MAJx2_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.C(n_384),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_378),
.B(n_384),
.Y(n_452)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_381),
.B(n_452),
.Y(n_451)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_383),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_389),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_387),
.B(n_390),
.C(n_392),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_392),
.Y(n_389)
);

NOR2x1_ASAP7_75t_L g407 ( 
.A(n_393),
.B(n_408),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_395),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g398 ( 
.A(n_394),
.B(n_395),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_403),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_401),
.B(n_403),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_410),
.A2(n_432),
.B(n_514),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_429),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_411),
.B(n_429),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_415),
.C(n_417),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_412),
.A2(n_413),
.B1(n_454),
.B2(n_455),
.Y(n_453)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g455 ( 
.A(n_415),
.B(n_417),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_419),
.C(n_425),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_418),
.A2(n_419),
.B1(n_420),
.B2(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_418),
.Y(n_437)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_423),
.Y(n_502)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_425),
.B(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_427),
.Y(n_507)
);

INVx5_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

AOI21x1_ASAP7_75t_SL g432 ( 
.A1(n_433),
.A2(n_456),
.B(n_513),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_453),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_434),
.B(n_453),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_438),
.C(n_451),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_435),
.B(n_472),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_438),
.B(n_451),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_444),
.C(n_447),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_439),
.B(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_447),
.Y(n_461)
);

INVx5_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

OAI21x1_ASAP7_75t_L g456 ( 
.A1(n_457),
.A2(n_473),
.B(n_512),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_471),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_458),
.B(n_471),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_462),
.C(n_469),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_SL g482 ( 
.A1(n_459),
.A2(n_460),
.B1(n_483),
.B2(n_485),
.Y(n_482)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_462),
.A2(n_469),
.B1(n_470),
.B2(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_462),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_465),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_463),
.A2(n_464),
.B1(n_465),
.B2(n_466),
.Y(n_476)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_474),
.A2(n_486),
.B(n_511),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_482),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_475),
.B(n_482),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.C(n_481),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_476),
.B(n_495),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_477),
.A2(n_478),
.B1(n_481),
.B2(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_481),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_483),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_487),
.A2(n_497),
.B(n_510),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_494),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_488),
.B(n_494),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_491),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_489),
.B(n_491),
.Y(n_503)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_498),
.A2(n_504),
.B(n_509),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_503),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_499),
.B(n_503),
.Y(n_509)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_508),
.Y(n_504)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);


endmodule