module fake_jpeg_15063_n_38 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_38);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_38;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

INVx5_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx4_ASAP7_75t_SL g15 ( 
.A(n_10),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

OA22x2_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_19),
.A2(n_20),
.B1(n_22),
.B2(n_15),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_17),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_15),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_22)
);

NAND3xp33_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_16),
.C(n_6),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_16),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_18),
.Y(n_27)
);

AOI322xp5_ASAP7_75t_L g28 ( 
.A1(n_27),
.A2(n_19),
.A3(n_15),
.B1(n_17),
.B2(n_18),
.C1(n_21),
.C2(n_5),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_29),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_5),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_25),
.B(n_24),
.Y(n_32)
);

NOR2xp67_ASAP7_75t_SL g35 ( 
.A(n_32),
.B(n_34),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_10),
.Y(n_34)
);

AOI322xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_31),
.C2(n_30),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_35),
.B1(n_33),
.B2(n_8),
.Y(n_38)
);


endmodule