module fake_jpeg_462_n_311 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_311);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_8),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_21),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_46),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_21),
.B(n_0),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_23),
.B(n_1),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_50),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_23),
.B(n_1),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_24),
.B(n_3),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_53),
.Y(n_90)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_52),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_24),
.B(n_3),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_60),
.Y(n_130)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_28),
.B(n_4),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_68),
.Y(n_95)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_73),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_72),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_28),
.B(n_5),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_75),
.Y(n_98)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_78),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_29),
.B(n_5),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_77),
.B(n_39),
.Y(n_103)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_81),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_82),
.Y(n_113)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_29),
.B(n_5),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_26),
.Y(n_83)
);

NOR2x1_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_47),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_85),
.Y(n_116)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_37),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_31),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_63),
.A2(n_26),
.B1(n_18),
.B2(n_36),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_91),
.A2(n_110),
.B1(n_120),
.B2(n_133),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_117),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_103),
.B(n_88),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_83),
.A2(n_37),
.B1(n_42),
.B2(n_40),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_107),
.A2(n_114),
.B1(n_124),
.B2(n_131),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_60),
.A2(n_18),
.B1(n_31),
.B2(n_36),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_112),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_48),
.A2(n_55),
.B1(n_86),
.B2(n_56),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_57),
.B(n_44),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_118),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_54),
.A2(n_36),
.B1(n_43),
.B2(n_33),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_66),
.B(n_39),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_128),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_58),
.A2(n_27),
.B1(n_43),
.B2(n_38),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_84),
.A2(n_25),
.B1(n_38),
.B2(n_33),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_125),
.A2(n_98),
.B(n_113),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_67),
.B(n_42),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_59),
.B(n_44),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_7),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_62),
.A2(n_27),
.B1(n_40),
.B2(n_17),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_71),
.B(n_6),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_135),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_78),
.A2(n_70),
.B1(n_87),
.B2(n_72),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_87),
.A2(n_17),
.B1(n_30),
.B2(n_9),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_134),
.A2(n_137),
.B1(n_139),
.B2(n_124),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_61),
.B(n_6),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_79),
.B(n_7),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_130),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_75),
.A2(n_30),
.B1(n_9),
.B2(n_10),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_48),
.A2(n_30),
.B1(n_13),
.B2(n_15),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_138),
.A2(n_117),
.B1(n_129),
.B2(n_125),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_141),
.B(n_176),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_131),
.A2(n_30),
.B1(n_13),
.B2(n_15),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_142),
.A2(n_159),
.B1(n_181),
.B2(n_144),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_15),
.B(n_89),
.C(n_90),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_143),
.B(n_146),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_145),
.A2(n_156),
.B1(n_162),
.B2(n_170),
.Y(n_190)
);

NOR2x1_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_95),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_154),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_152),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_102),
.B(n_94),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_173),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_109),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_155),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_94),
.A2(n_138),
.B1(n_126),
.B2(n_92),
.Y(n_156)
);

NAND2xp33_ASAP7_75t_SL g213 ( 
.A(n_157),
.B(n_165),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_126),
.A2(n_108),
.B1(n_121),
.B2(n_119),
.Y(n_159)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_103),
.A2(n_97),
.B1(n_116),
.B2(n_121),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_96),
.B(n_106),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_166),
.Y(n_201)
);

AND2x4_ASAP7_75t_L g165 ( 
.A(n_106),
.B(n_101),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_97),
.A2(n_105),
.B1(n_108),
.B2(n_121),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_105),
.Y(n_171)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_111),
.B(n_127),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_115),
.Y(n_174)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_111),
.B(n_127),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_179),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_123),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_115),
.Y(n_177)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_108),
.B(n_119),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_119),
.B(n_104),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_183),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_L g181 ( 
.A1(n_99),
.A2(n_126),
.B1(n_102),
.B2(n_91),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_104),
.A2(n_99),
.B1(n_130),
.B2(n_117),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_182),
.A2(n_149),
.B1(n_156),
.B2(n_172),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_104),
.B(n_117),
.Y(n_183)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_140),
.A2(n_104),
.A3(n_153),
.B1(n_141),
.B2(n_183),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_192),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_140),
.B(n_145),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_194),
.A2(n_181),
.B1(n_180),
.B2(n_179),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_173),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_204),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_199),
.A2(n_178),
.B1(n_171),
.B2(n_151),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_169),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_157),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_161),
.C(n_163),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_150),
.B(n_147),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_152),
.B(n_176),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_165),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_165),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_158),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_192),
.B(n_184),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_214),
.B(n_223),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_221),
.A2(n_234),
.B(n_237),
.Y(n_254)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_184),
.B(n_143),
.Y(n_223)
);

NOR3xp33_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_165),
.C(n_177),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_203),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_227),
.Y(n_251)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_226),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_203),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_202),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_187),
.B(n_185),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_230),
.B(n_197),
.Y(n_246)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_231),
.B(n_232),
.Y(n_239)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_188),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_174),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_205),
.B(n_202),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_190),
.A2(n_194),
.B1(n_187),
.B2(n_185),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_236),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_190),
.A2(n_204),
.B1(n_209),
.B2(n_189),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_209),
.A2(n_193),
.B(n_196),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_201),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_238),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_249),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_247),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_219),
.B(n_197),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_219),
.B(n_197),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_256),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_198),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_217),
.C(n_233),
.Y(n_259)
);

OAI32xp33_ASAP7_75t_L g256 ( 
.A1(n_216),
.A2(n_198),
.A3(n_199),
.B1(n_195),
.B2(n_186),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_228),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_257),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_261),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_216),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_240),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_264),
.Y(n_275)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_253),
.A2(n_214),
.B1(n_235),
.B2(n_236),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_268),
.B1(n_244),
.B2(n_254),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_229),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_267),
.C(n_272),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_233),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_253),
.A2(n_221),
.B1(n_234),
.B2(n_224),
.Y(n_268)
);

OAI321xp33_ASAP7_75t_L g269 ( 
.A1(n_241),
.A2(n_223),
.A3(n_237),
.B1(n_218),
.B2(n_215),
.C(n_225),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_269),
.B(n_270),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_242),
.B(n_227),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_232),
.C(n_231),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_258),
.A2(n_245),
.B1(n_256),
.B2(n_248),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_273),
.A2(n_283),
.B1(n_265),
.B2(n_268),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_246),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_262),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_271),
.A2(n_242),
.B(n_257),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_278),
.A2(n_258),
.B(n_254),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_260),
.B(n_241),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_279),
.B(n_281),
.Y(n_284)
);

BUFx24_ASAP7_75t_SL g281 ( 
.A(n_261),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_251),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_267),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_291),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_287),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_266),
.C(n_259),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_292),
.C(n_285),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_280),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_275),
.A2(n_250),
.B1(n_252),
.B2(n_239),
.Y(n_290)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_290),
.Y(n_298)
);

O2A1O1Ixp33_ASAP7_75t_L g291 ( 
.A1(n_273),
.A2(n_250),
.B(n_220),
.C(n_226),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_239),
.C(n_222),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_291),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_297),
.C(n_287),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_280),
.C(n_277),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_292),
.Y(n_299)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_299),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_274),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_301),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_284),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_302),
.A2(n_303),
.B(n_293),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_299),
.B(n_293),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_307),
.A2(n_308),
.B(n_304),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_252),
.C(n_206),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_309),
.B(n_310),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_307),
.A2(n_252),
.B(n_200),
.Y(n_310)
);


endmodule