module fake_jpeg_1359_n_28 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_28);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_28;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_15;

INVx2_ASAP7_75t_SL g9 ( 
.A(n_6),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_3),
.Y(n_12)
);

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_15),
.B(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_16),
.B1(n_10),
.B2(n_9),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_20),
.A2(n_10),
.B1(n_12),
.B2(n_4),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_1),
.B(n_3),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_19),
.C(n_20),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_23),
.A2(n_24),
.B1(n_22),
.B2(n_4),
.Y(n_25)
);

AOI21x1_ASAP7_75t_L g26 ( 
.A1(n_25),
.A2(n_5),
.B(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

BUFx24_ASAP7_75t_SL g28 ( 
.A(n_27),
.Y(n_28)
);


endmodule