module fake_netlist_1_1348_n_38 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_38);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
INVx1_ASAP7_75t_L g11 ( .A(n_5), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_6), .Y(n_12) );
CKINVDCx20_ASAP7_75t_R g13 ( .A(n_1), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_3), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_2), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_8), .Y(n_16) );
BUFx6f_ASAP7_75t_L g17 ( .A(n_5), .Y(n_17) );
NOR2xp33_ASAP7_75t_R g18 ( .A(n_15), .B(n_10), .Y(n_18) );
INVx4_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_12), .B(n_0), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_11), .B(n_0), .Y(n_21) );
NAND3xp33_ASAP7_75t_SL g22 ( .A(n_14), .B(n_1), .C(n_2), .Y(n_22) );
INVx4_ASAP7_75t_L g23 ( .A(n_19), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_19), .B(n_16), .Y(n_24) );
A2O1A1Ixp33_ASAP7_75t_L g25 ( .A1(n_21), .A2(n_17), .B(n_13), .C(n_4), .Y(n_25) );
AOI22xp33_ASAP7_75t_L g26 ( .A1(n_22), .A2(n_17), .B1(n_13), .B2(n_4), .Y(n_26) );
OR2x2_ASAP7_75t_L g27 ( .A(n_25), .B(n_20), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_23), .Y(n_28) );
HB1xp67_ASAP7_75t_L g29 ( .A(n_24), .Y(n_29) );
OAI211xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_26), .B(n_18), .C(n_23), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_31), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_30), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
NAND2xp5_ASAP7_75t_L g35 ( .A(n_33), .B(n_27), .Y(n_35) );
CKINVDCx5p33_ASAP7_75t_R g36 ( .A(n_34), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_36), .Y(n_37) );
AOI322xp5_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_17), .A3(n_35), .B1(n_34), .B2(n_3), .C1(n_9), .C2(n_7), .Y(n_38) );
endmodule