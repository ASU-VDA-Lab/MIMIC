module fake_jpeg_13656_n_531 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_531);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_531;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_17),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_17),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_2),
.A2(n_4),
.B(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_19),
.B(n_18),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_51),
.B(n_73),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_52),
.Y(n_131)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_54),
.Y(n_137)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_55),
.Y(n_138)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_56),
.Y(n_155)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_60),
.B(n_71),
.Y(n_110)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_65),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_29),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_66),
.B(n_102),
.Y(n_116)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_69),
.Y(n_161)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_23),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_72),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_19),
.B(n_18),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_74),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_30),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

BUFx4f_ASAP7_75t_SL g76 ( 
.A(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_76),
.B(n_79),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_77),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_44),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_80),
.B(n_83),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_20),
.B(n_16),
.Y(n_83)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_84),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_92),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_21),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_90),
.B(n_94),
.Y(n_133)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_93),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_39),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

NAND2xp33_ASAP7_75t_SL g159 ( 
.A(n_95),
.B(n_96),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

AOI21xp33_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_31),
.B(n_32),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_100),
.Y(n_135)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_27),
.Y(n_104)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_101),
.B(n_44),
.Y(n_147)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_59),
.A2(n_36),
.B1(n_49),
.B2(n_24),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g163 ( 
.A1(n_103),
.A2(n_35),
.B1(n_89),
.B2(n_95),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_84),
.A2(n_50),
.B1(n_48),
.B2(n_31),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_107),
.A2(n_112),
.B1(n_124),
.B2(n_132),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_66),
.B(n_28),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_108),
.B(n_144),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_97),
.A2(n_50),
.B1(n_48),
.B2(n_31),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_57),
.B(n_40),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_122),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_61),
.B(n_40),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_123),
.B(n_156),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_82),
.A2(n_50),
.B1(n_48),
.B2(n_43),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_82),
.A2(n_50),
.B1(n_48),
.B2(n_43),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_90),
.A2(n_50),
.B1(n_43),
.B2(n_38),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_136),
.A2(n_139),
.B1(n_143),
.B2(n_72),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_90),
.A2(n_38),
.B1(n_32),
.B2(n_46),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_98),
.A2(n_38),
.B1(n_32),
.B2(n_46),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_98),
.B(n_20),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_96),
.A2(n_40),
.B1(n_28),
.B2(n_36),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_145),
.A2(n_151),
.B1(n_160),
.B2(n_1),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_76),
.B(n_44),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_42),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_70),
.A2(n_49),
.B1(n_24),
.B2(n_33),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_65),
.B(n_37),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_63),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_91),
.A2(n_37),
.B1(n_35),
.B2(n_33),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_163),
.A2(n_178),
.B1(n_187),
.B2(n_212),
.Y(n_237)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_164),
.Y(n_230)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_168),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_126),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_169),
.B(n_186),
.Y(n_234)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_170),
.Y(n_265)
);

O2A1O1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_117),
.A2(n_56),
.B(n_76),
.C(n_75),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_171),
.B(n_189),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_105),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_172),
.Y(n_248)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_173),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_174),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_151),
.A2(n_92),
.B1(n_93),
.B2(n_77),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_175),
.A2(n_196),
.B1(n_198),
.B2(n_208),
.Y(n_264)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_176),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_122),
.A2(n_69),
.B1(n_74),
.B2(n_58),
.Y(n_178)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_179),
.Y(n_244)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_181),
.Y(n_249)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_182),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_127),
.B(n_53),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_183),
.B(n_184),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_42),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_106),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_116),
.A2(n_62),
.B1(n_64),
.B2(n_81),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_120),
.Y(n_188)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_188),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_135),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_190),
.B(n_197),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_191),
.Y(n_245)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_192),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_133),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_193),
.B(n_200),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_108),
.B(n_102),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_194),
.B(n_199),
.Y(n_236)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_128),
.Y(n_195)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_195),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_118),
.A2(n_87),
.B1(n_158),
.B2(n_101),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_144),
.B(n_42),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_118),
.A2(n_68),
.B1(n_99),
.B2(n_67),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_106),
.Y(n_200)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_113),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_201),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_203),
.C(n_211),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_116),
.B(n_88),
.C(n_86),
.Y(n_203)
);

INVx11_ASAP7_75t_L g204 ( 
.A(n_155),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_204),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_138),
.A2(n_55),
.B1(n_54),
.B2(n_52),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_205),
.A2(n_138),
.B1(n_131),
.B2(n_137),
.Y(n_251)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_128),
.Y(n_206)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_206),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_110),
.B(n_42),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_213),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_118),
.A2(n_42),
.B1(n_85),
.B2(n_39),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_209),
.B(n_210),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_104),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_159),
.A2(n_1),
.B(n_3),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_159),
.A2(n_39),
.B1(n_16),
.B2(n_78),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_129),
.B(n_1),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_114),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_214),
.B(n_14),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_129),
.B(n_39),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_215),
.B(n_220),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_140),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_216),
.A2(n_162),
.B1(n_138),
.B2(n_161),
.Y(n_242)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_134),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_221),
.Y(n_238)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_134),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_218),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_219),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_142),
.B(n_146),
.C(n_125),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_114),
.B(n_3),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_165),
.A2(n_140),
.B1(n_148),
.B2(n_119),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_228),
.A2(n_229),
.B1(n_239),
.B2(n_246),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_219),
.A2(n_177),
.B1(n_180),
.B2(n_171),
.Y(n_229)
);

FAx1_ASAP7_75t_SL g232 ( 
.A(n_165),
.B(n_137),
.CI(n_131),
.CON(n_232),
.SN(n_232)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_232),
.B(n_243),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_210),
.A2(n_178),
.B1(n_177),
.B2(n_212),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_233),
.A2(n_242),
.B1(n_259),
.B2(n_269),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_199),
.A2(n_148),
.B1(n_119),
.B2(n_158),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_221),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_203),
.A2(n_119),
.B1(n_161),
.B2(n_111),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_202),
.B(n_213),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_215),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_251),
.Y(n_274)
);

FAx1_ASAP7_75t_SL g253 ( 
.A(n_202),
.B(n_142),
.CI(n_146),
.CON(n_253),
.SN(n_253)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_253),
.B(n_258),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_189),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_187),
.A2(n_111),
.B1(n_157),
.B2(n_130),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_167),
.A2(n_130),
.B1(n_121),
.B2(n_113),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_262),
.A2(n_266),
.B1(n_270),
.B2(n_272),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_180),
.A2(n_141),
.B1(n_125),
.B2(n_109),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_263),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_194),
.A2(n_130),
.B1(n_121),
.B2(n_113),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_211),
.A2(n_121),
.B1(n_109),
.B2(n_155),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_166),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_273),
.Y(n_321)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_250),
.Y(n_275)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_275),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_276),
.B(n_318),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_234),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_278),
.B(n_279),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_254),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_250),
.Y(n_280)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_280),
.Y(n_343)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_281),
.Y(n_326)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_256),
.Y(n_282)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_282),
.Y(n_330)
);

NAND2xp33_ASAP7_75t_SL g283 ( 
.A(n_267),
.B(n_190),
.Y(n_283)
);

OAI21xp33_ASAP7_75t_L g335 ( 
.A1(n_283),
.A2(n_304),
.B(n_308),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_226),
.B(n_166),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_284),
.B(n_300),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_243),
.B(n_238),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_285),
.B(n_295),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_273),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_286),
.B(n_309),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_267),
.A2(n_214),
.B(n_186),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_288),
.A2(n_293),
.B(n_298),
.Y(n_338)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_256),
.Y(n_289)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_289),
.Y(n_334)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_257),
.Y(n_291)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_291),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_267),
.A2(n_200),
.B(n_209),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_231),
.A2(n_169),
.B(n_207),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_294),
.A2(n_320),
.B(n_272),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_238),
.B(n_220),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_261),
.B(n_217),
.C(n_188),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_296),
.B(n_297),
.C(n_303),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_247),
.B(n_192),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_224),
.A2(n_204),
.B(n_173),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_257),
.Y(n_299)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_299),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_225),
.B(n_170),
.Y(n_300)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_249),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_302),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_231),
.B(n_195),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_271),
.B(n_218),
.Y(n_304)
);

AO22x1_ASAP7_75t_L g305 ( 
.A1(n_232),
.A2(n_206),
.B1(n_179),
.B2(n_185),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_305),
.A2(n_317),
.B(n_242),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_224),
.A2(n_191),
.B1(n_182),
.B2(n_181),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_306),
.A2(n_268),
.B1(n_245),
.B2(n_249),
.Y(n_362)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_260),
.Y(n_307)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_307),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_261),
.B(n_176),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_260),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_230),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_310),
.B(n_312),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_246),
.A2(n_236),
.B1(n_264),
.B2(n_228),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_311),
.A2(n_240),
.B1(n_244),
.B2(n_201),
.Y(n_353)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_230),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_222),
.B(n_168),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_314),
.B(n_315),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_222),
.B(n_216),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_232),
.B(n_164),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_316),
.B(n_253),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_239),
.B(n_191),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_240),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_241),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_241),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_269),
.A2(n_7),
.B(n_8),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_304),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_325),
.B(n_327),
.Y(n_370)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_304),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_294),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_328),
.B(n_360),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_337),
.B(n_354),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_340),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_341),
.B(n_346),
.Y(n_377)
);

INVx11_ASAP7_75t_L g342 ( 
.A(n_319),
.Y(n_342)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_342),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_285),
.B(n_286),
.Y(n_346)
);

INVx8_ASAP7_75t_L g347 ( 
.A(n_281),
.Y(n_347)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_347),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_303),
.B(n_236),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_349),
.B(n_359),
.C(n_299),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_350),
.B(n_298),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_301),
.A2(n_262),
.B1(n_266),
.B2(n_237),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_351),
.A2(n_352),
.B1(n_362),
.B2(n_274),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_315),
.A2(n_237),
.B1(n_259),
.B2(n_253),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_353),
.A2(n_361),
.B1(n_317),
.B2(n_280),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_313),
.B(n_314),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_305),
.A2(n_248),
.B(n_268),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_355),
.A2(n_357),
.B(n_293),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_316),
.B(n_227),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_295),
.B(n_249),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_358),
.B(n_363),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_308),
.B(n_248),
.C(n_235),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_277),
.B(n_255),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_311),
.A2(n_201),
.B1(n_245),
.B2(n_244),
.Y(n_361)
);

AND2x6_ASAP7_75t_L g363 ( 
.A(n_305),
.B(n_265),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_342),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_364),
.B(n_384),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_365),
.A2(n_378),
.B1(n_324),
.B2(n_330),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_351),
.A2(n_290),
.B1(n_287),
.B2(n_321),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_366),
.A2(n_367),
.B1(n_368),
.B2(n_372),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_352),
.A2(n_290),
.B1(n_287),
.B2(n_322),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_348),
.B(n_308),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_369),
.B(n_385),
.C(n_387),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_348),
.B(n_296),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_371),
.B(n_393),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_353),
.A2(n_274),
.B1(n_317),
.B2(n_292),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_338),
.A2(n_292),
.B(n_288),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_373),
.B(n_396),
.Y(n_409)
);

AOI21x1_ASAP7_75t_L g426 ( 
.A1(n_374),
.A2(n_375),
.B(n_394),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_331),
.A2(n_276),
.B1(n_280),
.B2(n_297),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_346),
.B(n_275),
.Y(n_380)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_380),
.Y(n_400)
);

AO21x1_ASAP7_75t_L g382 ( 
.A1(n_363),
.A2(n_320),
.B(n_318),
.Y(n_382)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_382),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_323),
.B(n_312),
.Y(n_383)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_383),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_361),
.A2(n_310),
.B1(n_309),
.B2(n_307),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_349),
.B(n_291),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_358),
.B(n_331),
.C(n_344),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_388),
.B(n_357),
.C(n_332),
.Y(n_412)
);

AOI22x1_ASAP7_75t_L g389 ( 
.A1(n_357),
.A2(n_350),
.B1(n_355),
.B2(n_337),
.Y(n_389)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_389),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_323),
.B(n_289),
.Y(n_390)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_390),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_325),
.A2(n_282),
.B1(n_302),
.B2(n_252),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_391),
.B(n_399),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_344),
.B(n_227),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_338),
.B(n_255),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_357),
.A2(n_235),
.B(n_223),
.Y(n_395)
);

NOR3xp33_ASAP7_75t_L g401 ( 
.A(n_395),
.B(n_345),
.C(n_322),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_340),
.A2(n_359),
.B(n_335),
.Y(n_396)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_345),
.Y(n_398)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_398),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_333),
.A2(n_252),
.B1(n_223),
.B2(n_9),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_401),
.B(n_428),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_381),
.B(n_333),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_403),
.B(n_413),
.Y(n_445)
);

AND2x6_ASAP7_75t_L g410 ( 
.A(n_379),
.B(n_357),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_410),
.A2(n_420),
.B1(n_382),
.B2(n_370),
.Y(n_436)
);

XOR2x2_ASAP7_75t_L g411 ( 
.A(n_369),
.B(n_332),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_411),
.B(n_416),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_385),
.C(n_371),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_386),
.B(n_356),
.Y(n_413)
);

NOR3xp33_ASAP7_75t_L g416 ( 
.A(n_377),
.B(n_356),
.C(n_339),
.Y(n_416)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_376),
.Y(n_418)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_418),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_377),
.B(n_324),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_419),
.B(n_429),
.Y(n_438)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_376),
.Y(n_421)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_421),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_380),
.B(n_339),
.Y(n_422)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_422),
.Y(n_443)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_398),
.Y(n_423)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_423),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_388),
.B(n_326),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_425),
.Y(n_448)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_383),
.Y(n_427)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_427),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_390),
.B(n_336),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_387),
.B(n_326),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_402),
.A2(n_397),
.B1(n_375),
.B2(n_394),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_432),
.A2(n_405),
.B1(n_399),
.B2(n_406),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_433),
.B(n_434),
.C(n_439),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_408),
.B(n_397),
.C(n_396),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_408),
.B(n_379),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_435),
.B(n_447),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_436),
.B(n_449),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_424),
.B(n_393),
.C(n_378),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_407),
.A2(n_375),
.B1(n_374),
.B2(n_394),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_440),
.A2(n_432),
.B1(n_452),
.B2(n_453),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_418),
.Y(n_442)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_442),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_422),
.B(n_364),
.Y(n_446)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_446),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_424),
.B(n_389),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_417),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_417),
.B(n_384),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_450),
.B(n_451),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_423),
.B(n_395),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_411),
.B(n_389),
.C(n_373),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_452),
.B(n_455),
.C(n_426),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_409),
.A2(n_382),
.B(n_372),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_453),
.A2(n_426),
.B(n_404),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_412),
.B(n_420),
.C(n_414),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_456),
.B(n_458),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_433),
.B(n_402),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_435),
.B(n_414),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_459),
.B(n_462),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_439),
.B(n_404),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_463),
.B(n_464),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_434),
.B(n_406),
.C(n_427),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_445),
.B(n_413),
.Y(n_465)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_465),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_466),
.A2(n_467),
.B1(n_444),
.B2(n_442),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_419),
.Y(n_468)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_468),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_448),
.B(n_415),
.C(n_400),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_469),
.B(n_473),
.C(n_474),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_447),
.B(n_415),
.C(n_400),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_440),
.B(n_428),
.C(n_421),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_431),
.B(n_405),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_475),
.B(n_476),
.Y(n_492)
);

BUFx24_ASAP7_75t_SL g476 ( 
.A(n_437),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_446),
.Y(n_481)
);

OAI321xp33_ASAP7_75t_L g500 ( 
.A1(n_481),
.A2(n_483),
.A3(n_490),
.B1(n_484),
.B2(n_334),
.C(n_477),
.Y(n_500)
);

OAI321xp33_ASAP7_75t_L g483 ( 
.A1(n_472),
.A2(n_437),
.A3(n_454),
.B1(n_443),
.B2(n_450),
.C(n_451),
.Y(n_483)
);

NOR3xp33_ASAP7_75t_SL g484 ( 
.A(n_461),
.B(n_454),
.C(n_443),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_484),
.A2(n_367),
.B1(n_343),
.B2(n_329),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_474),
.A2(n_410),
.B(n_438),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_485),
.A2(n_489),
.B(n_460),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_486),
.B(n_463),
.Y(n_495)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_469),
.Y(n_487)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_487),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_464),
.B(n_444),
.C(n_441),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_488),
.B(n_343),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_473),
.A2(n_441),
.B(n_430),
.Y(n_489)
);

OAI321xp33_ASAP7_75t_L g490 ( 
.A1(n_471),
.A2(n_430),
.A3(n_336),
.B1(n_334),
.B2(n_330),
.C(n_392),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_482),
.A2(n_462),
.B1(n_460),
.B2(n_459),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_493),
.B(n_495),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_494),
.A2(n_485),
.B(n_489),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_457),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_501),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_480),
.B(n_458),
.C(n_392),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_498),
.B(n_504),
.C(n_505),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_481),
.Y(n_499)
);

AOI31xp67_ASAP7_75t_L g514 ( 
.A1(n_499),
.A2(n_500),
.A3(n_503),
.B(n_506),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_479),
.B(n_347),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_502),
.B(n_497),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_480),
.B(n_329),
.C(n_252),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_478),
.B(n_347),
.C(n_8),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_492),
.B(n_7),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_508),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_522)
);

AOI221xp5_ASAP7_75t_L g509 ( 
.A1(n_496),
.A2(n_494),
.B1(n_486),
.B2(n_502),
.C(n_495),
.Y(n_509)
);

NAND3xp33_ASAP7_75t_L g521 ( 
.A(n_509),
.B(n_510),
.C(n_511),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_496),
.A2(n_488),
.B(n_491),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_510),
.A2(n_513),
.B(n_509),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_512),
.B(n_515),
.Y(n_520)
);

AOI322xp5_ASAP7_75t_L g515 ( 
.A1(n_504),
.A2(n_491),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_7),
.C2(n_13),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_498),
.B(n_14),
.C(n_10),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_516),
.Y(n_519)
);

A2O1A1Ixp33_ASAP7_75t_L g517 ( 
.A1(n_514),
.A2(n_493),
.B(n_505),
.C(n_11),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_517),
.A2(n_518),
.B(n_516),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_521),
.B(n_10),
.Y(n_526)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_522),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_523),
.A2(n_524),
.B(n_526),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_520),
.A2(n_507),
.B(n_13),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_525),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_528),
.B(n_519),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_527),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_530),
.B(n_14),
.Y(n_531)
);


endmodule