module real_jpeg_16179_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx3_ASAP7_75t_L g94 ( 
.A(n_0),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_0),
.Y(n_101)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_0),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_1),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_1),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_1),
.A2(n_118),
.B1(n_310),
.B2(n_314),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_1),
.A2(n_118),
.B1(n_321),
.B2(n_323),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_2),
.A2(n_127),
.B1(n_132),
.B2(n_133),
.Y(n_126)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_2),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_2),
.A2(n_132),
.B1(n_187),
.B2(n_191),
.Y(n_186)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_3),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_3),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_3),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_3),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_4),
.A2(n_67),
.B1(n_71),
.B2(n_73),
.Y(n_66)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_5),
.A2(n_77),
.B1(n_82),
.B2(n_87),
.Y(n_76)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_5),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_5),
.A2(n_87),
.B1(n_212),
.B2(n_214),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_5),
.A2(n_87),
.B1(n_226),
.B2(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_5),
.A2(n_87),
.B1(n_251),
.B2(n_346),
.Y(n_345)
);

OAI22xp33_ASAP7_75t_L g196 ( 
.A1(n_6),
.A2(n_43),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_6),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_6),
.A2(n_197),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_6),
.A2(n_197),
.B1(n_296),
.B2(n_299),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_7),
.Y(n_330)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_8),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_8),
.Y(n_114)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_8),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_8),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_8),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_8),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_8),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_9),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_10),
.A2(n_177),
.B1(n_180),
.B2(n_183),
.Y(n_176)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_10),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_10),
.A2(n_183),
.B1(n_246),
.B2(n_251),
.Y(n_245)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_11),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_11),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_11),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_12),
.B(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_12),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_12),
.A2(n_34),
.B(n_208),
.Y(n_207)
);

OAI32xp33_ASAP7_75t_L g231 ( 
.A1(n_12),
.A2(n_232),
.A3(n_236),
.B1(n_239),
.B2(n_242),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_12),
.B(n_306),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_12),
.A2(n_48),
.B1(n_345),
.B2(n_348),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_12),
.A2(n_141),
.B1(n_369),
.B2(n_373),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_13),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g161 ( 
.A(n_14),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g206 ( 
.A(n_15),
.Y(n_206)
);

BUFx8_ASAP7_75t_L g210 ( 
.A(n_15),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_258),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_256),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_217),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_19),
.B(n_217),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_148),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_74),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_47),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_33),
.B1(n_37),
.B2(n_43),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_32),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AO21x2_ASAP7_75t_L g200 ( 
.A1(n_37),
.A2(n_143),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_39),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_40),
.Y(n_216)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_54),
.B1(n_65),
.B2(n_66),
.Y(n_47)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_48),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_48),
.A2(n_65),
.B1(n_295),
.B2(n_303),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_48),
.A2(n_320),
.B1(n_345),
.B2(n_355),
.Y(n_354)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_50),
.Y(n_139)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_53),
.Y(n_135)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_53),
.Y(n_281)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_53),
.Y(n_298)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_53),
.Y(n_302)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_53),
.Y(n_325)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_53),
.Y(n_342)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_55),
.A2(n_125),
.B1(n_126),
.B2(n_136),
.Y(n_124)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_63),
.Y(n_158)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_65),
.Y(n_255)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_69),
.Y(n_254)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_69),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_123),
.C(n_140),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_75),
.B(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_88),
.B1(n_115),
.B2(n_122),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_76),
.A2(n_88),
.B1(n_122),
.B2(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_82),
.Y(n_198)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AO22x2_ASAP7_75t_L g143 ( 
.A1(n_85),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_143)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_86),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_88),
.A2(n_115),
.B1(n_122),
.B2(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

OA21x2_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_98),
.B(n_105),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_97),
.Y(n_235)
);

INVxp33_ASAP7_75t_L g242 ( 
.A(n_98),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_106),
.B1(n_109),
.B2(n_112),
.Y(n_105)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_111),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_112),
.Y(n_225)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_114),
.Y(n_267)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_121),
.Y(n_377)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_122),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_123),
.A2(n_124),
.B1(n_140),
.B2(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_125),
.A2(n_126),
.B1(n_245),
.B2(n_255),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_125),
.A2(n_319),
.B1(n_326),
.B2(n_331),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_140),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_141),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_141),
.B(n_273),
.Y(n_272)
);

OAI21xp33_ASAP7_75t_SL g284 ( 
.A1(n_141),
.A2(n_272),
.B(n_285),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_141),
.B(n_327),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_141),
.B(n_184),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_142),
.A2(n_200),
.B1(n_207),
.B2(n_211),
.Y(n_199)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_199),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_194),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_176),
.B1(n_184),
.B2(n_185),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_151),
.A2(n_176),
.B1(n_184),
.B2(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_152),
.A2(n_284),
.B1(n_287),
.B2(n_292),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_152),
.A2(n_287),
.B1(n_292),
.B2(n_309),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_152),
.A2(n_224),
.B1(n_292),
.B2(n_309),
.Y(n_379)
);

AND2x2_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_164),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_157),
.B1(n_159),
.B2(n_162),
.Y(n_153)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_156),
.Y(n_280)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_160),
.Y(n_268)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_161),
.Y(n_250)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_161),
.Y(n_322)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_169),
.B1(n_172),
.B2(n_174),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_168),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_168),
.Y(n_313)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_173),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_175),
.Y(n_182)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_184),
.Y(n_292)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx8_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.C(n_229),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_218),
.A2(n_219),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_222),
.A2(n_229),
.B1(n_230),
.B2(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_222),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_243),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_231),
.A2(n_243),
.B1(n_244),
.B2(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_231),
.Y(n_364)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_241),
.Y(n_286)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_245),
.Y(n_303)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

OAI21x1_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_381),
.B(n_387),
.Y(n_258)
);

AOI21x1_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_360),
.B(n_380),
.Y(n_259)
);

OAI21x1_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_316),
.B(n_359),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_293),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_262),
.B(n_293),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_282),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_263),
.A2(n_282),
.B1(n_283),
.B2(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_263),
.Y(n_333)
);

OAI32xp33_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_268),
.A3(n_269),
.B1(n_272),
.B2(n_276),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_281),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_288),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_304),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_294),
.B(n_307),
.C(n_315),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_295),
.Y(n_331)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_307),
.B1(n_308),
.B2(n_315),
.Y(n_304)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_305),
.Y(n_315)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_334),
.B(n_358),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_332),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_318),
.B(n_332),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx6_ASAP7_75t_L g355 ( 
.A(n_329),
.Y(n_355)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_330),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_353),
.B(n_357),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_344),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_343),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_356),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_354),
.B(n_356),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

NOR2xp67_ASAP7_75t_SL g380 ( 
.A(n_361),
.B(n_362),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_365),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_363),
.B(n_366),
.C(n_379),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_366),
.A2(n_367),
.B1(n_378),
.B2(n_379),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_382),
.B(n_383),
.Y(n_387)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);


endmodule