module fake_jpeg_15542_n_262 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_262);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_262;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_152;
wire n_73;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_258;
wire n_96;

INVx11_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_11),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_2),
.B(n_10),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_39),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_40),
.B(n_46),
.Y(n_100)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_45),
.B(n_53),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_0),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_37),
.Y(n_49)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

HAxp5_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_1),
.CON(n_52),
.SN(n_52)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_21),
.B1(n_23),
.B2(n_22),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_28),
.B(n_1),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_1),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_26),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_58),
.A2(n_35),
.B1(n_30),
.B2(n_22),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_62),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_31),
.B(n_38),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_25),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_34),
.B1(n_26),
.B2(n_18),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_66),
.A2(n_76),
.B1(n_94),
.B2(n_4),
.Y(n_132)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_77),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_27),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_71),
.B(n_79),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_51),
.A2(n_34),
.B1(n_18),
.B2(n_16),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_27),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_27),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_80),
.B(n_81),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_38),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_84),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_31),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_39),
.B(n_32),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_86),
.Y(n_123)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_61),
.B(n_32),
.Y(n_87)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_41),
.B(n_21),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_91),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_43),
.B(n_29),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_42),
.B(n_30),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_99),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_48),
.A2(n_16),
.B1(n_18),
.B2(n_35),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_96),
.A2(n_19),
.B1(n_25),
.B2(n_33),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_50),
.B(n_19),
.Y(n_98)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_30),
.Y(n_99)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_29),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_103),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_45),
.B(n_29),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_42),
.A2(n_25),
.B1(n_37),
.B2(n_33),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_64),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_111),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_79),
.A2(n_23),
.B(n_22),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_108),
.A2(n_126),
.B(n_15),
.Y(n_162)
);

AND2x6_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_80),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_110),
.A2(n_125),
.B1(n_15),
.B2(n_100),
.Y(n_160)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_64),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_114),
.B(n_116),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_74),
.A2(n_25),
.B1(n_23),
.B2(n_19),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_67),
.B1(n_105),
.B2(n_92),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_117),
.B(n_120),
.Y(n_166)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_65),
.B1(n_86),
.B2(n_101),
.Y(n_151)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_71),
.B(n_2),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_33),
.B1(n_6),
.B2(n_7),
.Y(n_126)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_132),
.A2(n_69),
.B1(n_74),
.B2(n_78),
.Y(n_142)
);

INVx4_ASAP7_75t_SL g134 ( 
.A(n_92),
.Y(n_134)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_67),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_136),
.B(n_138),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_SL g152 ( 
.A1(n_137),
.A2(n_12),
.B(n_13),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_99),
.B(n_6),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_141),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_10),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_142),
.A2(n_152),
.B1(n_158),
.B2(n_162),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_143),
.B(n_159),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_119),
.B(n_103),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_145),
.B(n_149),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_105),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_148),
.A2(n_156),
.B(n_137),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_118),
.B(n_97),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_70),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_163),
.C(n_164),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_126),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_14),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_110),
.A2(n_65),
.B1(n_73),
.B2(n_72),
.Y(n_157)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

OAI22x1_ASAP7_75t_SL g158 ( 
.A1(n_131),
.A2(n_88),
.B1(n_73),
.B2(n_104),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_118),
.B(n_97),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_168),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_75),
.C(n_83),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_88),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_141),
.B(n_15),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_83),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_171),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_121),
.B(n_90),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_147),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_131),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_130),
.Y(n_172)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_174),
.A2(n_117),
.B1(n_138),
.B2(n_166),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_180),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_128),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_124),
.C(n_109),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_191),
.C(n_196),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_165),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_184),
.B(n_187),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_189),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_131),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

NOR3xp33_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_108),
.C(n_125),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_133),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_153),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_192),
.B(n_197),
.Y(n_211)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_195),
.A2(n_156),
.B(n_116),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_148),
.B(n_122),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_144),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_124),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_155),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_179),
.B(n_145),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_207),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_203),
.B1(n_212),
.B2(n_187),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_167),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_202),
.A2(n_210),
.B1(n_217),
.B2(n_174),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_160),
.B1(n_162),
.B2(n_154),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_157),
.C(n_154),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_208),
.C(n_215),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_178),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_180),
.C(n_176),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_199),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_SL g210 ( 
.A1(n_178),
.A2(n_142),
.B(n_143),
.C(n_129),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_175),
.A2(n_163),
.B1(n_156),
.B2(n_155),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_213),
.B(n_195),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_123),
.C(n_127),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_174),
.A2(n_144),
.B1(n_134),
.B2(n_146),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_216),
.Y(n_218)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_218),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_219),
.A2(n_220),
.B1(n_225),
.B2(n_226),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_224),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_198),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_222),
.A2(n_229),
.B(n_202),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_191),
.C(n_182),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_207),
.A2(n_173),
.B1(n_190),
.B2(n_196),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_211),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_228),
.A2(n_230),
.B1(n_214),
.B2(n_212),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_194),
.C(n_179),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_184),
.Y(n_231)
);

BUFx24_ASAP7_75t_SL g233 ( 
.A(n_231),
.Y(n_233)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_231),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_227),
.A2(n_210),
.B(n_205),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_238),
.A2(n_240),
.B(n_221),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_220),
.A2(n_210),
.B1(n_215),
.B2(n_204),
.Y(n_239)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_224),
.A2(n_210),
.B(n_183),
.Y(n_240)
);

AOI31xp67_ASAP7_75t_L g242 ( 
.A1(n_238),
.A2(n_240),
.A3(n_235),
.B(n_237),
.Y(n_242)
);

NAND2xp33_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_186),
.Y(n_254)
);

A2O1A1Ixp33_ASAP7_75t_SL g250 ( 
.A1(n_243),
.A2(n_248),
.B(n_233),
.C(n_111),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_236),
.B(n_185),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_246),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_247),
.C(n_243),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_R g246 ( 
.A1(n_234),
.A2(n_229),
.B1(n_225),
.B2(n_223),
.Y(n_246)
);

AOI21x1_ASAP7_75t_SL g248 ( 
.A1(n_234),
.A2(n_222),
.B(n_223),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_249),
.B(n_252),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_250),
.A2(n_248),
.B(n_185),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_183),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_242),
.B(n_188),
.Y(n_253)
);

OAI21x1_ASAP7_75t_L g258 ( 
.A1(n_253),
.A2(n_254),
.B(n_112),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_256),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_251),
.A2(n_120),
.B1(n_186),
.B2(n_139),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_258),
.A2(n_250),
.B(n_127),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_257),
.Y(n_261)
);

FAx1_ASAP7_75t_SL g262 ( 
.A(n_261),
.B(n_259),
.CI(n_139),
.CON(n_262),
.SN(n_262)
);


endmodule