module fake_aes_5543_n_449 (n_117, n_44, n_133, n_149, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_107, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_125, n_9, n_10, n_130, n_103, n_19, n_87, n_137, n_104, n_98, n_74, n_154, n_7, n_29, n_146, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_152, n_113, n_95, n_124, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_40, n_111, n_79, n_38, n_64, n_142, n_46, n_31, n_58, n_122, n_138, n_126, n_118, n_32, n_0, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_75, n_105, n_72, n_136, n_43, n_76, n_89, n_68, n_144, n_27, n_53, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_3, n_18, n_110, n_66, n_134, n_1, n_82, n_106, n_15, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_449);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_107;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_125;
input n_9;
input n_10;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_104;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_146;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_152;
input n_113;
input n_95;
input n_124;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_142;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_118;
input n_32;
input n_0;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_75;
input n_105;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_68;
input n_144;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_82;
input n_106;
input n_15;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_449;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_431;
wire n_161;
wire n_177;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_328;
wire n_229;
wire n_336;
wire n_448;
wire n_348;
wire n_252;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_232;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_384;
wire n_227;
wire n_231;
wire n_298;
wire n_411;
wire n_183;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_443;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_277;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_238;
wire n_318;
wire n_293;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_299;
wire n_338;
wire n_256;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_362;
wire n_259;
wire n_308;
wire n_412;
wire n_207;
wire n_224;
wire n_219;
wire n_214;
wire n_204;
wire n_430;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_379;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_388;
wire n_193;
wire n_273;
wire n_390;
wire n_245;
wire n_357;
wire n_260;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_178;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_283;
wire n_435;
wire n_216;
wire n_212;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_429;
wire n_233;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_203;
wire n_300;
wire n_158;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_335;
wire n_272;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_343;
wire n_291;
wire n_170;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_187;
wire n_375;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_223;
wire n_372;
wire n_194;
wire n_287;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_406;
wire n_395;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g156 ( .A(n_8), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_55), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_46), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_144), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_2), .Y(n_160) );
BUFx3_ASAP7_75t_L g161 ( .A(n_127), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_38), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_59), .Y(n_163) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_37), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_28), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_1), .Y(n_166) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_136), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_142), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_41), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_77), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_154), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_82), .Y(n_172) );
CKINVDCx16_ASAP7_75t_R g173 ( .A(n_109), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_112), .Y(n_174) );
INVxp67_ASAP7_75t_L g175 ( .A(n_151), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_50), .Y(n_176) );
INVx2_ASAP7_75t_SL g177 ( .A(n_141), .Y(n_177) );
NOR2xp67_ASAP7_75t_L g178 ( .A(n_130), .B(n_22), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_145), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_23), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_15), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_134), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_143), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_123), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_147), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_104), .Y(n_186) );
NOR2xp67_ASAP7_75t_L g187 ( .A(n_139), .B(n_80), .Y(n_187) );
INVx2_ASAP7_75t_SL g188 ( .A(n_129), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_66), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_94), .Y(n_190) );
BUFx10_ASAP7_75t_L g191 ( .A(n_97), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_69), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_118), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_132), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_101), .B(n_6), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_146), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_135), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_84), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_99), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_137), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_152), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_83), .Y(n_202) );
INVx2_ASAP7_75t_SL g203 ( .A(n_149), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_138), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_119), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_140), .B(n_87), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_74), .Y(n_207) );
INVxp67_ASAP7_75t_L g208 ( .A(n_133), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_45), .Y(n_209) );
INVxp67_ASAP7_75t_SL g210 ( .A(n_48), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_64), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_72), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_25), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_102), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_131), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_70), .Y(n_216) );
BUFx2_ASAP7_75t_L g217 ( .A(n_150), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_16), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_35), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_32), .Y(n_220) );
CKINVDCx14_ASAP7_75t_R g221 ( .A(n_63), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_116), .Y(n_222) );
NOR2xp67_ASAP7_75t_L g223 ( .A(n_92), .B(n_44), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_42), .Y(n_224) );
CKINVDCx16_ASAP7_75t_R g225 ( .A(n_24), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_128), .Y(n_226) );
INVxp67_ASAP7_75t_SL g227 ( .A(n_58), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_62), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_148), .Y(n_229) );
NOR2xp67_ASAP7_75t_L g230 ( .A(n_65), .B(n_68), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_86), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_73), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_113), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_21), .Y(n_234) );
INVxp67_ASAP7_75t_L g235 ( .A(n_53), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_81), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_47), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_43), .Y(n_238) );
INVx1_ASAP7_75t_SL g239 ( .A(n_71), .Y(n_239) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_157), .A2(n_11), .B(n_10), .Y(n_240) );
AND2x4_ASAP7_75t_L g241 ( .A(n_217), .B(n_0), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_219), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_166), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_177), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_188), .B(n_0), .Y(n_245) );
INVx3_ASAP7_75t_L g246 ( .A(n_191), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_203), .Y(n_247) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_156), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_164), .B(n_1), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_167), .B(n_2), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_163), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_168), .Y(n_252) );
INVx5_ASAP7_75t_L g253 ( .A(n_219), .Y(n_253) );
OAI21x1_ASAP7_75t_L g254 ( .A1(n_176), .A2(n_13), .B(n_12), .Y(n_254) );
INVx3_ASAP7_75t_L g255 ( .A(n_182), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_219), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_253), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_244), .Y(n_258) );
INVxp33_ASAP7_75t_L g259 ( .A(n_243), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_246), .B(n_173), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_247), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_255), .Y(n_262) );
INVx3_ASAP7_75t_L g263 ( .A(n_255), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_245), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_245), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_251), .B(n_225), .Y(n_266) );
AND2x6_ASAP7_75t_L g267 ( .A(n_241), .B(n_169), .Y(n_267) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_242), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_264), .A2(n_248), .B1(n_252), .B2(n_205), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_265), .A2(n_241), .B1(n_252), .B2(n_250), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_258), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_266), .B(n_249), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_257), .Y(n_273) );
O2A1O1Ixp5_ASAP7_75t_L g274 ( .A1(n_260), .A2(n_195), .B(n_227), .C(n_210), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_259), .B(n_158), .Y(n_275) );
A2O1A1Ixp33_ASAP7_75t_L g276 ( .A1(n_261), .A2(n_254), .B(n_208), .C(n_228), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_267), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_263), .B(n_159), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_267), .B(n_221), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_263), .B(n_162), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_262), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_267), .B(n_175), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g283 ( .A1(n_267), .A2(n_171), .B1(n_172), .B2(n_170), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_269), .B(n_160), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_269), .A2(n_229), .B1(n_237), .B2(n_215), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_272), .B(n_175), .Y(n_286) );
INVx3_ASAP7_75t_L g287 ( .A(n_277), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_275), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_270), .B(n_235), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_276), .A2(n_240), .B(n_206), .Y(n_290) );
O2A1O1Ixp33_ASAP7_75t_L g291 ( .A1(n_282), .A2(n_174), .B(n_181), .C(n_179), .Y(n_291) );
OAI21xp5_ASAP7_75t_L g292 ( .A1(n_274), .A2(n_240), .B(n_190), .Y(n_292) );
NOR2xp67_ASAP7_75t_L g293 ( .A(n_277), .B(n_14), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_271), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_281), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_282), .A2(n_193), .B(n_184), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_283), .B(n_165), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_273), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_279), .A2(n_198), .B(n_196), .Y(n_299) );
OA22x2_ASAP7_75t_L g300 ( .A1(n_278), .A2(n_200), .B1(n_201), .B2(n_199), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_290), .A2(n_280), .B(n_277), .Y(n_301) );
OAI21x1_ASAP7_75t_L g302 ( .A1(n_292), .A2(n_214), .B(n_211), .Y(n_302) );
NAND2x1p5_ASAP7_75t_L g303 ( .A(n_285), .B(n_239), .Y(n_303) );
INVxp67_ASAP7_75t_SL g304 ( .A(n_284), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_289), .B(n_3), .Y(n_305) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_287), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_296), .A2(n_220), .B(n_218), .Y(n_307) );
AO32x2_ASAP7_75t_L g308 ( .A1(n_300), .A2(n_242), .A3(n_256), .B1(n_187), .B2(n_178), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_295), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_298), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_288), .B(n_180), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_291), .B(n_299), .Y(n_312) );
AO32x2_ASAP7_75t_L g313 ( .A1(n_293), .A2(n_242), .A3(n_256), .B1(n_230), .B2(n_223), .Y(n_313) );
A2O1A1Ixp33_ASAP7_75t_L g314 ( .A1(n_297), .A2(n_232), .B(n_233), .C(n_231), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_294), .Y(n_315) );
OAI21x1_ASAP7_75t_L g316 ( .A1(n_290), .A2(n_236), .B(n_234), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_286), .B(n_238), .Y(n_317) );
OAI21x1_ASAP7_75t_L g318 ( .A1(n_316), .A2(n_226), .B(n_224), .Y(n_318) );
OA21x2_ASAP7_75t_L g319 ( .A1(n_302), .A2(n_185), .B(n_183), .Y(n_319) );
OAI21x1_ASAP7_75t_SL g320 ( .A1(n_301), .A2(n_3), .B(n_4), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_304), .B(n_4), .Y(n_321) );
OR2x6_ASAP7_75t_L g322 ( .A(n_303), .B(n_161), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_309), .Y(n_323) );
NOR2xp33_ASAP7_75t_R g324 ( .A(n_311), .B(n_5), .Y(n_324) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_306), .Y(n_325) );
A2O1A1Ixp33_ASAP7_75t_L g326 ( .A1(n_312), .A2(n_189), .B(n_192), .C(n_186), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_315), .B(n_5), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_310), .Y(n_328) );
AO31x2_ASAP7_75t_L g329 ( .A1(n_314), .A2(n_268), .A3(n_17), .B(n_18), .Y(n_329) );
AO31x2_ASAP7_75t_L g330 ( .A1(n_307), .A2(n_268), .A3(n_19), .B(n_20), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_305), .Y(n_331) );
INVx3_ASAP7_75t_L g332 ( .A(n_306), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_317), .A2(n_268), .B(n_197), .Y(n_333) );
OR2x6_ASAP7_75t_L g334 ( .A(n_308), .B(n_7), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_313), .Y(n_335) );
OAI21x1_ASAP7_75t_SL g336 ( .A1(n_312), .A2(n_8), .B(n_9), .Y(n_336) );
A2O1A1Ixp33_ASAP7_75t_L g337 ( .A1(n_312), .A2(n_202), .B(n_204), .C(n_194), .Y(n_337) );
AO21x2_ASAP7_75t_L g338 ( .A1(n_302), .A2(n_27), .B(n_26), .Y(n_338) );
OAI21x1_ASAP7_75t_L g339 ( .A1(n_316), .A2(n_30), .B(n_29), .Y(n_339) );
OAI21x1_ASAP7_75t_L g340 ( .A1(n_316), .A2(n_33), .B(n_31), .Y(n_340) );
OAI21xp5_ASAP7_75t_L g341 ( .A1(n_321), .A2(n_209), .B(n_207), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_328), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_320), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_320), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_324), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_336), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_332), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_327), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_334), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_334), .Y(n_350) );
OAI21x1_ASAP7_75t_L g351 ( .A1(n_318), .A2(n_36), .B(n_34), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_339), .Y(n_352) );
INVx3_ASAP7_75t_L g353 ( .A(n_340), .Y(n_353) );
INVx2_ASAP7_75t_SL g354 ( .A(n_329), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_330), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_338), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_319), .Y(n_357) );
INVxp67_ASAP7_75t_R g358 ( .A(n_326), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_333), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_337), .Y(n_360) );
OA21x2_ASAP7_75t_L g361 ( .A1(n_335), .A2(n_213), .B(n_212), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_331), .B(n_216), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_323), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_323), .Y(n_364) );
NAND2x1p5_ASAP7_75t_L g365 ( .A(n_325), .B(n_39), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_323), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_323), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_323), .B(n_40), .Y(n_368) );
INVx4_ASAP7_75t_SL g369 ( .A(n_322), .Y(n_369) );
AND2x4_ASAP7_75t_SL g370 ( .A(n_322), .B(n_222), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_323), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_366), .B(n_367), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_342), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_369), .B(n_49), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_363), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_364), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_370), .A2(n_51), .B1(n_52), .B2(n_54), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_364), .B(n_56), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_349), .A2(n_57), .B1(n_60), .B2(n_61), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_345), .B(n_155), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_371), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_350), .B(n_67), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_368), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_344), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_343), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_355), .Y(n_386) );
INVxp67_ASAP7_75t_SL g387 ( .A(n_357), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_352), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_348), .A2(n_75), .B1(n_76), .B2(n_78), .C(n_79), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_346), .B(n_359), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_347), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g392 ( .A1(n_358), .A2(n_360), .B1(n_362), .B2(n_341), .Y(n_392) );
BUFx3_ASAP7_75t_L g393 ( .A(n_365), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_356), .B(n_153), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_351), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_353), .Y(n_396) );
INVx3_ASAP7_75t_L g397 ( .A(n_361), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_354), .B(n_85), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_376), .B(n_88), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_375), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_373), .B(n_89), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_372), .B(n_90), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_381), .Y(n_403) );
AND2x4_ASAP7_75t_SL g404 ( .A(n_383), .B(n_91), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_384), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_386), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_391), .B(n_93), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_388), .B(n_95), .Y(n_408) );
AND2x4_ASAP7_75t_SL g409 ( .A(n_374), .B(n_96), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_382), .B(n_98), .Y(n_410) );
INVx3_ASAP7_75t_L g411 ( .A(n_393), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_390), .B(n_100), .Y(n_412) );
INVxp67_ASAP7_75t_L g413 ( .A(n_397), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_387), .Y(n_414) );
INVx3_ASAP7_75t_L g415 ( .A(n_398), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_385), .Y(n_416) );
AND2x4_ASAP7_75t_L g417 ( .A(n_385), .B(n_103), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_378), .B(n_105), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_396), .B(n_106), .Y(n_419) );
AND3x1_ASAP7_75t_L g420 ( .A(n_411), .B(n_380), .C(n_392), .Y(n_420) );
AND2x2_ASAP7_75t_SL g421 ( .A(n_409), .B(n_394), .Y(n_421) );
NOR2xp67_ASAP7_75t_L g422 ( .A(n_414), .B(n_413), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_400), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_403), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_406), .B(n_405), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_416), .Y(n_426) );
BUFx2_ASAP7_75t_L g427 ( .A(n_419), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_425), .Y(n_428) );
AND2x2_ASAP7_75t_SL g429 ( .A(n_421), .B(n_409), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_426), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_423), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_424), .B(n_415), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_428), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_429), .A2(n_420), .B1(n_422), .B2(n_427), .Y(n_434) );
OAI31xp33_ASAP7_75t_L g435 ( .A1(n_434), .A2(n_432), .A3(n_430), .B(n_431), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_433), .Y(n_436) );
NAND4xp25_ASAP7_75t_L g437 ( .A(n_435), .B(n_377), .C(n_379), .D(n_402), .Y(n_437) );
NAND3xp33_ASAP7_75t_L g438 ( .A(n_436), .B(n_389), .C(n_412), .Y(n_438) );
NOR2xp33_ASAP7_75t_SL g439 ( .A(n_437), .B(n_410), .Y(n_439) );
AOI211xp5_ASAP7_75t_L g440 ( .A1(n_439), .A2(n_438), .B(n_418), .C(n_407), .Y(n_440) );
OAI221xp5_ASAP7_75t_SL g441 ( .A1(n_440), .A2(n_408), .B1(n_399), .B2(n_401), .C(n_395), .Y(n_441) );
NOR3xp33_ASAP7_75t_L g442 ( .A(n_441), .B(n_417), .C(n_419), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_442), .B(n_404), .Y(n_443) );
INVx2_ASAP7_75t_SL g444 ( .A(n_443), .Y(n_444) );
AOI31xp33_ASAP7_75t_L g445 ( .A1(n_444), .A2(n_107), .A3(n_108), .B(n_110), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_445), .A2(n_111), .B1(n_114), .B2(n_115), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_446), .B(n_117), .Y(n_447) );
AOI221xp5_ASAP7_75t_L g448 ( .A1(n_447), .A2(n_120), .B1(n_121), .B2(n_122), .C(n_124), .Y(n_448) );
AO21x2_ASAP7_75t_L g449 ( .A1(n_448), .A2(n_125), .B(n_126), .Y(n_449) );
endmodule