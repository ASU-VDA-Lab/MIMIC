module fake_jpeg_2972_n_126 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_126);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_39),
.Y(n_50)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_54),
.Y(n_64)
);

INVx2_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_0),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_47),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_65),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_50),
.A2(n_47),
.B1(n_39),
.B2(n_37),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_49),
.B1(n_55),
.B2(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_61),
.B(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_52),
.B(n_42),
.C(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_67),
.B(n_73),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_20),
.Y(n_91)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_59),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

AOI221xp5_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_75),
.B1(n_36),
.B2(n_46),
.C(n_44),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_36),
.Y(n_73)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_49),
.B1(n_41),
.B2(n_38),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_41),
.Y(n_80)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_80),
.B(n_6),
.Y(n_102)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_22),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_38),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_67),
.C(n_70),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_86),
.A2(n_74),
.B1(n_76),
.B2(n_72),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_1),
.B(n_2),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_5),
.B(n_6),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_3),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_90),
.B(n_23),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_84),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_98),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_95),
.B(n_96),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_82),
.B(n_5),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_100),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_72),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

OA21x2_ASAP7_75t_SL g111 ( 
.A1(n_101),
.A2(n_102),
.B(n_103),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_7),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_7),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_104),
.A2(n_105),
.B(n_106),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_8),
.Y(n_105)
);

OAI321xp33_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_92),
.A3(n_89),
.B1(n_27),
.B2(n_28),
.C(n_34),
.Y(n_107)
);

OAI322xp33_ASAP7_75t_L g116 ( 
.A1(n_107),
.A2(n_9),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_15),
.C2(n_17),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_95),
.A2(n_83),
.B1(n_81),
.B2(n_11),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_109),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_81),
.B(n_10),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_115),
.A2(n_9),
.B(n_12),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_118),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_97),
.C(n_25),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_110),
.C(n_111),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_114),
.B(n_113),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_108),
.C(n_121),
.Y(n_123)
);

AOI322xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_115),
.A3(n_119),
.B1(n_109),
.B2(n_30),
.C1(n_31),
.C2(n_33),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_21),
.C(n_24),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_13),
.Y(n_126)
);


endmodule