module fake_aes_6617_n_1232 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_280, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1232);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1232;
wire n_963;
wire n_1034;
wire n_949;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_677;
wire n_756;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_994;
wire n_930;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_795;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_713;
wire n_457;
wire n_736;
wire n_287;
wire n_606;
wire n_332;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_791;
wire n_707;
wire n_603;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_336;
wire n_464;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_366;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_313;
wire n_322;
wire n_427;
wire n_703;
wire n_415;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_416;
wire n_536;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_998;
wire n_604;
wire n_755;
wire n_848;
wire n_1031;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1195;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1114;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_924;
wire n_378;
wire n_441;
wire n_335;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_491;
INVx2_ASAP7_75t_L g287 ( .A(n_238), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_143), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_203), .Y(n_289) );
INVxp67_ASAP7_75t_SL g290 ( .A(n_23), .Y(n_290) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_99), .Y(n_291) );
BUFx3_ASAP7_75t_L g292 ( .A(n_92), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_74), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_205), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g295 ( .A(n_104), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_122), .Y(n_296) );
INVxp67_ASAP7_75t_SL g297 ( .A(n_232), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_116), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_33), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_211), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_7), .Y(n_301) );
CKINVDCx16_ASAP7_75t_R g302 ( .A(n_189), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_140), .Y(n_303) );
BUFx8_ASAP7_75t_SL g304 ( .A(n_163), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_36), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_37), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_68), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_286), .Y(n_308) );
CKINVDCx20_ASAP7_75t_R g309 ( .A(n_23), .Y(n_309) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_110), .Y(n_310) );
CKINVDCx14_ASAP7_75t_R g311 ( .A(n_282), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_72), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_270), .Y(n_313) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_47), .Y(n_314) );
CKINVDCx16_ASAP7_75t_R g315 ( .A(n_222), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_172), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_38), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_62), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_137), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_219), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_208), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_192), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_262), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_141), .Y(n_324) );
INVxp67_ASAP7_75t_SL g325 ( .A(n_114), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_239), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_186), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_8), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_252), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_250), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_247), .Y(n_331) );
BUFx3_ASAP7_75t_L g332 ( .A(n_214), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_277), .Y(n_333) );
INVxp67_ASAP7_75t_SL g334 ( .A(n_98), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_76), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_127), .Y(n_336) );
INVxp67_ASAP7_75t_SL g337 ( .A(n_161), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_10), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_221), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_198), .Y(n_340) );
CKINVDCx20_ASAP7_75t_R g341 ( .A(n_202), .Y(n_341) );
INVx1_ASAP7_75t_SL g342 ( .A(n_265), .Y(n_342) );
BUFx5_ASAP7_75t_L g343 ( .A(n_66), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_190), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_111), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_78), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_183), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_5), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_72), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_169), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_228), .Y(n_351) );
CKINVDCx16_ASAP7_75t_R g352 ( .A(n_134), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_242), .Y(n_353) );
BUFx8_ASAP7_75t_SL g354 ( .A(n_27), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_28), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_158), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_117), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_244), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_142), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_260), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_188), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_181), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_124), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_179), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_206), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_121), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_126), .Y(n_367) );
BUFx3_ASAP7_75t_L g368 ( .A(n_261), .Y(n_368) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_108), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_253), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_14), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_2), .Y(n_372) );
CKINVDCx20_ASAP7_75t_R g373 ( .A(n_174), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_240), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_16), .B(n_3), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_182), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_82), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_113), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_275), .Y(n_379) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_37), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_112), .Y(n_381) );
CKINVDCx20_ASAP7_75t_R g382 ( .A(n_153), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_272), .Y(n_383) );
BUFx5_ASAP7_75t_L g384 ( .A(n_185), .Y(n_384) );
INVxp67_ASAP7_75t_SL g385 ( .A(n_109), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_194), .Y(n_386) );
BUFx5_ASAP7_75t_L g387 ( .A(n_271), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_45), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_168), .Y(n_389) );
CKINVDCx20_ASAP7_75t_R g390 ( .A(n_35), .Y(n_390) );
INVx1_ASAP7_75t_SL g391 ( .A(n_115), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_52), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_218), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_268), .Y(n_394) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_278), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_80), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_167), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_87), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_57), .Y(n_399) );
INVxp67_ASAP7_75t_L g400 ( .A(n_274), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_148), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_187), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_258), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_233), .Y(n_404) );
BUFx3_ASAP7_75t_L g405 ( .A(n_84), .Y(n_405) );
NOR2xp67_ASAP7_75t_L g406 ( .A(n_209), .B(n_234), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_284), .Y(n_407) );
CKINVDCx20_ASAP7_75t_R g408 ( .A(n_269), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_14), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_159), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_173), .Y(n_411) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_285), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_6), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_56), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_254), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_207), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_246), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_251), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_229), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_164), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_58), .Y(n_421) );
INVx1_ASAP7_75t_SL g422 ( .A(n_171), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_36), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_256), .Y(n_424) );
INVxp67_ASAP7_75t_SL g425 ( .A(n_102), .Y(n_425) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_118), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_170), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_26), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_11), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_105), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_15), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_160), .Y(n_432) );
NOR2xp67_ASAP7_75t_L g433 ( .A(n_49), .B(n_93), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g434 ( .A(n_210), .Y(n_434) );
BUFx3_ASAP7_75t_L g435 ( .A(n_24), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_73), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_24), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_226), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_263), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_86), .Y(n_440) );
BUFx2_ASAP7_75t_L g441 ( .A(n_225), .Y(n_441) );
BUFx2_ASAP7_75t_L g442 ( .A(n_40), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_237), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_107), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_74), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_38), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_62), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_162), .Y(n_448) );
INVxp67_ASAP7_75t_L g449 ( .A(n_77), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_11), .Y(n_450) );
AND2x4_ASAP7_75t_L g451 ( .A(n_324), .B(n_0), .Y(n_451) );
BUFx3_ASAP7_75t_L g452 ( .A(n_289), .Y(n_452) );
OAI22xp5_ASAP7_75t_SL g453 ( .A1(n_390), .A2(n_2), .B1(n_0), .B2(n_1), .Y(n_453) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_291), .Y(n_454) );
AND2x4_ASAP7_75t_L g455 ( .A(n_324), .B(n_1), .Y(n_455) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_291), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_384), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_395), .B(n_3), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_384), .Y(n_459) );
OA21x2_ASAP7_75t_L g460 ( .A1(n_287), .A2(n_85), .B(n_83), .Y(n_460) );
BUFx3_ASAP7_75t_L g461 ( .A(n_289), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_395), .B(n_4), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_314), .A2(n_6), .B1(n_4), .B2(n_5), .Y(n_463) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_291), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_384), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_314), .B(n_8), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_435), .B(n_9), .Y(n_467) );
BUFx3_ASAP7_75t_L g468 ( .A(n_292), .Y(n_468) );
BUFx2_ASAP7_75t_L g469 ( .A(n_442), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_441), .B(n_9), .Y(n_470) );
BUFx3_ASAP7_75t_L g471 ( .A(n_292), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_435), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_384), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_311), .B(n_10), .Y(n_474) );
INVx4_ASAP7_75t_L g475 ( .A(n_332), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_311), .B(n_12), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_354), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_354), .Y(n_478) );
NOR2xp33_ASAP7_75t_SL g479 ( .A(n_302), .B(n_283), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_343), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_343), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_449), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_384), .Y(n_483) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_291), .Y(n_484) );
OAI21x1_ASAP7_75t_L g485 ( .A1(n_287), .A2(n_89), .B(n_88), .Y(n_485) );
BUFx8_ASAP7_75t_L g486 ( .A(n_384), .Y(n_486) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_299), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_387), .B(n_13), .Y(n_488) );
AOI22xp5_ASAP7_75t_SL g489 ( .A1(n_390), .A2(n_17), .B1(n_15), .B2(n_16), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_472), .B(n_315), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_457), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_457), .Y(n_492) );
NOR2x1p5_ASAP7_75t_L g493 ( .A(n_458), .B(n_290), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_457), .Y(n_494) );
BUFx3_ASAP7_75t_L g495 ( .A(n_452), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_459), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_459), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_459), .Y(n_498) );
INVxp33_ASAP7_75t_SL g499 ( .A(n_477), .Y(n_499) );
BUFx4f_ASAP7_75t_L g500 ( .A(n_467), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_486), .B(n_352), .Y(n_501) );
INVx5_ASAP7_75t_L g502 ( .A(n_475), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_465), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_465), .Y(n_504) );
INVx2_ASAP7_75t_SL g505 ( .A(n_486), .Y(n_505) );
OAI22x1_ASAP7_75t_L g506 ( .A1(n_463), .A2(n_305), .B1(n_306), .B2(n_301), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_465), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_473), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_472), .B(n_343), .Y(n_509) );
INVx3_ASAP7_75t_L g510 ( .A(n_467), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_473), .Y(n_511) );
BUFx4f_ASAP7_75t_L g512 ( .A(n_467), .Y(n_512) );
INVx2_ASAP7_75t_SL g513 ( .A(n_486), .Y(n_513) );
INVx2_ASAP7_75t_SL g514 ( .A(n_486), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_473), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_475), .B(n_312), .Y(n_516) );
BUFx10_ASAP7_75t_L g517 ( .A(n_451), .Y(n_517) );
NOR2x1p5_ASAP7_75t_L g518 ( .A(n_458), .B(n_317), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_483), .Y(n_519) );
INVx3_ASAP7_75t_L g520 ( .A(n_467), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_483), .Y(n_521) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_454), .Y(n_522) );
AND2x4_ASAP7_75t_L g523 ( .A(n_451), .B(n_450), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_487), .B(n_400), .Y(n_524) );
BUFx10_ASAP7_75t_L g525 ( .A(n_451), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_483), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_480), .Y(n_527) );
INVx2_ASAP7_75t_SL g528 ( .A(n_474), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_480), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_469), .B(n_343), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_481), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_481), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_454), .Y(n_533) );
INVx2_ASAP7_75t_SL g534 ( .A(n_474), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_485), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_475), .B(n_318), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_485), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_485), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_452), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_509), .Y(n_540) );
INVx4_ASAP7_75t_L g541 ( .A(n_517), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_509), .Y(n_542) );
INVx2_ASAP7_75t_SL g543 ( .A(n_493), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_490), .B(n_451), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_495), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_500), .A2(n_455), .B1(n_466), .B2(n_476), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_530), .B(n_455), .Y(n_547) );
INVxp67_ASAP7_75t_SL g548 ( .A(n_500), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_530), .B(n_455), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_524), .B(n_487), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_528), .B(n_534), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_500), .A2(n_460), .B(n_488), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_528), .B(n_455), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_539), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_512), .A2(n_466), .B1(n_476), .B2(n_462), .Y(n_555) );
INVx5_ASAP7_75t_L g556 ( .A(n_502), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_534), .B(n_523), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_523), .B(n_469), .Y(n_558) );
INVx2_ASAP7_75t_SL g559 ( .A(n_493), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_512), .A2(n_408), .B1(n_295), .B2(n_463), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_523), .B(n_482), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_523), .B(n_482), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_517), .Y(n_563) );
AOI221xp5_ASAP7_75t_L g564 ( .A1(n_506), .A2(n_462), .B1(n_478), .B2(n_477), .C(n_470), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_516), .B(n_470), .Y(n_565) );
OAI21xp5_ASAP7_75t_L g566 ( .A1(n_535), .A2(n_538), .B(n_537), .Y(n_566) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_505), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_525), .Y(n_568) );
BUFx3_ASAP7_75t_L g569 ( .A(n_499), .Y(n_569) );
INVx3_ASAP7_75t_L g570 ( .A(n_525), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_505), .B(n_479), .Y(n_571) );
OR2x6_ASAP7_75t_L g572 ( .A(n_506), .B(n_478), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_536), .B(n_452), .Y(n_573) );
XOR2xp5_ASAP7_75t_L g574 ( .A(n_501), .B(n_489), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_510), .B(n_475), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_525), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_518), .B(n_461), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_510), .A2(n_468), .B1(n_471), .B2(n_461), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_518), .B(n_468), .Y(n_579) );
INVx3_ASAP7_75t_L g580 ( .A(n_510), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_513), .B(n_468), .Y(n_581) );
INVxp67_ASAP7_75t_L g582 ( .A(n_513), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_520), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_520), .B(n_489), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_520), .B(n_471), .Y(n_585) );
NOR2x2_ASAP7_75t_L g586 ( .A(n_494), .B(n_453), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_491), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_514), .B(n_471), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_529), .B(n_300), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_514), .B(n_288), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_529), .B(n_294), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_531), .B(n_303), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_502), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_531), .A2(n_295), .B1(n_408), .B2(n_453), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_535), .A2(n_341), .B1(n_373), .B2(n_310), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_492), .B(n_298), .Y(n_596) );
NAND2x1p5_ASAP7_75t_L g597 ( .A(n_502), .B(n_375), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g598 ( .A(n_492), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_496), .Y(n_599) );
NAND2x1p5_ASAP7_75t_L g600 ( .A(n_502), .B(n_293), .Y(n_600) );
OAI22xp5_ASAP7_75t_SL g601 ( .A1(n_537), .A2(n_309), .B1(n_412), .B2(n_382), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_497), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_527), .B(n_313), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_502), .B(n_308), .Y(n_604) );
INVx4_ASAP7_75t_L g605 ( .A(n_527), .Y(n_605) );
NOR3xp33_ASAP7_75t_L g606 ( .A(n_498), .B(n_414), .C(n_409), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_532), .B(n_319), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_532), .B(n_320), .Y(n_608) );
INVx3_ASAP7_75t_L g609 ( .A(n_511), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_498), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_511), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_519), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g613 ( .A1(n_538), .A2(n_460), .B(n_322), .Y(n_613) );
INVx3_ASAP7_75t_L g614 ( .A(n_519), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_503), .A2(n_460), .B(n_322), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_504), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_507), .B(n_323), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_507), .B(n_423), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_508), .B(n_436), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_508), .B(n_437), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_515), .A2(n_439), .B1(n_426), .B2(n_328), .Y(n_621) );
NAND2x1p5_ASAP7_75t_L g622 ( .A(n_515), .B(n_307), .Y(n_622) );
OR2x6_ASAP7_75t_L g623 ( .A(n_521), .B(n_335), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_521), .B(n_321), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_526), .A2(n_346), .B1(n_348), .B2(n_338), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_526), .B(n_330), .Y(n_626) );
OR2x6_ASAP7_75t_L g627 ( .A(n_601), .B(n_349), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_546), .A2(n_371), .B1(n_372), .B2(n_355), .Y(n_628) );
BUFx2_ASAP7_75t_L g629 ( .A(n_569), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_541), .B(n_326), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g631 ( .A1(n_566), .A2(n_460), .B(n_325), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_560), .B(n_377), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_605), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_565), .B(n_388), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_550), .B(n_304), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_552), .A2(n_460), .B(n_334), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_555), .B(n_392), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_567), .B(n_327), .Y(n_638) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_623), .Y(n_639) );
NOR2x1_ASAP7_75t_L g640 ( .A(n_558), .B(n_396), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_613), .A2(n_337), .B(n_297), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_567), .B(n_331), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_573), .A2(n_425), .B(n_385), .Y(n_643) );
NOR2xp33_ASAP7_75t_R g644 ( .A(n_593), .B(n_333), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_582), .B(n_336), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_582), .B(n_350), .Y(n_646) );
OAI21xp5_ASAP7_75t_L g647 ( .A1(n_615), .A2(n_340), .B(n_339), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_544), .A2(n_345), .B(n_344), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_584), .A2(n_413), .B1(n_421), .B2(n_399), .Y(n_649) );
AND2x2_ASAP7_75t_SL g650 ( .A(n_594), .B(n_304), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_550), .B(n_428), .Y(n_651) );
AND2x4_ASAP7_75t_L g652 ( .A(n_623), .B(n_429), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_585), .A2(n_351), .B(n_347), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_555), .B(n_431), .Y(n_654) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_556), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_551), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_557), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_546), .A2(n_445), .B1(n_447), .B2(n_446), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_580), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_598), .A2(n_380), .B1(n_356), .B2(n_357), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g661 ( .A1(n_571), .A2(n_358), .B(n_353), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_571), .A2(n_360), .B(n_359), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_588), .A2(n_362), .B(n_361), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_561), .B(n_316), .Y(n_664) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_623), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_606), .A2(n_363), .B1(n_367), .B2(n_366), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_562), .B(n_342), .Y(n_667) );
BUFx12f_ASAP7_75t_L g668 ( .A(n_572), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_581), .A2(n_381), .B(n_379), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_581), .A2(n_389), .B(n_386), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_575), .A2(n_394), .B(n_393), .Y(n_671) );
O2A1O1Ixp33_ASAP7_75t_L g672 ( .A1(n_547), .A2(n_398), .B(n_401), .C(n_397), .Y(n_672) );
O2A1O1Ixp33_ASAP7_75t_L g673 ( .A1(n_549), .A2(n_410), .B(n_415), .C(n_403), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_543), .B(n_391), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_548), .A2(n_380), .B1(n_417), .B2(n_416), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_548), .A2(n_380), .B1(n_424), .B2(n_419), .Y(n_676) );
O2A1O1Ixp33_ASAP7_75t_L g677 ( .A1(n_540), .A2(n_438), .B(n_440), .C(n_430), .Y(n_677) );
O2A1O1Ixp33_ASAP7_75t_L g678 ( .A1(n_542), .A2(n_444), .B(n_364), .C(n_365), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_621), .B(n_343), .Y(n_679) );
INVx3_ASAP7_75t_L g680 ( .A(n_570), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_622), .A2(n_433), .B1(n_380), .B2(n_364), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_622), .Y(n_682) );
OR2x2_ASAP7_75t_L g683 ( .A(n_595), .B(n_17), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_597), .A2(n_378), .B1(n_383), .B2(n_376), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_583), .A2(n_370), .B(n_296), .Y(n_685) );
O2A1O1Ixp33_ASAP7_75t_SL g686 ( .A1(n_577), .A2(n_422), .B(n_374), .C(n_370), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_618), .B(n_343), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_606), .A2(n_402), .B1(n_407), .B2(n_404), .Y(n_688) );
O2A1O1Ixp33_ASAP7_75t_L g689 ( .A1(n_553), .A2(n_432), .B(n_427), .C(n_368), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_559), .B(n_411), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_580), .Y(n_691) );
CKINVDCx8_ASAP7_75t_R g692 ( .A(n_572), .Y(n_692) );
NOR2x1_ASAP7_75t_L g693 ( .A(n_572), .B(n_332), .Y(n_693) );
INVx3_ASAP7_75t_L g694 ( .A(n_600), .Y(n_694) );
OR2x6_ASAP7_75t_L g695 ( .A(n_597), .B(n_406), .Y(n_695) );
BUFx2_ASAP7_75t_L g696 ( .A(n_619), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_563), .B(n_418), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_620), .B(n_420), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_609), .Y(n_699) );
BUFx3_ASAP7_75t_L g700 ( .A(n_600), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_568), .A2(n_533), .B(n_405), .Y(n_701) );
CKINVDCx8_ASAP7_75t_R g702 ( .A(n_556), .Y(n_702) );
AOI21xp5_ASAP7_75t_L g703 ( .A1(n_576), .A2(n_591), .B(n_596), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_574), .B(n_18), .Y(n_704) );
BUFx2_ASAP7_75t_L g705 ( .A(n_586), .Y(n_705) );
O2A1O1Ixp33_ASAP7_75t_SL g706 ( .A1(n_579), .A2(n_387), .B(n_90), .C(n_91), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_587), .A2(n_443), .B1(n_448), .B2(n_434), .Y(n_707) );
AO21x2_ASAP7_75t_L g708 ( .A1(n_617), .A2(n_387), .B(n_369), .Y(n_708) );
INVxp67_ASAP7_75t_L g709 ( .A(n_589), .Y(n_709) );
NAND3xp33_ASAP7_75t_L g710 ( .A(n_625), .B(n_369), .C(n_329), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_592), .B(n_387), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_592), .B(n_387), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_599), .B(n_19), .Y(n_713) );
A2O1A1Ixp33_ASAP7_75t_L g714 ( .A1(n_603), .A2(n_369), .B(n_329), .C(n_454), .Y(n_714) );
A2O1A1Ixp33_ASAP7_75t_L g715 ( .A1(n_603), .A2(n_329), .B(n_456), .C(n_454), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_602), .A2(n_329), .B1(n_456), .B2(n_454), .Y(n_716) );
INVx4_ASAP7_75t_L g717 ( .A(n_556), .Y(n_717) );
NOR3xp33_ASAP7_75t_L g718 ( .A(n_564), .B(n_19), .C(n_20), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_610), .B(n_20), .Y(n_719) );
O2A1O1Ixp33_ASAP7_75t_L g720 ( .A1(n_617), .A2(n_25), .B(n_21), .C(n_22), .Y(n_720) );
BUFx6f_ASAP7_75t_L g721 ( .A(n_609), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_614), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_616), .B(n_21), .Y(n_723) );
NAND2xp5_ASAP7_75t_SL g724 ( .A(n_590), .B(n_456), .Y(n_724) );
NAND2xp5_ASAP7_75t_SL g725 ( .A(n_624), .B(n_456), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_554), .Y(n_726) );
AOI21x1_ASAP7_75t_L g727 ( .A1(n_626), .A2(n_522), .B(n_464), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_625), .B(n_22), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_614), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_607), .B(n_25), .Y(n_730) );
AND2x2_ASAP7_75t_L g731 ( .A(n_607), .B(n_26), .Y(n_731) );
BUFx8_ASAP7_75t_L g732 ( .A(n_611), .Y(n_732) );
OA22x2_ASAP7_75t_L g733 ( .A1(n_545), .A2(n_29), .B1(n_27), .B2(n_28), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g734 ( .A1(n_608), .A2(n_484), .B1(n_464), .B2(n_31), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_608), .B(n_29), .Y(n_735) );
NAND2xp5_ASAP7_75t_SL g736 ( .A(n_578), .B(n_484), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g737 ( .A(n_578), .B(n_484), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_612), .B(n_30), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_604), .Y(n_739) );
O2A1O1Ixp33_ASAP7_75t_SL g740 ( .A1(n_571), .A2(n_145), .B(n_281), .C(n_280), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_551), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_546), .A2(n_30), .B1(n_31), .B2(n_32), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_565), .B(n_32), .Y(n_743) );
O2A1O1Ixp33_ASAP7_75t_L g744 ( .A1(n_561), .A2(n_33), .B(n_34), .C(n_35), .Y(n_744) );
OAI321xp33_ASAP7_75t_L g745 ( .A1(n_551), .A2(n_34), .A3(n_39), .B1(n_40), .B2(n_41), .C(n_42), .Y(n_745) );
CKINVDCx5p33_ASAP7_75t_R g746 ( .A(n_569), .Y(n_746) );
OAI21xp5_ASAP7_75t_L g747 ( .A1(n_566), .A2(n_95), .B(n_94), .Y(n_747) );
A2O1A1Ixp33_ASAP7_75t_L g748 ( .A1(n_544), .A2(n_42), .B(n_43), .C(n_44), .Y(n_748) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_623), .Y(n_749) );
OAI21xp5_ASAP7_75t_L g750 ( .A1(n_566), .A2(n_97), .B(n_96), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_605), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g752 ( .A(n_541), .B(n_44), .Y(n_752) );
O2A1O1Ixp33_ASAP7_75t_L g753 ( .A1(n_561), .A2(n_45), .B(n_46), .C(n_47), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_584), .A2(n_46), .B1(n_48), .B2(n_49), .Y(n_754) );
O2A1O1Ixp33_ASAP7_75t_L g755 ( .A1(n_561), .A2(n_48), .B(n_50), .C(n_51), .Y(n_755) );
AO21x1_ASAP7_75t_L g756 ( .A1(n_747), .A2(n_101), .B(n_100), .Y(n_756) );
OAI22x1_ASAP7_75t_L g757 ( .A1(n_754), .A2(n_50), .B1(n_51), .B2(n_52), .Y(n_757) );
NAND3x1_ASAP7_75t_L g758 ( .A(n_704), .B(n_53), .C(n_54), .Y(n_758) );
OAI21xp5_ASAP7_75t_L g759 ( .A1(n_631), .A2(n_106), .B(n_103), .Y(n_759) );
AOI221xp5_ASAP7_75t_SL g760 ( .A1(n_672), .A2(n_53), .B1(n_54), .B2(n_55), .C(n_56), .Y(n_760) );
BUFx2_ASAP7_75t_L g761 ( .A(n_732), .Y(n_761) );
AO31x2_ASAP7_75t_L g762 ( .A1(n_714), .A2(n_55), .A3(n_57), .B(n_58), .Y(n_762) );
OAI22x1_ASAP7_75t_L g763 ( .A1(n_705), .A2(n_59), .B1(n_60), .B2(n_61), .Y(n_763) );
AO22x2_ASAP7_75t_L g764 ( .A1(n_683), .A2(n_59), .B1(n_60), .B2(n_61), .Y(n_764) );
CKINVDCx12_ASAP7_75t_R g765 ( .A(n_627), .Y(n_765) );
BUFx10_ASAP7_75t_L g766 ( .A(n_746), .Y(n_766) );
INVxp67_ASAP7_75t_SL g767 ( .A(n_732), .Y(n_767) );
AOI21xp5_ASAP7_75t_L g768 ( .A1(n_647), .A2(n_176), .B(n_279), .Y(n_768) );
AOI21xp5_ASAP7_75t_L g769 ( .A1(n_647), .A2(n_175), .B(n_276), .Y(n_769) );
AO22x1_ASAP7_75t_L g770 ( .A1(n_635), .A2(n_63), .B1(n_64), .B2(n_65), .Y(n_770) );
BUFx3_ASAP7_75t_L g771 ( .A(n_629), .Y(n_771) );
AOI21xp5_ASAP7_75t_L g772 ( .A1(n_725), .A2(n_177), .B(n_273), .Y(n_772) );
INVx3_ASAP7_75t_L g773 ( .A(n_702), .Y(n_773) );
AOI21xp5_ASAP7_75t_L g774 ( .A1(n_724), .A2(n_166), .B(n_267), .Y(n_774) );
OAI21xp33_ASAP7_75t_SL g775 ( .A1(n_682), .A2(n_66), .B(n_67), .Y(n_775) );
AO31x2_ASAP7_75t_L g776 ( .A1(n_715), .A2(n_69), .A3(n_70), .B(n_71), .Y(n_776) );
BUFx3_ASAP7_75t_L g777 ( .A(n_655), .Y(n_777) );
O2A1O1Ixp33_ASAP7_75t_SL g778 ( .A1(n_736), .A2(n_737), .B(n_750), .C(n_747), .Y(n_778) );
AO31x2_ASAP7_75t_L g779 ( .A1(n_681), .A2(n_71), .A3(n_73), .B(n_75), .Y(n_779) );
AOI21xp5_ASAP7_75t_L g780 ( .A1(n_661), .A2(n_178), .B(n_266), .Y(n_780) );
AOI21xp5_ASAP7_75t_L g781 ( .A1(n_662), .A2(n_663), .B(n_743), .Y(n_781) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_639), .A2(n_75), .B1(n_76), .B2(n_77), .Y(n_782) );
BUFx6f_ASAP7_75t_L g783 ( .A(n_655), .Y(n_783) );
OAI22xp5_ASAP7_75t_L g784 ( .A1(n_665), .A2(n_78), .B1(n_79), .B2(n_80), .Y(n_784) );
AOI22xp33_ASAP7_75t_SL g785 ( .A1(n_650), .A2(n_79), .B1(n_81), .B2(n_82), .Y(n_785) );
CKINVDCx11_ASAP7_75t_R g786 ( .A(n_692), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_741), .B(n_81), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_627), .A2(n_119), .B1(n_120), .B2(n_123), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_726), .Y(n_789) );
OR2x2_ASAP7_75t_L g790 ( .A(n_632), .B(n_125), .Y(n_790) );
BUFx6f_ASAP7_75t_L g791 ( .A(n_655), .Y(n_791) );
AOI221x1_ASAP7_75t_L g792 ( .A1(n_681), .A2(n_128), .B1(n_129), .B2(n_130), .C(n_131), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_718), .A2(n_132), .B1(n_133), .B2(n_135), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_713), .Y(n_794) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_749), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_657), .B(n_136), .Y(n_796) );
CKINVDCx9p33_ASAP7_75t_R g797 ( .A(n_728), .Y(n_797) );
OAI21xp5_ASAP7_75t_L g798 ( .A1(n_641), .A2(n_138), .B(n_139), .Y(n_798) );
NOR2xp33_ASAP7_75t_L g799 ( .A(n_651), .B(n_144), .Y(n_799) );
A2O1A1Ixp33_ASAP7_75t_L g800 ( .A1(n_648), .A2(n_146), .B(n_147), .C(n_149), .Y(n_800) );
A2O1A1Ixp33_ASAP7_75t_L g801 ( .A1(n_678), .A2(n_150), .B(n_151), .C(n_152), .Y(n_801) );
INVx4_ASAP7_75t_L g802 ( .A(n_700), .Y(n_802) );
AOI221x1_ASAP7_75t_L g803 ( .A1(n_742), .A2(n_154), .B1(n_155), .B2(n_156), .C(n_157), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_719), .Y(n_804) );
OR2x2_ASAP7_75t_L g805 ( .A(n_634), .B(n_165), .Y(n_805) );
AOI21xp5_ASAP7_75t_L g806 ( .A1(n_671), .A2(n_180), .B(n_184), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_723), .Y(n_807) );
AOI21xp5_ASAP7_75t_L g808 ( .A1(n_687), .A2(n_191), .B(n_193), .Y(n_808) );
CKINVDCx5p33_ASAP7_75t_R g809 ( .A(n_668), .Y(n_809) );
BUFx3_ASAP7_75t_L g810 ( .A(n_717), .Y(n_810) );
CKINVDCx11_ASAP7_75t_R g811 ( .A(n_695), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_649), .B(n_195), .Y(n_812) );
OR2x2_ASAP7_75t_L g813 ( .A(n_652), .B(n_196), .Y(n_813) );
A2O1A1Ixp33_ASAP7_75t_L g814 ( .A1(n_677), .A2(n_197), .B(n_199), .C(n_200), .Y(n_814) );
NOR2xp67_ASAP7_75t_L g815 ( .A(n_666), .B(n_201), .Y(n_815) );
BUFx3_ASAP7_75t_L g816 ( .A(n_694), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g817 ( .A(n_695), .Y(n_817) );
AOI211x1_ASAP7_75t_L g818 ( .A1(n_628), .A2(n_204), .B(n_212), .C(n_213), .Y(n_818) );
OAI21xp33_ASAP7_75t_SL g819 ( .A1(n_730), .A2(n_735), .B(n_731), .Y(n_819) );
NOR2xp67_ASAP7_75t_L g820 ( .A(n_688), .B(n_215), .Y(n_820) );
OR2x2_ASAP7_75t_L g821 ( .A(n_658), .B(n_216), .Y(n_821) );
BUFx3_ASAP7_75t_L g822 ( .A(n_694), .Y(n_822) );
O2A1O1Ixp33_ASAP7_75t_L g823 ( .A1(n_748), .A2(n_217), .B(n_220), .C(n_223), .Y(n_823) );
AOI21xp5_ASAP7_75t_L g824 ( .A1(n_711), .A2(n_224), .B(n_227), .Y(n_824) );
AOI31xp67_ASAP7_75t_L g825 ( .A1(n_712), .A2(n_230), .A3(n_231), .B(n_235), .Y(n_825) );
INVx1_ASAP7_75t_SL g826 ( .A(n_752), .Y(n_826) );
NAND4xp25_ASAP7_75t_L g827 ( .A(n_640), .B(n_236), .C(n_241), .D(n_243), .Y(n_827) );
OAI21xp5_ASAP7_75t_L g828 ( .A1(n_653), .A2(n_245), .B(n_248), .Y(n_828) );
AOI21xp5_ASAP7_75t_L g829 ( .A1(n_701), .A2(n_249), .B(n_255), .Y(n_829) );
AND2x2_ASAP7_75t_L g830 ( .A(n_664), .B(n_257), .Y(n_830) );
HB1xp67_ASAP7_75t_L g831 ( .A(n_633), .Y(n_831) );
BUFx6f_ASAP7_75t_L g832 ( .A(n_721), .Y(n_832) );
O2A1O1Ixp33_ASAP7_75t_SL g833 ( .A1(n_738), .A2(n_259), .B(n_264), .C(n_689), .Y(n_833) );
BUFx2_ASAP7_75t_L g834 ( .A(n_751), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_679), .B(n_637), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_699), .Y(n_836) );
O2A1O1Ixp33_ASAP7_75t_L g837 ( .A1(n_654), .A2(n_755), .B(n_753), .C(n_744), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_733), .Y(n_838) );
OR2x2_ASAP7_75t_L g839 ( .A(n_667), .B(n_698), .Y(n_839) );
BUFx6f_ASAP7_75t_L g840 ( .A(n_721), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_638), .B(n_642), .Y(n_841) );
NAND3xp33_ASAP7_75t_L g842 ( .A(n_710), .B(n_734), .C(n_693), .Y(n_842) );
AOI21xp5_ASAP7_75t_L g843 ( .A1(n_669), .A2(n_670), .B(n_643), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_680), .B(n_674), .Y(n_844) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_680), .A2(n_675), .B1(n_676), .B2(n_660), .Y(n_845) );
OAI22xp5_ASAP7_75t_L g846 ( .A1(n_721), .A2(n_722), .B1(n_729), .B2(n_645), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_720), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_646), .B(n_707), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_690), .B(n_659), .Y(n_849) );
AO31x2_ASAP7_75t_L g850 ( .A1(n_685), .A2(n_716), .A3(n_739), .B(n_691), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_697), .Y(n_851) );
O2A1O1Ixp33_ASAP7_75t_L g852 ( .A1(n_686), .A2(n_745), .B(n_630), .C(n_706), .Y(n_852) );
OAI21x1_ASAP7_75t_L g853 ( .A1(n_708), .A2(n_740), .B(n_745), .Y(n_853) );
NOR2xp33_ASAP7_75t_SL g854 ( .A(n_708), .B(n_732), .Y(n_854) );
A2O1A1Ixp33_ASAP7_75t_L g855 ( .A1(n_672), .A2(n_673), .B(n_709), .C(n_703), .Y(n_855) );
INVx2_ASAP7_75t_SL g856 ( .A(n_732), .Y(n_856) );
AOI21xp5_ASAP7_75t_L g857 ( .A1(n_636), .A2(n_566), .B(n_571), .Y(n_857) );
AOI21xp5_ASAP7_75t_L g858 ( .A1(n_636), .A2(n_566), .B(n_571), .Y(n_858) );
AOI21xp5_ASAP7_75t_L g859 ( .A1(n_636), .A2(n_566), .B(n_571), .Y(n_859) );
CKINVDCx11_ASAP7_75t_R g860 ( .A(n_629), .Y(n_860) );
INVx3_ASAP7_75t_L g861 ( .A(n_702), .Y(n_861) );
CKINVDCx11_ASAP7_75t_R g862 ( .A(n_629), .Y(n_862) );
NAND2x1p5_ASAP7_75t_L g863 ( .A(n_629), .B(n_700), .Y(n_863) );
NAND3xp33_ASAP7_75t_SL g864 ( .A(n_635), .B(n_644), .C(n_564), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_656), .Y(n_865) );
NOR4xp25_ASAP7_75t_L g866 ( .A(n_745), .B(n_742), .C(n_678), .D(n_744), .Y(n_866) );
AO31x2_ASAP7_75t_L g867 ( .A1(n_636), .A2(n_631), .A3(n_613), .B(n_615), .Y(n_867) );
BUFx2_ASAP7_75t_R g868 ( .A(n_746), .Y(n_868) );
INVx4_ASAP7_75t_L g869 ( .A(n_700), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_656), .Y(n_870) );
INVx3_ASAP7_75t_SL g871 ( .A(n_746), .Y(n_871) );
NAND3xp33_ASAP7_75t_L g872 ( .A(n_635), .B(n_550), .C(n_651), .Y(n_872) );
A2O1A1Ixp33_ASAP7_75t_L g873 ( .A1(n_672), .A2(n_673), .B(n_709), .C(n_703), .Y(n_873) );
NAND3xp33_ASAP7_75t_SL g874 ( .A(n_635), .B(n_644), .C(n_564), .Y(n_874) );
NAND2xp5_ASAP7_75t_SL g875 ( .A(n_684), .B(n_505), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_709), .A2(n_546), .B1(n_598), .B2(n_555), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_709), .B(n_584), .Y(n_877) );
INVx1_ASAP7_75t_SL g878 ( .A(n_629), .Y(n_878) );
AOI21xp5_ASAP7_75t_L g879 ( .A1(n_636), .A2(n_566), .B(n_571), .Y(n_879) );
AND2x4_ASAP7_75t_L g880 ( .A(n_682), .B(n_656), .Y(n_880) );
AND2x2_ASAP7_75t_L g881 ( .A(n_696), .B(n_584), .Y(n_881) );
A2O1A1Ixp33_ASAP7_75t_L g882 ( .A1(n_672), .A2(n_673), .B(n_709), .C(n_703), .Y(n_882) );
NOR2xp67_ASAP7_75t_SL g883 ( .A(n_639), .B(n_569), .Y(n_883) );
AOI21xp5_ASAP7_75t_L g884 ( .A1(n_636), .A2(n_566), .B(n_571), .Y(n_884) );
NOR2x1_ASAP7_75t_SL g885 ( .A(n_695), .B(n_623), .Y(n_885) );
OAI21x1_ASAP7_75t_L g886 ( .A1(n_727), .A2(n_613), .B(n_566), .Y(n_886) );
BUFx4_ASAP7_75t_SL g887 ( .A(n_746), .Y(n_887) );
OR2x6_ASAP7_75t_L g888 ( .A(n_629), .B(n_627), .Y(n_888) );
AND2x6_ASAP7_75t_L g889 ( .A(n_700), .B(n_682), .Y(n_889) );
AOI21xp5_ASAP7_75t_L g890 ( .A1(n_636), .A2(n_566), .B(n_571), .Y(n_890) );
AND2x4_ASAP7_75t_L g891 ( .A(n_682), .B(n_656), .Y(n_891) );
OAI21xp5_ASAP7_75t_SL g892 ( .A1(n_635), .A2(n_594), .B(n_595), .Y(n_892) );
OAI21x1_ASAP7_75t_L g893 ( .A1(n_727), .A2(n_613), .B(n_566), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_877), .B(n_865), .Y(n_894) );
AND2x4_ASAP7_75t_L g895 ( .A(n_880), .B(n_891), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_870), .B(n_881), .Y(n_896) );
BUFx8_ASAP7_75t_L g897 ( .A(n_761), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_892), .B(n_880), .Y(n_898) );
INVx4_ASAP7_75t_L g899 ( .A(n_889), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_891), .B(n_876), .Y(n_900) );
CKINVDCx20_ASAP7_75t_R g901 ( .A(n_860), .Y(n_901) );
AO21x2_ASAP7_75t_L g902 ( .A1(n_778), .A2(n_853), .B(n_759), .Y(n_902) );
AO31x2_ASAP7_75t_L g903 ( .A1(n_756), .A2(n_890), .A3(n_884), .B(n_857), .Y(n_903) );
AO21x2_ASAP7_75t_L g904 ( .A1(n_879), .A2(n_852), .B(n_833), .Y(n_904) );
INVx2_ASAP7_75t_L g905 ( .A(n_789), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_789), .Y(n_906) );
OAI21xp5_ASAP7_75t_L g907 ( .A1(n_872), .A2(n_873), .B(n_855), .Y(n_907) );
NOR2xp33_ASAP7_75t_SL g908 ( .A(n_868), .B(n_767), .Y(n_908) );
INVx3_ASAP7_75t_L g909 ( .A(n_889), .Y(n_909) );
AOI21xp5_ASAP7_75t_L g910 ( .A1(n_819), .A2(n_781), .B(n_882), .Y(n_910) );
BUFx2_ASAP7_75t_L g911 ( .A(n_771), .Y(n_911) );
NOR2x1_ASAP7_75t_SL g912 ( .A(n_783), .B(n_791), .Y(n_912) );
NOR2xp33_ASAP7_75t_L g913 ( .A(n_864), .B(n_874), .Y(n_913) );
INVx4_ASAP7_75t_SL g914 ( .A(n_871), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_839), .B(n_835), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_838), .Y(n_916) );
INVx3_ASAP7_75t_L g917 ( .A(n_889), .Y(n_917) );
AND2x4_ASAP7_75t_L g918 ( .A(n_889), .B(n_885), .Y(n_918) );
AOI21xp5_ASAP7_75t_L g919 ( .A1(n_843), .A2(n_837), .B(n_796), .Y(n_919) );
AO21x2_ASAP7_75t_L g920 ( .A1(n_842), .A2(n_866), .B(n_847), .Y(n_920) );
NAND2x1p5_ASAP7_75t_L g921 ( .A(n_856), .B(n_802), .Y(n_921) );
OA21x2_ASAP7_75t_L g922 ( .A1(n_803), .A2(n_792), .B(n_798), .Y(n_922) );
INVx3_ASAP7_75t_L g923 ( .A(n_810), .Y(n_923) );
AND2x2_ASAP7_75t_L g924 ( .A(n_764), .B(n_888), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_836), .Y(n_925) );
AND2x4_ASAP7_75t_L g926 ( .A(n_802), .B(n_869), .Y(n_926) );
BUFx2_ASAP7_75t_L g927 ( .A(n_888), .Y(n_927) );
AO31x2_ASAP7_75t_L g928 ( .A1(n_768), .A2(n_769), .A3(n_801), .B(n_814), .Y(n_928) );
AO31x2_ASAP7_75t_L g929 ( .A1(n_800), .A2(n_757), .A3(n_794), .B(n_807), .Y(n_929) );
OAI21x1_ASAP7_75t_SL g930 ( .A1(n_828), .A2(n_821), .B(n_813), .Y(n_930) );
AO31x2_ASAP7_75t_L g931 ( .A1(n_804), .A2(n_829), .A3(n_824), .B(n_799), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_787), .Y(n_932) );
AO31x2_ASAP7_75t_L g933 ( .A1(n_808), .A2(n_806), .A3(n_845), .B(n_846), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_779), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_795), .B(n_848), .Y(n_935) );
NAND3xp33_ASAP7_75t_L g936 ( .A(n_760), .B(n_818), .C(n_785), .Y(n_936) );
AO31x2_ASAP7_75t_L g937 ( .A1(n_780), .A2(n_772), .A3(n_782), .B(n_784), .Y(n_937) );
OA21x2_ASAP7_75t_L g938 ( .A1(n_774), .A2(n_827), .B(n_793), .Y(n_938) );
BUFx4f_ASAP7_75t_SL g939 ( .A(n_766), .Y(n_939) );
NAND2x1p5_ASAP7_75t_L g940 ( .A(n_869), .B(n_878), .Y(n_940) );
AOI21xp5_ASAP7_75t_L g941 ( .A1(n_805), .A2(n_849), .B(n_823), .Y(n_941) );
OA21x2_ASAP7_75t_L g942 ( .A1(n_812), .A2(n_815), .B(n_820), .Y(n_942) );
INVxp67_ASAP7_75t_L g943 ( .A(n_883), .Y(n_943) );
OA21x2_ASAP7_75t_L g944 ( .A1(n_867), .A2(n_844), .B(n_830), .Y(n_944) );
BUFx2_ASAP7_75t_L g945 ( .A(n_863), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_779), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_850), .Y(n_947) );
AOI21xp5_ASAP7_75t_L g948 ( .A1(n_875), .A2(n_841), .B(n_826), .Y(n_948) );
OAI21x1_ASAP7_75t_L g949 ( .A1(n_773), .A2(n_861), .B(n_788), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_790), .B(n_764), .Y(n_950) );
INVx3_ASAP7_75t_L g951 ( .A(n_777), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_851), .B(n_834), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_831), .B(n_822), .Y(n_953) );
AO21x2_ASAP7_75t_L g954 ( .A1(n_825), .A2(n_776), .B(n_762), .Y(n_954) );
INVx2_ASAP7_75t_L g955 ( .A(n_776), .Y(n_955) );
OA21x2_ASAP7_75t_L g956 ( .A1(n_776), .A2(n_762), .B(n_854), .Y(n_956) );
NOR2xp33_ASAP7_75t_L g957 ( .A(n_817), .B(n_765), .Y(n_957) );
AOI21xp5_ASAP7_75t_L g958 ( .A1(n_832), .A2(n_840), .B(n_775), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_762), .Y(n_959) );
AOI21x1_ASAP7_75t_L g960 ( .A1(n_770), .A2(n_763), .B(n_797), .Y(n_960) );
BUFx2_ASAP7_75t_R g961 ( .A(n_809), .Y(n_961) );
BUFx6f_ASAP7_75t_L g962 ( .A(n_832), .Y(n_962) );
INVx1_ASAP7_75t_L g963 ( .A(n_840), .Y(n_963) );
OAI21x1_ASAP7_75t_L g964 ( .A1(n_840), .A2(n_758), .B(n_816), .Y(n_964) );
INVx1_ASAP7_75t_L g965 ( .A(n_811), .Y(n_965) );
OAI21x1_ASAP7_75t_SL g966 ( .A1(n_786), .A2(n_887), .B(n_862), .Y(n_966) );
CKINVDCx6p67_ASAP7_75t_R g967 ( .A(n_766), .Y(n_967) );
AND2x2_ASAP7_75t_L g968 ( .A(n_881), .B(n_696), .Y(n_968) );
A2O1A1Ixp33_ASAP7_75t_L g969 ( .A1(n_819), .A2(n_837), .B(n_872), .C(n_855), .Y(n_969) );
AOI21xp5_ASAP7_75t_L g970 ( .A1(n_778), .A2(n_858), .B(n_857), .Y(n_970) );
CKINVDCx5p33_ASAP7_75t_R g971 ( .A(n_887), .Y(n_971) );
AO31x2_ASAP7_75t_L g972 ( .A1(n_756), .A2(n_858), .A3(n_859), .B(n_857), .Y(n_972) );
AOI21xp5_ASAP7_75t_L g973 ( .A1(n_778), .A2(n_858), .B(n_857), .Y(n_973) );
INVx2_ASAP7_75t_SL g974 ( .A(n_761), .Y(n_974) );
OR2x2_ASAP7_75t_L g975 ( .A(n_881), .B(n_696), .Y(n_975) );
HB1xp67_ASAP7_75t_L g976 ( .A(n_761), .Y(n_976) );
AO21x2_ASAP7_75t_L g977 ( .A1(n_778), .A2(n_853), .B(n_857), .Y(n_977) );
NOR2xp33_ASAP7_75t_L g978 ( .A(n_892), .B(n_872), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_789), .Y(n_979) );
AND2x2_ASAP7_75t_L g980 ( .A(n_881), .B(n_696), .Y(n_980) );
CKINVDCx20_ASAP7_75t_R g981 ( .A(n_860), .Y(n_981) );
INVx4_ASAP7_75t_L g982 ( .A(n_889), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_877), .B(n_584), .Y(n_983) );
INVx1_ASAP7_75t_L g984 ( .A(n_789), .Y(n_984) );
AO31x2_ASAP7_75t_L g985 ( .A1(n_756), .A2(n_858), .A3(n_859), .B(n_857), .Y(n_985) );
OA21x2_ASAP7_75t_L g986 ( .A1(n_853), .A2(n_893), .B(n_886), .Y(n_986) );
NAND2x1p5_ASAP7_75t_L g987 ( .A(n_761), .B(n_856), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_789), .Y(n_988) );
OR2x2_ASAP7_75t_L g989 ( .A(n_881), .B(n_696), .Y(n_989) );
AOI21xp5_ASAP7_75t_L g990 ( .A1(n_778), .A2(n_858), .B(n_857), .Y(n_990) );
HB1xp67_ASAP7_75t_L g991 ( .A(n_761), .Y(n_991) );
INVx4_ASAP7_75t_L g992 ( .A(n_889), .Y(n_992) );
INVx2_ASAP7_75t_L g993 ( .A(n_865), .Y(n_993) );
OR2x2_ASAP7_75t_L g994 ( .A(n_881), .B(n_696), .Y(n_994) );
AOI21xp5_ASAP7_75t_L g995 ( .A1(n_778), .A2(n_858), .B(n_857), .Y(n_995) );
AOI21xp5_ASAP7_75t_L g996 ( .A1(n_778), .A2(n_858), .B(n_857), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_877), .B(n_584), .Y(n_997) );
OAI21xp5_ASAP7_75t_L g998 ( .A1(n_872), .A2(n_873), .B(n_855), .Y(n_998) );
NOR2xp33_ASAP7_75t_L g999 ( .A(n_892), .B(n_872), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g1000 ( .A(n_877), .B(n_584), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_881), .B(n_696), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_877), .B(n_584), .Y(n_1002) );
OR2x6_ASAP7_75t_L g1003 ( .A(n_761), .B(n_856), .Y(n_1003) );
NAND3xp33_ASAP7_75t_L g1004 ( .A(n_872), .B(n_760), .C(n_819), .Y(n_1004) );
A2O1A1Ixp33_ASAP7_75t_L g1005 ( .A1(n_819), .A2(n_837), .B(n_872), .C(n_855), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_789), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_789), .Y(n_1007) );
NAND2x1p5_ASAP7_75t_L g1008 ( .A(n_761), .B(n_856), .Y(n_1008) );
HB1xp67_ASAP7_75t_L g1009 ( .A(n_761), .Y(n_1009) );
NAND2x1p5_ASAP7_75t_L g1010 ( .A(n_761), .B(n_856), .Y(n_1010) );
NAND2x1p5_ASAP7_75t_L g1011 ( .A(n_761), .B(n_856), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_915), .B(n_983), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_905), .B(n_925), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_997), .B(n_1000), .Y(n_1014) );
AND2x4_ASAP7_75t_SL g1015 ( .A(n_899), .B(n_982), .Y(n_1015) );
INVx2_ASAP7_75t_L g1016 ( .A(n_906), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_993), .Y(n_1017) );
HB1xp67_ASAP7_75t_L g1018 ( .A(n_911), .Y(n_1018) );
HB1xp67_ASAP7_75t_L g1019 ( .A(n_895), .Y(n_1019) );
OR2x2_ASAP7_75t_L g1020 ( .A(n_975), .B(n_989), .Y(n_1020) );
HB1xp67_ASAP7_75t_L g1021 ( .A(n_895), .Y(n_1021) );
OR2x2_ASAP7_75t_L g1022 ( .A(n_994), .B(n_896), .Y(n_1022) );
OAI22xp33_ASAP7_75t_L g1023 ( .A1(n_950), .A2(n_908), .B1(n_992), .B2(n_899), .Y(n_1023) );
OR2x6_ASAP7_75t_L g1024 ( .A(n_982), .B(n_992), .Y(n_1024) );
OA21x2_ASAP7_75t_L g1025 ( .A1(n_970), .A2(n_990), .B(n_973), .Y(n_1025) );
BUFx2_ASAP7_75t_L g1026 ( .A(n_926), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_906), .B(n_979), .Y(n_1027) );
OA21x2_ASAP7_75t_L g1028 ( .A1(n_995), .A2(n_996), .B(n_910), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_978), .A2(n_999), .B1(n_913), .B2(n_898), .Y(n_1029) );
INVx2_ASAP7_75t_L g1030 ( .A(n_979), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_984), .B(n_988), .Y(n_1031) );
INVx4_ASAP7_75t_L g1032 ( .A(n_918), .Y(n_1032) );
INVx2_ASAP7_75t_L g1033 ( .A(n_984), .Y(n_1033) );
BUFx2_ASAP7_75t_L g1034 ( .A(n_926), .Y(n_1034) );
INVx1_ASAP7_75t_SL g1035 ( .A(n_945), .Y(n_1035) );
AND2x4_ASAP7_75t_L g1036 ( .A(n_918), .B(n_909), .Y(n_1036) );
BUFx3_ASAP7_75t_L g1037 ( .A(n_921), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_1006), .B(n_1007), .Y(n_1038) );
OAI211xp5_ASAP7_75t_SL g1039 ( .A1(n_965), .A2(n_1002), .B(n_935), .C(n_894), .Y(n_1039) );
BUFx2_ASAP7_75t_L g1040 ( .A(n_1003), .Y(n_1040) );
AOI322xp5_ASAP7_75t_L g1041 ( .A1(n_924), .A2(n_981), .A3(n_901), .B1(n_980), .B2(n_968), .C1(n_1001), .C2(n_965), .Y(n_1041) );
AO21x1_ASAP7_75t_SL g1042 ( .A1(n_900), .A2(n_963), .B(n_953), .Y(n_1042) );
INVx2_ASAP7_75t_L g1043 ( .A(n_947), .Y(n_1043) );
BUFx4f_ASAP7_75t_L g1044 ( .A(n_917), .Y(n_1044) );
OR2x2_ASAP7_75t_L g1045 ( .A(n_916), .B(n_934), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_952), .Y(n_1046) );
INVx1_ASAP7_75t_L g1047 ( .A(n_916), .Y(n_1047) );
HB1xp67_ASAP7_75t_L g1048 ( .A(n_940), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_932), .B(n_907), .Y(n_1049) );
INVx2_ASAP7_75t_SL g1050 ( .A(n_987), .Y(n_1050) );
INVx2_ASAP7_75t_L g1051 ( .A(n_986), .Y(n_1051) );
BUFx3_ASAP7_75t_L g1052 ( .A(n_1008), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_934), .Y(n_1053) );
INVx2_ASAP7_75t_SL g1054 ( .A(n_1010), .Y(n_1054) );
OAI21xp5_ASAP7_75t_L g1055 ( .A1(n_936), .A2(n_941), .B(n_969), .Y(n_1055) );
OR2x6_ASAP7_75t_L g1056 ( .A(n_964), .B(n_930), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_946), .Y(n_1057) );
OR2x2_ASAP7_75t_L g1058 ( .A(n_920), .B(n_959), .Y(n_1058) );
AND2x4_ASAP7_75t_L g1059 ( .A(n_912), .B(n_949), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_932), .B(n_998), .Y(n_1060) );
BUFx2_ASAP7_75t_L g1061 ( .A(n_897), .Y(n_1061) );
INVx1_ASAP7_75t_L g1062 ( .A(n_923), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_923), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_1005), .B(n_929), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_1004), .A2(n_927), .B1(n_944), .B2(n_959), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_944), .A2(n_991), .B1(n_1009), .B2(n_976), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_929), .B(n_955), .Y(n_1067) );
AO21x2_ASAP7_75t_L g1068 ( .A1(n_919), .A2(n_954), .B(n_977), .Y(n_1068) );
HB1xp67_ASAP7_75t_L g1069 ( .A(n_974), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_960), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_929), .B(n_912), .Y(n_1071) );
BUFx3_ASAP7_75t_L g1072 ( .A(n_1011), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_943), .Y(n_1073) );
OR2x2_ASAP7_75t_L g1074 ( .A(n_956), .B(n_951), .Y(n_1074) );
INVx1_ASAP7_75t_L g1075 ( .A(n_951), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_954), .B(n_956), .Y(n_1076) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_942), .A2(n_957), .B1(n_948), .B2(n_922), .Y(n_1077) );
AND2x4_ASAP7_75t_L g1078 ( .A(n_962), .B(n_958), .Y(n_1078) );
OR2x2_ASAP7_75t_L g1079 ( .A(n_903), .B(n_985), .Y(n_1079) );
HB1xp67_ASAP7_75t_L g1080 ( .A(n_914), .Y(n_1080) );
AOI21xp5_ASAP7_75t_L g1081 ( .A1(n_904), .A2(n_922), .B(n_938), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_962), .B(n_937), .Y(n_1082) );
INVx5_ASAP7_75t_L g1083 ( .A(n_1024), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1053), .Y(n_1084) );
INVx6_ASAP7_75t_L g1085 ( .A(n_1032), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_1027), .B(n_985), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_1027), .B(n_985), .Y(n_1087) );
INVx2_ASAP7_75t_L g1088 ( .A(n_1043), .Y(n_1088) );
HB1xp67_ASAP7_75t_L g1089 ( .A(n_1018), .Y(n_1089) );
AND2x4_ASAP7_75t_L g1090 ( .A(n_1082), .B(n_972), .Y(n_1090) );
BUFx8_ASAP7_75t_L g1091 ( .A(n_1061), .Y(n_1091) );
HB1xp67_ASAP7_75t_L g1092 ( .A(n_1026), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_1031), .B(n_972), .Y(n_1093) );
INVx2_ASAP7_75t_SL g1094 ( .A(n_1032), .Y(n_1094) );
NAND2xp5_ASAP7_75t_L g1095 ( .A(n_1049), .B(n_967), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_1031), .B(n_972), .Y(n_1096) );
INVx2_ASAP7_75t_SL g1097 ( .A(n_1032), .Y(n_1097) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1057), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1099 ( .A(n_1049), .B(n_937), .Y(n_1099) );
BUFx3_ASAP7_75t_L g1100 ( .A(n_1034), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1038), .B(n_902), .Y(n_1101) );
BUFx2_ASAP7_75t_L g1102 ( .A(n_1059), .Y(n_1102) );
NAND2xp5_ASAP7_75t_L g1103 ( .A(n_1060), .B(n_937), .Y(n_1103) );
INVx2_ASAP7_75t_L g1104 ( .A(n_1051), .Y(n_1104) );
NAND2xp33_ASAP7_75t_SL g1105 ( .A(n_1080), .B(n_971), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_1064), .B(n_933), .Y(n_1106) );
NAND2xp5_ASAP7_75t_L g1107 ( .A(n_1060), .B(n_939), .Y(n_1107) );
OR2x2_ASAP7_75t_L g1108 ( .A(n_1045), .B(n_931), .Y(n_1108) );
HB1xp67_ASAP7_75t_L g1109 ( .A(n_1048), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1016), .Y(n_1110) );
HB1xp67_ASAP7_75t_L g1111 ( .A(n_1013), .Y(n_1111) );
NOR2xp33_ASAP7_75t_L g1112 ( .A(n_1012), .B(n_961), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_1016), .B(n_931), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1030), .B(n_931), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1033), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_1029), .B(n_966), .Y(n_1116) );
AND2x4_ASAP7_75t_L g1117 ( .A(n_1082), .B(n_928), .Y(n_1117) );
AND2x4_ASAP7_75t_L g1118 ( .A(n_1071), .B(n_1078), .Y(n_1118) );
INVx2_ASAP7_75t_L g1119 ( .A(n_1025), .Y(n_1119) );
INVx5_ASAP7_75t_L g1120 ( .A(n_1024), .Y(n_1120) );
AOI22xp5_ASAP7_75t_L g1121 ( .A1(n_1029), .A2(n_1039), .B1(n_1014), .B2(n_1046), .Y(n_1121) );
AND2x4_ASAP7_75t_L g1122 ( .A(n_1071), .B(n_1056), .Y(n_1122) );
BUFx2_ASAP7_75t_SL g1123 ( .A(n_1083), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_1086), .B(n_1067), .Y(n_1124) );
HB1xp67_ASAP7_75t_L g1125 ( .A(n_1089), .Y(n_1125) );
NOR3xp33_ASAP7_75t_L g1126 ( .A(n_1116), .B(n_1073), .C(n_1070), .Y(n_1126) );
INVx2_ASAP7_75t_L g1127 ( .A(n_1104), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1087), .B(n_1066), .Y(n_1128) );
AND2x4_ASAP7_75t_L g1129 ( .A(n_1118), .B(n_1056), .Y(n_1129) );
HB1xp67_ASAP7_75t_L g1130 ( .A(n_1092), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_1087), .B(n_1058), .Y(n_1131) );
BUFx2_ASAP7_75t_L g1132 ( .A(n_1102), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_1093), .B(n_1076), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_1096), .B(n_1076), .Y(n_1134) );
NAND2xp5_ASAP7_75t_SL g1135 ( .A(n_1083), .B(n_1023), .Y(n_1135) );
OR2x2_ASAP7_75t_L g1136 ( .A(n_1111), .B(n_1079), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g1137 ( .A(n_1096), .B(n_1066), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1084), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1084), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1106), .B(n_1065), .Y(n_1140) );
NOR2x1_ASAP7_75t_L g1141 ( .A(n_1100), .B(n_1037), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1106), .B(n_1065), .Y(n_1142) );
BUFx2_ASAP7_75t_L g1143 ( .A(n_1102), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1101), .B(n_1074), .Y(n_1144) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_1121), .A2(n_1021), .B1(n_1019), .B2(n_1042), .Y(n_1145) );
BUFx3_ASAP7_75t_L g1146 ( .A(n_1085), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1101), .B(n_1068), .Y(n_1147) );
BUFx2_ASAP7_75t_SL g1148 ( .A(n_1083), .Y(n_1148) );
OR2x2_ASAP7_75t_L g1149 ( .A(n_1099), .B(n_1020), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_1090), .B(n_1047), .Y(n_1150) );
INVxp67_ASAP7_75t_L g1151 ( .A(n_1109), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1090), .B(n_1077), .Y(n_1152) );
AOI21xp5_ASAP7_75t_L g1153 ( .A1(n_1119), .A2(n_1081), .B(n_1055), .Y(n_1153) );
OR2x2_ASAP7_75t_L g1154 ( .A(n_1103), .B(n_1022), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1117), .B(n_1028), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1138), .Y(n_1156) );
INVx2_ASAP7_75t_L g1157 ( .A(n_1127), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1138), .Y(n_1158) );
INVx2_ASAP7_75t_L g1159 ( .A(n_1127), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1139), .Y(n_1160) );
NAND2xp5_ASAP7_75t_L g1161 ( .A(n_1149), .B(n_1121), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1133), .B(n_1117), .Y(n_1162) );
NOR2x1_ASAP7_75t_L g1163 ( .A(n_1141), .B(n_1040), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1164 ( .A(n_1154), .B(n_1098), .Y(n_1164) );
OR2x2_ASAP7_75t_L g1165 ( .A(n_1136), .B(n_1108), .Y(n_1165) );
OR2x2_ASAP7_75t_L g1166 ( .A(n_1136), .B(n_1108), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1133), .B(n_1113), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1134), .B(n_1114), .Y(n_1168) );
INVxp67_ASAP7_75t_SL g1169 ( .A(n_1125), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1131), .B(n_1110), .Y(n_1170) );
CKINVDCx16_ASAP7_75t_R g1171 ( .A(n_1123), .Y(n_1171) );
OR2x2_ASAP7_75t_L g1172 ( .A(n_1131), .B(n_1088), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1144), .B(n_1122), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1124), .B(n_1122), .Y(n_1174) );
NAND2x1p5_ASAP7_75t_L g1175 ( .A(n_1135), .B(n_1083), .Y(n_1175) );
NAND2x1p5_ASAP7_75t_L g1176 ( .A(n_1146), .B(n_1083), .Y(n_1176) );
NOR2xp33_ASAP7_75t_L g1177 ( .A(n_1151), .B(n_1112), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_1130), .B(n_1115), .Y(n_1178) );
INVxp67_ASAP7_75t_L g1179 ( .A(n_1169), .Y(n_1179) );
NOR2x1_ASAP7_75t_L g1180 ( .A(n_1163), .B(n_1123), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1178), .Y(n_1181) );
INVx2_ASAP7_75t_L g1182 ( .A(n_1172), .Y(n_1182) );
INVx2_ASAP7_75t_SL g1183 ( .A(n_1171), .Y(n_1183) );
INVx2_ASAP7_75t_L g1184 ( .A(n_1157), .Y(n_1184) );
OR2x6_ASAP7_75t_L g1185 ( .A(n_1175), .B(n_1148), .Y(n_1185) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1156), .Y(n_1186) );
NOR2xp33_ASAP7_75t_L g1187 ( .A(n_1177), .B(n_1091), .Y(n_1187) );
INVx1_ASAP7_75t_SL g1188 ( .A(n_1170), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_1164), .B(n_1147), .Y(n_1189) );
AND2x4_ASAP7_75t_L g1190 ( .A(n_1174), .B(n_1129), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1158), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1160), .Y(n_1192) );
OAI221xp5_ASAP7_75t_SL g1193 ( .A1(n_1161), .A2(n_1041), .B1(n_1145), .B2(n_1095), .C(n_1107), .Y(n_1193) );
NAND2x1p5_ASAP7_75t_L g1194 ( .A(n_1176), .B(n_1120), .Y(n_1194) );
INVx2_ASAP7_75t_L g1195 ( .A(n_1159), .Y(n_1195) );
OAI21xp5_ASAP7_75t_L g1196 ( .A1(n_1179), .A2(n_1126), .B(n_1175), .Y(n_1196) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1186), .Y(n_1197) );
NAND2xp5_ASAP7_75t_L g1198 ( .A(n_1181), .B(n_1167), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1188), .B(n_1167), .Y(n_1199) );
NOR2xp33_ASAP7_75t_R g1200 ( .A(n_1183), .B(n_1105), .Y(n_1200) );
AOI211xp5_ASAP7_75t_SL g1201 ( .A1(n_1193), .A2(n_1137), .B(n_1128), .C(n_1152), .Y(n_1201) );
AOI22xp5_ASAP7_75t_L g1202 ( .A1(n_1189), .A2(n_1150), .B1(n_1162), .B2(n_1173), .Y(n_1202) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1191), .Y(n_1203) );
INVx2_ASAP7_75t_L g1204 ( .A(n_1184), .Y(n_1204) );
HB1xp67_ASAP7_75t_L g1205 ( .A(n_1195), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1182), .B(n_1168), .Y(n_1206) );
A2O1A1Ixp33_ASAP7_75t_L g1207 ( .A1(n_1201), .A2(n_1187), .B(n_1180), .C(n_1190), .Y(n_1207) );
AOI21xp5_ASAP7_75t_L g1208 ( .A1(n_1196), .A2(n_1185), .B(n_1194), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1197), .Y(n_1209) );
INVx1_ASAP7_75t_SL g1210 ( .A(n_1200), .Y(n_1210) );
OAI22xp5_ASAP7_75t_L g1211 ( .A1(n_1202), .A2(n_1176), .B1(n_1166), .B2(n_1165), .Y(n_1211) );
NOR3xp33_ASAP7_75t_L g1212 ( .A(n_1198), .B(n_1069), .C(n_1054), .Y(n_1212) );
AOI222xp33_ASAP7_75t_L g1213 ( .A1(n_1199), .A2(n_1091), .B1(n_1192), .B2(n_1142), .C1(n_1140), .C2(n_1155), .Y(n_1213) );
AOI21x1_ASAP7_75t_L g1214 ( .A1(n_1205), .A2(n_1143), .B(n_1132), .Y(n_1214) );
NOR3xp33_ASAP7_75t_L g1215 ( .A(n_1203), .B(n_1050), .C(n_1035), .Y(n_1215) );
AOI21xp33_ASAP7_75t_SL g1216 ( .A1(n_1206), .A2(n_1097), .B(n_1094), .Y(n_1216) );
NOR3xp33_ASAP7_75t_L g1217 ( .A(n_1204), .B(n_1063), .C(n_1062), .Y(n_1217) );
AOI21xp5_ASAP7_75t_L g1218 ( .A1(n_1204), .A2(n_1097), .B(n_1094), .Y(n_1218) );
OAI211xp5_ASAP7_75t_L g1219 ( .A1(n_1210), .A2(n_1207), .B(n_1208), .C(n_1213), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1209), .Y(n_1220) );
O2A1O1Ixp33_ASAP7_75t_L g1221 ( .A1(n_1215), .A2(n_1212), .B(n_1211), .C(n_1216), .Y(n_1221) );
NAND4xp25_ASAP7_75t_L g1222 ( .A(n_1219), .B(n_1052), .C(n_1072), .D(n_1037), .Y(n_1222) );
NOR3xp33_ASAP7_75t_L g1223 ( .A(n_1221), .B(n_1214), .C(n_1218), .Y(n_1223) );
NAND4xp25_ASAP7_75t_L g1224 ( .A(n_1222), .B(n_1072), .C(n_1052), .D(n_1220), .Y(n_1224) );
AND2x4_ASAP7_75t_L g1225 ( .A(n_1223), .B(n_1217), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1225), .Y(n_1226) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1226), .Y(n_1227) );
AOI22x1_ASAP7_75t_SL g1228 ( .A1(n_1227), .A2(n_1224), .B1(n_1075), .B2(n_1017), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1228), .Y(n_1229) );
XOR2x2_ASAP7_75t_L g1230 ( .A(n_1229), .B(n_1036), .Y(n_1230) );
AOI21xp5_ASAP7_75t_L g1231 ( .A1(n_1230), .A2(n_1044), .B(n_1015), .Y(n_1231) );
AOI21xp5_ASAP7_75t_L g1232 ( .A1(n_1231), .A2(n_1044), .B(n_1153), .Y(n_1232) );
endmodule