module real_jpeg_13344_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_297, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_297;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_233;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_249;
wire n_78;
wire n_286;
wire n_166;
wire n_221;
wire n_292;
wire n_176;
wire n_215;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_150;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_213;
wire n_179;
wire n_167;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;

BUFx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_3),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_3),
.B(n_38),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_3),
.B(n_162),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_3),
.A2(n_42),
.B(n_80),
.C(n_208),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_3),
.A2(n_59),
.B1(n_60),
.B2(n_133),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_3),
.B(n_29),
.C(n_63),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_3),
.B(n_81),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_L g247 ( 
.A1(n_3),
.A2(n_93),
.B(n_233),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_3),
.A2(n_42),
.B1(n_43),
.B2(n_133),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_6),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_6),
.A2(n_38),
.B1(n_39),
.B2(n_139),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_6),
.A2(n_59),
.B1(n_60),
.B2(n_139),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_139),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_7),
.A2(n_38),
.B1(n_39),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_7),
.A2(n_52),
.B1(n_59),
.B2(n_60),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_7),
.A2(n_42),
.B1(n_43),
.B2(n_52),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_52),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_8),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_8),
.A2(n_42),
.B1(n_43),
.B2(n_58),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_58),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_83),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_10),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_10),
.A2(n_59),
.B1(n_60),
.B2(n_83),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_83),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_83),
.Y(n_153)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_11),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_12),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_41)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_12),
.A2(n_38),
.B1(n_39),
.B2(n_45),
.Y(n_49)
);

NAND2xp33_ASAP7_75t_SL g150 ( 
.A(n_12),
.B(n_43),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_13),
.A2(n_34),
.B1(n_59),
.B2(n_60),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_14),
.A2(n_38),
.B1(n_39),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_14),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_14),
.A2(n_42),
.B1(n_43),
.B2(n_102),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_14),
.A2(n_59),
.B1(n_60),
.B2(n_102),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_102),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_15),
.A2(n_59),
.B1(n_60),
.B2(n_68),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_15),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_68),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_15),
.A2(n_42),
.B1(n_43),
.B2(n_68),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_16),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_16),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_16),
.A2(n_40),
.B1(n_59),
.B2(n_60),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_16),
.A2(n_28),
.B1(n_29),
.B2(n_40),
.Y(n_164)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_123),
.B1(n_293),
.B2(n_294),
.Y(n_18)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_19),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_121),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_105),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_21),
.B(n_105),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_71),
.C(n_87),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_22),
.A2(n_23),
.B1(n_71),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_54),
.B2(n_70),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_35),
.B1(n_36),
.B2(n_53),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_26),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_26),
.A2(n_36),
.B(n_70),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_26),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_31),
.B(n_32),
.Y(n_26)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_27),
.A2(n_31),
.B1(n_92),
.B2(n_155),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_27),
.B(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_27),
.A2(n_31),
.B1(n_237),
.B2(n_239),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_28),
.A2(n_29),
.B1(n_63),
.B2(n_64),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_28),
.B(n_249),
.Y(n_248)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_31),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_31),
.B(n_211),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_33),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_90)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B(n_46),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_37),
.A2(n_41),
.B1(n_48),
.B2(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_39),
.A2(n_48),
.B(n_133),
.C(n_134),
.Y(n_132)
);

AOI32xp33_ASAP7_75t_L g149 ( 
.A1(n_39),
.A2(n_42),
.A3(n_45),
.B1(n_135),
.B2(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_41),
.B(n_51),
.Y(n_104)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_41),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_41),
.A2(n_46),
.B(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_41),
.A2(n_48),
.B1(n_101),
.B2(n_179),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_42),
.A2(n_43),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_48),
.A2(n_101),
.B(n_103),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_61),
.B1(n_66),
.B2(n_69),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_57),
.A2(n_61),
.B1(n_69),
.B2(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_59),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

AO22x1_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_60),
.B1(n_79),
.B2(n_80),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_59),
.B(n_223),
.Y(n_222)
);

OAI21xp33_ASAP7_75t_L g208 ( 
.A1(n_60),
.A2(n_79),
.B(n_133),
.Y(n_208)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_61),
.A2(n_69),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_61),
.B(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_61),
.A2(n_69),
.B1(n_97),
.B2(n_143),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_61),
.A2(n_69),
.B1(n_203),
.B2(n_261),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_65),
.A2(n_67),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_65),
.A2(n_142),
.B(n_144),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_65),
.A2(n_144),
.B(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_65),
.B(n_133),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_69),
.B(n_145),
.Y(n_204)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_71),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_75),
.B(n_86),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_75),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_73),
.A2(n_202),
.B(n_204),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_73),
.A2(n_204),
.B(n_221),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_74),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_76),
.A2(n_82),
.B1(n_84),
.B2(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_76),
.A2(n_84),
.B1(n_138),
.B2(n_140),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_76),
.A2(n_140),
.B(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_76),
.A2(n_177),
.B(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_77),
.A2(n_81),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_77),
.B(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_81),
.B(n_159),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_84),
.A2(n_138),
.B(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_84),
.A2(n_99),
.B(n_158),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

FAx1_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_106),
.CI(n_107),
.CON(n_105),
.SN(n_105)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_87),
.B(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_98),
.C(n_100),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_88),
.A2(n_89),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_95),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_90),
.A2(n_95),
.B1(n_96),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_90),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_93),
.A2(n_94),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_93),
.A2(n_94),
.B1(n_153),
.B2(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_93),
.A2(n_232),
.B(n_233),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_94),
.A2(n_164),
.B(n_210),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_94),
.A2(n_210),
.B(n_238),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_94),
.B(n_133),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_98),
.B(n_100),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_104),
.B(n_132),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g295 ( 
.A(n_105),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.Y(n_107)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_113),
.B1(n_114),
.B2(n_116),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_109),
.Y(n_116)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_123),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_287),
.B(n_292),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_275),
.B(n_286),
.Y(n_125)
);

OAI321xp33_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_182),
.A3(n_194),
.B1(n_273),
.B2(n_274),
.C(n_297),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_165),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_128),
.B(n_165),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_147),
.C(n_156),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_129),
.B(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_136),
.B2(n_146),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_137),
.C(n_141),
.Y(n_171)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_141),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_147),
.B(n_156),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_152),
.Y(n_181)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.C(n_163),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_157),
.B(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_160),
.A2(n_161),
.B1(n_163),
.B2(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_163),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_172),
.B2(n_173),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_171),
.C(n_172),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_170),
.Y(n_192)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_181),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_180),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_180),
.C(n_181),
.Y(n_193)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_178),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_183),
.B(n_184),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_193),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_186),
.B(n_188),
.C(n_193),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_190),
.B(n_191),
.C(n_192),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_214),
.B(n_272),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_212),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_196),
.B(n_212),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_201),
.C(n_205),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_197),
.A2(n_198),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_201),
.A2(n_205),
.B1(n_206),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_201),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_207),
.B(n_209),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_265),
.B(n_271),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_253),
.B(n_264),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_234),
.B(n_252),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_224),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_218),
.B(n_224),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_222),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_219),
.A2(n_220),
.B1(n_222),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_222),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_231),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_229),
.C(n_231),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_230),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_232),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_242),
.B(n_251),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_240),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_236),
.B(n_240),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_246),
.B(n_250),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_244),
.B(n_245),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_254),
.B(n_255),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_260),
.C(n_263),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_257)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_258),
.Y(n_263)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_260),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_266),
.B(n_267),
.Y(n_271)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_285),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_285),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_280),
.C(n_281),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_289),
.Y(n_292)
);


endmodule