module real_jpeg_6200_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_11;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_9;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g91 ( 
.A(n_0),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_4),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_4),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_5),
.B(n_20),
.Y(n_19)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_5),
.B(n_58),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_5),
.A2(n_29),
.B1(n_98),
.B2(n_100),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_5),
.B(n_112),
.C(n_113),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_6),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_7),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_7),
.A2(n_38),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_68),
.Y(n_8)
);

AOI21xp5_ASAP7_75t_L g9 ( 
.A1(n_10),
.A2(n_43),
.B(n_67),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_23),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_19),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_14),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B(n_30),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_25),
.B(n_33),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_25),
.A2(n_71),
.B1(n_72),
.B2(n_81),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_36),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_57),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_57),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_53),
.B(n_56),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_58),
.B(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_117),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_82),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_70),
.B(n_82),
.Y(n_118)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_108),
.B1(n_115),
.B2(n_116),
.Y(n_82)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_97),
.B(n_103),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_92),
.B1(n_94),
.B2(n_96),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);


endmodule