module real_jpeg_5328_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_1),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_2),
.A2(n_126),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_2),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_2),
.A2(n_140),
.B1(n_173),
.B2(n_176),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_2),
.A2(n_140),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_2),
.A2(n_30),
.B1(n_140),
.B2(n_300),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_3),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_3),
.A2(n_40),
.B1(n_73),
.B2(n_75),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_3),
.A2(n_40),
.B1(n_114),
.B2(n_117),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_3),
.A2(n_40),
.B1(n_175),
.B2(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_4),
.A2(n_21),
.B1(n_22),
.B2(n_26),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_4),
.A2(n_21),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_5),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_6),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_6),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g315 ( 
.A(n_6),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_7),
.Y(n_123)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_7),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_7),
.Y(n_166)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_8),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_9),
.Y(n_116)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_9),
.Y(n_117)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_9),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_9),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_9),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_10),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_10),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_10),
.A2(n_51),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_10),
.A2(n_51),
.B1(n_184),
.B2(n_187),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_10),
.B(n_127),
.Y(n_236)
);

O2A1O1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_10),
.A2(n_82),
.B(n_260),
.C(n_267),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_10),
.B(n_290),
.C(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_10),
.B(n_80),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_10),
.B(n_37),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_10),
.B(n_63),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g290 ( 
.A(n_11),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_227),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_225),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_199),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_16),
.B(n_199),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_143),
.C(n_178),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_17),
.B(n_178),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_78),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_18),
.B(n_111),
.C(n_141),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_44),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_19),
.B(n_44),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_28),
.B(n_35),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_20),
.A2(n_149),
.B(n_152),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_29),
.B(n_38),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_29),
.A2(n_183),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_29),
.B(n_183),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_29),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_31),
.Y(n_187)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_31),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_32),
.Y(n_292)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_35),
.B(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_35),
.B(n_298),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_71),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_45),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_53),
.Y(n_45)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_46),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_49),
.Y(n_193)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_49),
.Y(n_266)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_50),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_50),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_51),
.B(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_51),
.A2(n_120),
.B(n_159),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_L g260 ( 
.A1(n_51),
.A2(n_261),
.B(n_264),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_53),
.B(n_72),
.Y(n_198)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_53),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_53),
.B(n_275),
.Y(n_274)
);

NOR2x1_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_63),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_57),
.B1(n_59),
.B2(n_62),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AO22x2_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_64),
.B1(n_66),
.B2(n_69),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_63),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_63),
.B(n_275),
.Y(n_294)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_71),
.A2(n_191),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_71),
.B(n_274),
.Y(n_303)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_77),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_111),
.B1(n_141),
.B2(n_142),
.Y(n_78)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_91),
.B(n_105),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_80),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_80),
.B(n_172),
.Y(n_249)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_81),
.B(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_84),
.Y(n_276)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_91),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_91),
.B(n_105),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_92),
.B(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_96),
.B1(n_99),
.B2(n_101),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_95),
.Y(n_263)
);

AOI32xp33_ASAP7_75t_L g153 ( 
.A1(n_96),
.A2(n_154),
.A3(n_155),
.B1(n_158),
.B2(n_161),
.Y(n_153)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_98),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_104),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_104),
.Y(n_269)
);

INVxp67_ASAP7_75t_SL g170 ( 
.A(n_105),
.Y(n_170)
);

INVx6_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_137),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_118),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_127),
.Y(n_145)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_138),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_118),
.B(n_207),
.Y(n_243)
);

NOR2x1_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_127),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_122),
.B1(n_124),
.B2(n_126),
.Y(n_119)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_127),
.B(n_207),
.Y(n_206)
);

AO22x2_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_130),
.B1(n_133),
.B2(n_135),
.Y(n_127)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_137),
.B(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_143),
.B(n_359),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.C(n_167),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_144),
.B(n_167),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_146),
.B(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_147),
.B(n_356),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_153),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_148),
.B(n_153),
.Y(n_240)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp33_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_171),
.B(n_209),
.Y(n_234)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_189),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_189),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_188),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_180),
.B(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_186),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_188),
.B(n_312),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B(n_198),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_190),
.A2(n_222),
.B(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_190),
.B(n_252),
.Y(n_273)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_198),
.B(n_294),
.Y(n_336)
);

BUFx24_ASAP7_75t_SL g364 ( 
.A(n_199),
.Y(n_364)
);

FAx1_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_216),
.CI(n_224),
.CON(n_199),
.SN(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_215),
.Y(n_208)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_210),
.Y(n_248)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_215),
.B(n_249),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_220),
.B1(n_221),
.B2(n_223),
.Y(n_216)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_217),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_217),
.A2(n_223),
.B1(n_259),
.B2(n_339),
.Y(n_338)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_348),
.B(n_361),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_280),
.B(n_347),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_254),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_230),
.B(n_254),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_241),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_239),
.B2(n_240),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_233),
.B(n_239),
.C(n_241),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.C(n_237),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_256),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_235),
.A2(n_236),
.B1(n_237),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_238),
.B(n_313),
.Y(n_324)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_242),
.B(n_245),
.C(n_251),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_250),
.B1(n_251),
.B2(n_253),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_245),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_249),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.C(n_270),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_255),
.B(n_343),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_258),
.A2(n_270),
.B1(n_271),
.B2(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_258),
.Y(n_344)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_259),
.Y(n_339)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx8_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_SL g264 ( 
.A(n_265),
.Y(n_264)
);

INVx8_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_341),
.B(n_346),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_331),
.B(n_340),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_307),
.B(n_330),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_295),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_284),
.B(n_295),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_293),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_285),
.A2(n_286),
.B1(n_293),
.B2(n_310),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_293),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_302),
.Y(n_295)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_296),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_302)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_303),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_304),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_304),
.B(n_305),
.C(n_333),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_308),
.A2(n_316),
.B(n_329),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_311),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_311),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_325),
.B(n_328),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_324),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_323),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx6_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_326),
.B(n_327),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_334),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_334),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_338),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_336),
.B(n_337),
.C(n_338),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_345),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_342),
.B(n_345),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_357),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_350),
.B(n_351),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_355),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_353),
.B(n_354),
.C(n_355),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_357),
.A2(n_362),
.B(n_363),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_360),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_358),
.B(n_360),
.Y(n_363)
);


endmodule