module fake_netlist_6_4693_n_942 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_942);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_942;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_209;
wire n_680;
wire n_760;
wire n_741;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_718;
wire n_517;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_491;
wire n_878;
wire n_772;
wire n_656;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_844;
wire n_343;
wire n_886;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_859;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_24),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_115),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_138),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_1),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_63),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_29),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_68),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_3),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_142),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_108),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_14),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_24),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_184),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_180),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_27),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_134),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_86),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_99),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_2),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_0),
.Y(n_212)
);

BUFx10_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_55),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_164),
.Y(n_215)
);

HB1xp67_ASAP7_75t_SL g216 ( 
.A(n_53),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_74),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_174),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_132),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_8),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_147),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_27),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_179),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_83),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_42),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_118),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_157),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_183),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_41),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_69),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_173),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_100),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_19),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_67),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_14),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_103),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_106),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_95),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_22),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_188),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_6),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_165),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_78),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_49),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_105),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_88),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_168),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_178),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_111),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_171),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_1),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_112),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_65),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_130),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_123),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_125),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_23),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_29),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_82),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_0),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_154),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_47),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_159),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_52),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_135),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_116),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_60),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_31),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_62),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_3),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_36),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_110),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_2),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_113),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_144),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_21),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_175),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_177),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_71),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_186),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_153),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_126),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_151),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_39),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_30),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_8),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_70),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_185),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_221),
.B(n_4),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_268),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_268),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_190),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_268),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_194),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_268),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_198),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_201),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_202),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_201),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_206),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_212),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_251),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_220),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_251),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_196),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_211),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_222),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_233),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_225),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_239),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_257),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_235),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_241),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_271),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_258),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_197),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_273),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_285),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_270),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_276),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_191),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_218),
.B(n_4),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_242),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_191),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_283),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_283),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_197),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_242),
.B(n_5),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_193),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_204),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_208),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_210),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_284),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_217),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_211),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_217),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_224),
.Y(n_337)
);

INVxp33_ASAP7_75t_L g338 ( 
.A(n_216),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_229),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_226),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_244),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_244),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_227),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_230),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_263),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_232),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_234),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_204),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_263),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_238),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_229),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_267),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_267),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_195),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_240),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_354),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_336),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_292),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_290),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_R g360 ( 
.A(n_292),
.B(n_192),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_336),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_342),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_291),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_316),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_293),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_321),
.B(n_246),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_295),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_338),
.B(n_294),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_329),
.Y(n_369)
);

INVx5_ASAP7_75t_L g370 ( 
.A(n_299),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_342),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_323),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_349),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_324),
.Y(n_374)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_299),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_310),
.B(n_274),
.Y(n_376)
);

AND2x6_ASAP7_75t_L g377 ( 
.A(n_323),
.B(n_250),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_348),
.B(n_298),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_327),
.B(n_260),
.Y(n_379)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_317),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_298),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_349),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_325),
.B(n_248),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_334),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_352),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_341),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_317),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_331),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_352),
.Y(n_389)
);

OAI21x1_ASAP7_75t_L g390 ( 
.A1(n_289),
.A2(n_277),
.B(n_259),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_353),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_353),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_326),
.B(n_282),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_332),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_300),
.Y(n_395)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_300),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_301),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_301),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_343),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_344),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_303),
.A2(n_200),
.B1(n_260),
.B2(n_286),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_346),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_330),
.B(n_204),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_297),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_319),
.B(n_207),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_R g406 ( 
.A(n_303),
.B(n_307),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_347),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_297),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_350),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_345),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_306),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_330),
.B(n_199),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_307),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_393),
.B(n_312),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_374),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_369),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_368),
.B(n_309),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_375),
.B(n_355),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_388),
.Y(n_419)
);

AND3x2_ASAP7_75t_L g420 ( 
.A(n_381),
.B(n_322),
.C(n_296),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_375),
.B(n_337),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_375),
.B(n_337),
.Y(n_422)
);

INVx5_ASAP7_75t_L g423 ( 
.A(n_377),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_404),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_363),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_365),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_412),
.B(n_309),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_387),
.Y(n_428)
);

INVx5_ASAP7_75t_L g429 ( 
.A(n_377),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_404),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_387),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_393),
.B(n_340),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_401),
.B(n_335),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_356),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_394),
.Y(n_435)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_377),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_393),
.B(n_374),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_404),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_404),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_376),
.B(n_340),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_399),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_360),
.B(n_311),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_408),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_380),
.B(n_311),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_387),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_378),
.B(n_315),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_400),
.Y(n_447)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_377),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_387),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_408),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_402),
.B(n_313),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_407),
.B(n_302),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_405),
.B(n_315),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_380),
.B(n_333),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_396),
.B(n_286),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_408),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_403),
.B(n_406),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_409),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_408),
.Y(n_459)
);

BUFx6f_ASAP7_75t_SL g460 ( 
.A(n_396),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_390),
.A2(n_328),
.B1(n_383),
.B2(n_366),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_380),
.Y(n_462)
);

OR2x2_ASAP7_75t_L g463 ( 
.A(n_358),
.B(n_339),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_359),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_396),
.B(n_333),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_413),
.B(n_296),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_359),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_411),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_367),
.Y(n_469)
);

NOR2x1p5_ASAP7_75t_L g470 ( 
.A(n_395),
.B(n_318),
.Y(n_470)
);

NOR2x1p5_ASAP7_75t_L g471 ( 
.A(n_397),
.B(n_413),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_398),
.A2(n_320),
.B1(n_255),
.B2(n_254),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_367),
.B(n_351),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_371),
.B(n_207),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_373),
.B(n_305),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_382),
.B(n_207),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_372),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_372),
.B(n_302),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_370),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_389),
.B(n_213),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_370),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_370),
.Y(n_482)
);

OR2x6_ASAP7_75t_L g483 ( 
.A(n_390),
.B(n_314),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_444),
.B(n_391),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_462),
.B(n_427),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_433),
.B(n_379),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_440),
.B(n_203),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_469),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_440),
.B(n_308),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_461),
.B(n_458),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_458),
.B(n_205),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_469),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_465),
.B(n_392),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_416),
.B(n_209),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_419),
.B(n_214),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_415),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_446),
.B(n_357),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_483),
.A2(n_454),
.B1(n_453),
.B2(n_457),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_477),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_475),
.B(n_417),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_477),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_415),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_455),
.A2(n_269),
.B1(n_215),
.B2(n_219),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_478),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_435),
.B(n_223),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_434),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_437),
.B(n_308),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_441),
.B(n_228),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_476),
.B(n_357),
.Y(n_509)
);

AO22x1_ASAP7_75t_L g510 ( 
.A1(n_414),
.A2(n_250),
.B1(n_377),
.B2(n_362),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_478),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_475),
.B(n_361),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_473),
.B(n_361),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_447),
.B(n_231),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_437),
.B(n_236),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_432),
.A2(n_377),
.B(n_243),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_464),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_467),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_431),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_483),
.A2(n_275),
.B1(n_237),
.B2(n_245),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_418),
.B(n_247),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_424),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_414),
.B(n_362),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_483),
.A2(n_279),
.B1(n_249),
.B2(n_266),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_421),
.A2(n_422),
.B(n_428),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_483),
.A2(n_250),
.B1(n_213),
.B2(n_288),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_425),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_414),
.B(n_425),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_451),
.A2(n_280),
.B1(n_252),
.B2(n_253),
.Y(n_529)
);

NOR3xp33_ASAP7_75t_L g530 ( 
.A(n_466),
.B(n_468),
.C(n_463),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_468),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_426),
.B(n_256),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_428),
.A2(n_370),
.B(n_250),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_452),
.B(n_304),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_426),
.B(n_261),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_472),
.B(n_385),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_442),
.B(n_385),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_470),
.Y(n_538)
);

BUFx6f_ASAP7_75t_SL g539 ( 
.A(n_451),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_424),
.Y(n_540)
);

OAI221xp5_ASAP7_75t_L g541 ( 
.A1(n_452),
.A2(n_304),
.B1(n_262),
.B2(n_264),
.C(n_265),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_449),
.B(n_272),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_430),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_430),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_431),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_449),
.B(n_278),
.Y(n_546)
);

NAND2xp33_ASAP7_75t_L g547 ( 
.A(n_423),
.B(n_281),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_438),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_445),
.B(n_287),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_451),
.A2(n_213),
.B1(n_288),
.B2(n_411),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_438),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_445),
.B(n_370),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_445),
.B(n_288),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_439),
.B(n_43),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_522),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_531),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_485),
.B(n_439),
.Y(n_557)
);

BUFx4f_ASAP7_75t_SL g558 ( 
.A(n_523),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_499),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_496),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_511),
.B(n_443),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_501),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_501),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_488),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_511),
.B(n_443),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_499),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_496),
.B(n_502),
.Y(n_567)
);

BUFx8_ASAP7_75t_SL g568 ( 
.A(n_506),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_506),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_527),
.B(n_450),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_513),
.B(n_463),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_527),
.B(n_450),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_R g573 ( 
.A(n_538),
.B(n_434),
.Y(n_573)
);

AND3x1_ASAP7_75t_SL g574 ( 
.A(n_541),
.B(n_471),
.C(n_433),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_504),
.B(n_456),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_522),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_488),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_502),
.B(n_456),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_492),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_L g580 ( 
.A1(n_490),
.A2(n_448),
.B(n_436),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_539),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_540),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_504),
.B(n_431),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_545),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_492),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_545),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_540),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_544),
.Y(n_588)
);

INVx6_ASAP7_75t_L g589 ( 
.A(n_545),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_525),
.A2(n_448),
.B(n_436),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_484),
.B(n_356),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_543),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_544),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_507),
.B(n_420),
.Y(n_594)
);

NAND3xp33_ASAP7_75t_SL g595 ( 
.A(n_503),
.B(n_384),
.C(n_364),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_518),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_548),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_507),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_500),
.B(n_474),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_548),
.Y(n_600)
);

NOR3xp33_ASAP7_75t_SL g601 ( 
.A(n_512),
.B(n_480),
.C(n_384),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_498),
.B(n_436),
.Y(n_602)
);

NAND2xp33_ASAP7_75t_SL g603 ( 
.A(n_539),
.B(n_460),
.Y(n_603)
);

AND3x1_ASAP7_75t_SL g604 ( 
.A(n_530),
.B(n_386),
.C(n_364),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_518),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_489),
.B(n_448),
.Y(n_606)
);

AND2x6_ASAP7_75t_L g607 ( 
.A(n_489),
.B(n_431),
.Y(n_607)
);

BUFx12f_ASAP7_75t_SL g608 ( 
.A(n_534),
.Y(n_608)
);

NOR3xp33_ASAP7_75t_SL g609 ( 
.A(n_536),
.B(n_410),
.C(n_386),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_543),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_517),
.Y(n_611)
);

BUFx10_ASAP7_75t_L g612 ( 
.A(n_537),
.Y(n_612)
);

OAI21xp5_ASAP7_75t_L g613 ( 
.A1(n_602),
.A2(n_528),
.B(n_516),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_566),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_590),
.A2(n_545),
.B(n_519),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_599),
.A2(n_497),
.B1(n_493),
.B2(n_520),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_598),
.B(n_534),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_566),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_568),
.Y(n_619)
);

AO31x2_ASAP7_75t_L g620 ( 
.A1(n_557),
.A2(n_551),
.A3(n_554),
.B(n_517),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_580),
.A2(n_545),
.B(n_547),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_606),
.A2(n_547),
.B(n_515),
.Y(n_622)
);

OAI21x1_ASAP7_75t_L g623 ( 
.A1(n_570),
.A2(n_551),
.B(n_552),
.Y(n_623)
);

CKINVDCx11_ASAP7_75t_R g624 ( 
.A(n_569),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_596),
.B(n_487),
.Y(n_625)
);

OAI21x1_ASAP7_75t_L g626 ( 
.A1(n_572),
.A2(n_549),
.B(n_546),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_608),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g628 ( 
.A1(n_561),
.A2(n_521),
.B(n_491),
.Y(n_628)
);

INVxp67_ASAP7_75t_SL g629 ( 
.A(n_584),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_605),
.B(n_532),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_591),
.B(n_535),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_583),
.A2(n_542),
.B(n_429),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_565),
.A2(n_586),
.B(n_584),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_584),
.A2(n_429),
.B(n_423),
.Y(n_634)
);

OAI22x1_ASAP7_75t_L g635 ( 
.A1(n_571),
.A2(n_509),
.B1(n_503),
.B2(n_486),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_559),
.B(n_529),
.Y(n_636)
);

OAI21xp5_ASAP7_75t_L g637 ( 
.A1(n_575),
.A2(n_529),
.B(n_495),
.Y(n_637)
);

AO21x1_ASAP7_75t_L g638 ( 
.A1(n_563),
.A2(n_524),
.B(n_553),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_563),
.B(n_494),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_584),
.A2(n_429),
.B(n_423),
.Y(n_640)
);

OAI21x1_ASAP7_75t_L g641 ( 
.A1(n_555),
.A2(n_533),
.B(n_508),
.Y(n_641)
);

OAI21x1_ASAP7_75t_L g642 ( 
.A1(n_555),
.A2(n_582),
.B(n_576),
.Y(n_642)
);

AO31x2_ASAP7_75t_L g643 ( 
.A1(n_592),
.A2(n_610),
.A3(n_564),
.B(n_585),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_L g644 ( 
.A1(n_562),
.A2(n_514),
.B(n_505),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_584),
.A2(n_429),
.B(n_423),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_556),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_SL g647 ( 
.A1(n_586),
.A2(n_539),
.B(n_460),
.Y(n_647)
);

OAI21xp33_ASAP7_75t_L g648 ( 
.A1(n_573),
.A2(n_550),
.B(n_486),
.Y(n_648)
);

OAI21x1_ASAP7_75t_L g649 ( 
.A1(n_555),
.A2(n_526),
.B(n_482),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_562),
.B(n_538),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_567),
.B(n_410),
.Y(n_651)
);

OAI21x1_ASAP7_75t_SL g652 ( 
.A1(n_585),
.A2(n_482),
.B(n_481),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_564),
.A2(n_460),
.B1(n_431),
.B2(n_459),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_589),
.Y(n_654)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_608),
.Y(n_655)
);

A2O1A1Ixp33_ASAP7_75t_L g656 ( 
.A1(n_611),
.A2(n_479),
.B(n_510),
.C(n_459),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_586),
.A2(n_429),
.B(n_423),
.Y(n_657)
);

OAI21x1_ASAP7_75t_L g658 ( 
.A1(n_576),
.A2(n_510),
.B(n_459),
.Y(n_658)
);

NOR3xp33_ASAP7_75t_L g659 ( 
.A(n_595),
.B(n_5),
.C(n_6),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_594),
.B(n_7),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_592),
.A2(n_459),
.B1(n_91),
.B2(n_92),
.Y(n_661)
);

OAI21x1_ASAP7_75t_L g662 ( 
.A1(n_576),
.A2(n_459),
.B(n_90),
.Y(n_662)
);

OAI21x1_ASAP7_75t_L g663 ( 
.A1(n_662),
.A2(n_610),
.B(n_593),
.Y(n_663)
);

AOI21x1_ASAP7_75t_L g664 ( 
.A1(n_621),
.A2(n_579),
.B(n_577),
.Y(n_664)
);

AO21x2_ASAP7_75t_L g665 ( 
.A1(n_613),
.A2(n_588),
.B(n_587),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_646),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_654),
.Y(n_667)
);

NOR2x1_ASAP7_75t_SL g668 ( 
.A(n_653),
.B(n_586),
.Y(n_668)
);

AO21x2_ASAP7_75t_L g669 ( 
.A1(n_638),
.A2(n_588),
.B(n_587),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_631),
.B(n_612),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_643),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_615),
.A2(n_586),
.B(n_603),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_643),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_643),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_659),
.A2(n_635),
.B1(n_594),
.B2(n_616),
.Y(n_675)
);

A2O1A1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_637),
.A2(n_601),
.B(n_609),
.C(n_594),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_624),
.Y(n_677)
);

BUFx12f_ASAP7_75t_L g678 ( 
.A(n_624),
.Y(n_678)
);

OA21x2_ASAP7_75t_L g679 ( 
.A1(n_623),
.A2(n_600),
.B(n_597),
.Y(n_679)
);

O2A1O1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_659),
.A2(n_556),
.B(n_560),
.C(n_567),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_648),
.A2(n_558),
.B1(n_612),
.B2(n_567),
.Y(n_681)
);

OAI21x1_ASAP7_75t_L g682 ( 
.A1(n_642),
.A2(n_593),
.B(n_582),
.Y(n_682)
);

OAI21x1_ASAP7_75t_L g683 ( 
.A1(n_658),
.A2(n_593),
.B(n_582),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_617),
.B(n_612),
.Y(n_684)
);

AOI221xp5_ASAP7_75t_L g685 ( 
.A1(n_625),
.A2(n_569),
.B1(n_581),
.B2(n_603),
.C(n_560),
.Y(n_685)
);

AO31x2_ASAP7_75t_L g686 ( 
.A1(n_656),
.A2(n_600),
.A3(n_597),
.B(n_574),
.Y(n_686)
);

NAND3xp33_ASAP7_75t_L g687 ( 
.A(n_636),
.B(n_630),
.C(n_639),
.Y(n_687)
);

OA21x2_ASAP7_75t_L g688 ( 
.A1(n_656),
.A2(n_578),
.B(n_607),
.Y(n_688)
);

NAND3xp33_ASAP7_75t_L g689 ( 
.A(n_644),
.B(n_581),
.C(n_578),
.Y(n_689)
);

OAI21x1_ASAP7_75t_L g690 ( 
.A1(n_641),
.A2(n_607),
.B(n_589),
.Y(n_690)
);

OR2x2_ASAP7_75t_L g691 ( 
.A(n_643),
.B(n_614),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_L g692 ( 
.A1(n_650),
.A2(n_629),
.B1(n_618),
.B2(n_646),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_660),
.B(n_578),
.Y(n_693)
);

OAI21x1_ASAP7_75t_L g694 ( 
.A1(n_633),
.A2(n_622),
.B(n_626),
.Y(n_694)
);

NOR2xp67_ASAP7_75t_L g695 ( 
.A(n_654),
.B(n_44),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_SL g696 ( 
.A(n_619),
.B(n_568),
.Y(n_696)
);

OA21x2_ASAP7_75t_L g697 ( 
.A1(n_628),
.A2(n_607),
.B(n_604),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_629),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_651),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_649),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_627),
.B(n_607),
.Y(n_701)
);

O2A1O1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_661),
.A2(n_607),
.B(n_9),
.C(n_10),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_620),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_652),
.Y(n_704)
);

A2O1A1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_632),
.A2(n_607),
.B(n_589),
.C(n_10),
.Y(n_705)
);

NOR3xp33_ASAP7_75t_L g706 ( 
.A(n_651),
.B(n_7),
.C(n_9),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_647),
.A2(n_589),
.B(n_96),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_706),
.A2(n_627),
.B1(n_655),
.B2(n_619),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_666),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_675),
.A2(n_655),
.B1(n_12),
.B2(n_13),
.Y(n_710)
);

AOI21xp33_ASAP7_75t_L g711 ( 
.A1(n_680),
.A2(n_620),
.B(n_12),
.Y(n_711)
);

HB1xp67_ASAP7_75t_L g712 ( 
.A(n_666),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_671),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_667),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_670),
.A2(n_657),
.B1(n_645),
.B2(n_640),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_699),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_701),
.B(n_693),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_699),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_698),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_677),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_701),
.B(n_620),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_693),
.B(n_620),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_672),
.A2(n_634),
.B(n_97),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_698),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_687),
.A2(n_11),
.B1(n_13),
.B2(n_15),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_667),
.B(n_45),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_681),
.A2(n_11),
.B1(n_15),
.B2(n_16),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_687),
.B(n_16),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_R g729 ( 
.A(n_696),
.B(n_189),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_684),
.B(n_17),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_667),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_667),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_689),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_676),
.B(n_18),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_667),
.Y(n_735)
);

AND2x6_ASAP7_75t_L g736 ( 
.A(n_671),
.B(n_46),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_695),
.B(n_48),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_674),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_685),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_692),
.B(n_20),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_695),
.B(n_50),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_689),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_742)
);

AOI21xp33_ASAP7_75t_L g743 ( 
.A1(n_702),
.A2(n_23),
.B(n_25),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_697),
.A2(n_678),
.B1(n_691),
.B2(n_704),
.Y(n_744)
);

OAI22xp33_ASAP7_75t_L g745 ( 
.A1(n_678),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_SL g746 ( 
.A1(n_697),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_697),
.B(n_31),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_674),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_691),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_SL g750 ( 
.A1(n_697),
.A2(n_668),
.B1(n_707),
.B2(n_688),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_SL g751 ( 
.A1(n_668),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_673),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_SL g753 ( 
.A1(n_688),
.A2(n_704),
.B1(n_700),
.B2(n_673),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_686),
.B(n_32),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_686),
.Y(n_755)
);

OR2x6_ASAP7_75t_L g756 ( 
.A(n_705),
.B(n_51),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_686),
.B(n_33),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_739),
.A2(n_700),
.B1(n_688),
.B2(n_703),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_710),
.A2(n_700),
.B1(n_688),
.B2(n_703),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_721),
.B(n_703),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_720),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_710),
.A2(n_669),
.B1(n_665),
.B2(n_663),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_721),
.B(n_686),
.Y(n_763)
);

OAI221xp5_ASAP7_75t_L g764 ( 
.A1(n_708),
.A2(n_733),
.B1(n_725),
.B2(n_743),
.C(n_751),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_749),
.B(n_669),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_712),
.Y(n_766)
);

OAI211xp5_ASAP7_75t_SL g767 ( 
.A1(n_708),
.A2(n_686),
.B(n_35),
.C(n_36),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_734),
.A2(n_669),
.B1(n_665),
.B2(n_663),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_733),
.A2(n_665),
.B1(n_694),
.B2(n_690),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_725),
.A2(n_694),
.B1(n_690),
.B2(n_679),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_730),
.A2(n_664),
.B1(n_679),
.B2(n_37),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_709),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_724),
.B(n_679),
.Y(n_773)
);

HB1xp67_ASAP7_75t_L g774 ( 
.A(n_709),
.Y(n_774)
);

AOI221xp5_ASAP7_75t_L g775 ( 
.A1(n_745),
.A2(n_742),
.B1(n_727),
.B2(n_730),
.C(n_711),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_756),
.A2(n_679),
.B1(n_682),
.B2(n_683),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_756),
.A2(n_682),
.B1(n_683),
.B2(n_664),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_719),
.B(n_34),
.Y(n_778)
);

AOI222xp33_ASAP7_75t_L g779 ( 
.A1(n_728),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.C1(n_39),
.C2(n_40),
.Y(n_779)
);

AOI21x1_ASAP7_75t_L g780 ( 
.A1(n_723),
.A2(n_728),
.B(n_715),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_756),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_717),
.A2(n_42),
.B1(n_54),
.B2(n_56),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_717),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_783)
);

AOI211xp5_ASAP7_75t_L g784 ( 
.A1(n_747),
.A2(n_61),
.B(n_64),
.C(n_66),
.Y(n_784)
);

OAI221xp5_ASAP7_75t_L g785 ( 
.A1(n_746),
.A2(n_72),
.B1(n_73),
.B2(n_75),
.C(n_76),
.Y(n_785)
);

AO21x2_ASAP7_75t_L g786 ( 
.A1(n_747),
.A2(n_77),
.B(n_79),
.Y(n_786)
);

OAI221xp5_ASAP7_75t_L g787 ( 
.A1(n_740),
.A2(n_80),
.B1(n_81),
.B2(n_84),
.C(n_85),
.Y(n_787)
);

OAI22xp33_ASAP7_75t_L g788 ( 
.A1(n_716),
.A2(n_87),
.B1(n_89),
.B2(n_93),
.Y(n_788)
);

OA21x2_ASAP7_75t_L g789 ( 
.A1(n_744),
.A2(n_755),
.B(n_752),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_713),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_721),
.B(n_94),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_713),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_SL g793 ( 
.A1(n_729),
.A2(n_98),
.B1(n_101),
.B2(n_102),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_738),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_790),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_766),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_790),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_792),
.B(n_754),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_792),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_763),
.B(n_744),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_763),
.B(n_753),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_794),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_764),
.A2(n_722),
.B1(n_717),
.B2(n_736),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_794),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_794),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_773),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_773),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_772),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_760),
.B(n_722),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_760),
.B(n_722),
.Y(n_810)
);

BUFx12f_ASAP7_75t_L g811 ( 
.A(n_761),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_789),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_774),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_789),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_789),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_789),
.Y(n_816)
);

INVxp67_ASAP7_75t_L g817 ( 
.A(n_765),
.Y(n_817)
);

OAI211xp5_ASAP7_75t_L g818 ( 
.A1(n_779),
.A2(n_729),
.B(n_757),
.C(n_750),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_765),
.B(n_748),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_758),
.B(n_748),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_768),
.B(n_738),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_772),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_769),
.B(n_732),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_818),
.A2(n_781),
.B1(n_784),
.B2(n_785),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_796),
.B(n_772),
.Y(n_825)
);

NAND2xp33_ASAP7_75t_R g826 ( 
.A(n_798),
.B(n_791),
.Y(n_826)
);

OAI221xp5_ASAP7_75t_L g827 ( 
.A1(n_818),
.A2(n_775),
.B1(n_784),
.B2(n_779),
.C(n_793),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_813),
.B(n_786),
.Y(n_828)
);

AOI221xp5_ASAP7_75t_L g829 ( 
.A1(n_798),
.A2(n_771),
.B1(n_785),
.B2(n_767),
.C(n_778),
.Y(n_829)
);

NAND4xp25_ASAP7_75t_L g830 ( 
.A(n_803),
.B(n_778),
.C(n_771),
.D(n_759),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_809),
.B(n_791),
.Y(n_831)
);

AOI221xp5_ASAP7_75t_L g832 ( 
.A1(n_806),
.A2(n_787),
.B1(n_786),
.B2(n_788),
.C(n_782),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_795),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_817),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_795),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_806),
.B(n_786),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_807),
.B(n_770),
.Y(n_837)
);

AOI222xp33_ASAP7_75t_L g838 ( 
.A1(n_800),
.A2(n_736),
.B1(n_762),
.B2(n_783),
.C1(n_791),
.C2(n_741),
.Y(n_838)
);

INVxp67_ASAP7_75t_L g839 ( 
.A(n_807),
.Y(n_839)
);

OAI221xp5_ASAP7_75t_L g840 ( 
.A1(n_817),
.A2(n_718),
.B1(n_780),
.B2(n_808),
.C(n_823),
.Y(n_840)
);

NAND3xp33_ASAP7_75t_L g841 ( 
.A(n_823),
.B(n_777),
.C(n_776),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_834),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_834),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_839),
.B(n_801),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_833),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_839),
.B(n_801),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_835),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_836),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_825),
.B(n_801),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_837),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_831),
.B(n_800),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_827),
.B(n_811),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_828),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_850),
.B(n_800),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_845),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_850),
.B(n_841),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_845),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_847),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_847),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_854),
.B(n_844),
.Y(n_860)
);

NAND2xp33_ASAP7_75t_R g861 ( 
.A(n_856),
.B(n_852),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_854),
.B(n_844),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_855),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_857),
.B(n_849),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_860),
.B(n_846),
.Y(n_865)
);

AOI222xp33_ASAP7_75t_L g866 ( 
.A1(n_860),
.A2(n_824),
.B1(n_829),
.B2(n_832),
.C1(n_846),
.C2(n_840),
.Y(n_866)
);

NAND2xp33_ASAP7_75t_SL g867 ( 
.A(n_861),
.B(n_826),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_862),
.B(n_849),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_862),
.B(n_853),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_865),
.Y(n_870)
);

OAI31xp33_ASAP7_75t_SL g871 ( 
.A1(n_867),
.A2(n_830),
.A3(n_863),
.B(n_853),
.Y(n_871)
);

A2O1A1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_868),
.A2(n_864),
.B(n_848),
.C(n_842),
.Y(n_872)
);

OAI21xp33_ASAP7_75t_L g873 ( 
.A1(n_866),
.A2(n_848),
.B(n_838),
.Y(n_873)
);

HAxp5_ASAP7_75t_SL g874 ( 
.A(n_871),
.B(n_870),
.CON(n_874),
.SN(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_872),
.B(n_869),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_873),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_873),
.B(n_858),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_870),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_876),
.B(n_811),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_878),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_877),
.B(n_811),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_877),
.Y(n_882)
);

OAI221xp5_ASAP7_75t_L g883 ( 
.A1(n_874),
.A2(n_842),
.B1(n_843),
.B2(n_859),
.C(n_858),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_875),
.Y(n_884)
);

OAI322xp33_ASAP7_75t_L g885 ( 
.A1(n_876),
.A2(n_859),
.A3(n_812),
.B1(n_814),
.B2(n_816),
.C1(n_720),
.C2(n_815),
.Y(n_885)
);

NOR2x1_ASAP7_75t_L g886 ( 
.A(n_877),
.B(n_847),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_883),
.A2(n_791),
.B1(n_808),
.B2(n_823),
.Y(n_887)
);

AOI221xp5_ASAP7_75t_L g888 ( 
.A1(n_882),
.A2(n_812),
.B1(n_814),
.B2(n_816),
.C(n_815),
.Y(n_888)
);

OAI211xp5_ASAP7_75t_L g889 ( 
.A1(n_884),
.A2(n_780),
.B(n_822),
.C(n_808),
.Y(n_889)
);

AOI221xp5_ASAP7_75t_L g890 ( 
.A1(n_885),
.A2(n_815),
.B1(n_851),
.B2(n_741),
.C(n_737),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_879),
.A2(n_736),
.B(n_726),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_881),
.A2(n_736),
.B1(n_851),
.B2(n_821),
.Y(n_892)
);

AOI221xp5_ASAP7_75t_L g893 ( 
.A1(n_880),
.A2(n_737),
.B1(n_741),
.B2(n_797),
.C(n_799),
.Y(n_893)
);

OAI221xp5_ASAP7_75t_L g894 ( 
.A1(n_886),
.A2(n_799),
.B1(n_797),
.B2(n_821),
.C(n_802),
.Y(n_894)
);

AOI211xp5_ASAP7_75t_L g895 ( 
.A1(n_883),
.A2(n_726),
.B(n_737),
.C(n_821),
.Y(n_895)
);

NAND2x1p5_ASAP7_75t_L g896 ( 
.A(n_879),
.B(n_726),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_896),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_894),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_895),
.Y(n_899)
);

AOI211xp5_ASAP7_75t_SL g900 ( 
.A1(n_887),
.A2(n_889),
.B(n_890),
.C(n_892),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_891),
.Y(n_901)
);

NOR3xp33_ASAP7_75t_L g902 ( 
.A(n_893),
.B(n_714),
.C(n_731),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_888),
.A2(n_736),
.B1(n_820),
.B2(n_714),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_896),
.B(n_810),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_887),
.B(n_731),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_896),
.Y(n_906)
);

NAND2xp33_ASAP7_75t_SL g907 ( 
.A(n_897),
.B(n_732),
.Y(n_907)
);

AND3x2_ASAP7_75t_L g908 ( 
.A(n_899),
.B(n_906),
.C(n_898),
.Y(n_908)
);

NOR4xp75_ASAP7_75t_L g909 ( 
.A(n_905),
.B(n_735),
.C(n_820),
.D(n_810),
.Y(n_909)
);

NOR3xp33_ASAP7_75t_SL g910 ( 
.A(n_904),
.B(n_104),
.C(n_107),
.Y(n_910)
);

AOI221xp5_ASAP7_75t_L g911 ( 
.A1(n_901),
.A2(n_735),
.B1(n_802),
.B2(n_804),
.C(n_820),
.Y(n_911)
);

AOI211xp5_ASAP7_75t_SL g912 ( 
.A1(n_902),
.A2(n_804),
.B(n_819),
.C(n_117),
.Y(n_912)
);

NAND3xp33_ASAP7_75t_SL g913 ( 
.A(n_901),
.B(n_810),
.C(n_809),
.Y(n_913)
);

INVx4_ASAP7_75t_L g914 ( 
.A(n_900),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_903),
.B(n_809),
.Y(n_915)
);

NAND4xp25_ASAP7_75t_L g916 ( 
.A(n_914),
.B(n_819),
.C(n_805),
.D(n_119),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_907),
.A2(n_805),
.B(n_819),
.Y(n_917)
);

INVxp33_ASAP7_75t_SL g918 ( 
.A(n_908),
.Y(n_918)
);

NOR3xp33_ASAP7_75t_L g919 ( 
.A(n_915),
.B(n_109),
.C(n_114),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_910),
.A2(n_805),
.B1(n_121),
.B2(n_122),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_912),
.B(n_120),
.Y(n_921)
);

NAND4xp75_ASAP7_75t_L g922 ( 
.A(n_911),
.B(n_124),
.C(n_127),
.D(n_128),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_909),
.B(n_129),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_918),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_920),
.Y(n_925)
);

INVxp67_ASAP7_75t_L g926 ( 
.A(n_923),
.Y(n_926)
);

O2A1O1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_921),
.A2(n_913),
.B(n_133),
.C(n_136),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_924),
.Y(n_928)
);

OR2x2_ASAP7_75t_L g929 ( 
.A(n_926),
.B(n_916),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_925),
.B(n_919),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_927),
.A2(n_917),
.B1(n_922),
.B2(n_139),
.Y(n_931)
);

OAI22x1_ASAP7_75t_L g932 ( 
.A1(n_928),
.A2(n_131),
.B1(n_137),
.B2(n_140),
.Y(n_932)
);

NAND3xp33_ASAP7_75t_L g933 ( 
.A(n_930),
.B(n_141),
.C(n_143),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_SL g934 ( 
.A1(n_933),
.A2(n_929),
.B1(n_931),
.B2(n_148),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_932),
.B(n_145),
.Y(n_935)
);

AO221x1_ASAP7_75t_L g936 ( 
.A1(n_934),
.A2(n_146),
.B1(n_149),
.B2(n_150),
.C(n_152),
.Y(n_936)
);

AOI221xp5_ASAP7_75t_L g937 ( 
.A1(n_935),
.A2(n_187),
.B1(n_158),
.B2(n_160),
.C(n_161),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_936),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_937),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_L g940 ( 
.A1(n_938),
.A2(n_939),
.B1(n_162),
.B2(n_166),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_940),
.A2(n_155),
.B1(n_167),
.B2(n_169),
.Y(n_941)
);

AOI211xp5_ASAP7_75t_L g942 ( 
.A1(n_941),
.A2(n_170),
.B(n_172),
.C(n_176),
.Y(n_942)
);


endmodule