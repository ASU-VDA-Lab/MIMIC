module fake_jpeg_705_n_200 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_200);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_200;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_18),
.B(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx4f_ASAP7_75t_SL g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx16f_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_47),
.B1(n_44),
.B2(n_43),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_60),
.B1(n_65),
.B2(n_56),
.Y(n_94)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_81),
.Y(n_93)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_64),
.Y(n_84)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_69),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_85),
.B(n_90),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_81),
.A2(n_51),
.B1(n_74),
.B2(n_61),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_72),
.B1(n_63),
.B2(n_59),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_73),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_57),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_95),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_65),
.B1(n_71),
.B2(n_70),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_58),
.Y(n_95)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_40),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_93),
.A2(n_70),
.B1(n_61),
.B2(n_74),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_101),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_95),
.A2(n_71),
.B1(n_60),
.B2(n_66),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_67),
.C(n_70),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_109),
.C(n_100),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_109),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_65),
.B1(n_68),
.B2(n_63),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_98),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_86),
.A2(n_72),
.B(n_68),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_87),
.B1(n_97),
.B2(n_88),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_39),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_96),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_112),
.B(n_36),
.Y(n_119)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_59),
.C(n_1),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_111),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_118),
.A2(n_134),
.B1(n_136),
.B2(n_6),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_119),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_133),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_127),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_110),
.B(n_0),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_124),
.B(n_128),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_114),
.B(n_0),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_59),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_5),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_1),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_2),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_137),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_3),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_3),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_139),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_117),
.B(n_4),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_4),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_7),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_132),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_159),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_131),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_148),
.C(n_149),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_146),
.B(n_122),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_38),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_152),
.C(n_12),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_125),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_126),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_5),
.B(n_6),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_37),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_153),
.A2(n_154),
.B1(n_158),
.B2(n_161),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_121),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_134),
.A2(n_34),
.B1(n_33),
.B2(n_27),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_132),
.A2(n_25),
.B1(n_21),
.B2(n_10),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_120),
.B(n_8),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_163),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_136),
.A2(n_17),
.B1(n_10),
.B2(n_11),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_160),
.Y(n_165)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_151),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_173),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_157),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_169),
.B(n_174),
.Y(n_180)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_172),
.B(n_175),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_9),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_12),
.C(n_13),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_178),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_150),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_170),
.Y(n_179)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

A2O1A1O1Ixp25_ASAP7_75t_L g182 ( 
.A1(n_166),
.A2(n_143),
.B(n_155),
.C(n_152),
.D(n_161),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_182),
.A2(n_184),
.B1(n_171),
.B2(n_173),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_164),
.B1(n_167),
.B2(n_158),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_189),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_183),
.A2(n_176),
.B1(n_168),
.B2(n_175),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_190),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_181),
.A2(n_177),
.B(n_14),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_191),
.A2(n_185),
.B(n_180),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_194),
.A2(n_191),
.B(n_187),
.Y(n_196)
);

NOR2xp67_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_186),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_L g197 ( 
.A(n_195),
.B(n_196),
.C(n_193),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_197),
.A2(n_179),
.B1(n_14),
.B2(n_15),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_13),
.B(n_15),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_16),
.Y(n_200)
);


endmodule