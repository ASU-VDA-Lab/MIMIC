module fake_jpeg_29400_n_433 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_433);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_433;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_2),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_11),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_54),
.Y(n_95)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_50),
.Y(n_128)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

CKINVDCx9p33_ASAP7_75t_R g53 ( 
.A(n_30),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_53),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_29),
.B(n_0),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_26),
.B(n_11),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_65),
.Y(n_99)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_64),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_36),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_68),
.B(n_73),
.Y(n_116)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_72),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_36),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx4f_ASAP7_75t_SL g138 ( 
.A(n_75),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_26),
.B(n_18),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_78),
.B(n_80),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_36),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_82),
.Y(n_109)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_36),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_38),
.B(n_18),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_38),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_87),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_90),
.B(n_92),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_21),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_94),
.B(n_97),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_21),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_53),
.A2(n_45),
.B1(n_20),
.B2(n_23),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_103),
.B(n_112),
.Y(n_157)
);

AOI21xp33_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_24),
.B(n_23),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_113),
.B(n_122),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_62),
.A2(n_32),
.B1(n_39),
.B2(n_43),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_121),
.A2(n_134),
.B1(n_58),
.B2(n_45),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_85),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_82),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_132),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_69),
.A2(n_32),
.B1(n_39),
.B2(n_43),
.Y(n_134)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

INVx3_ASAP7_75t_SL g197 ( 
.A(n_140),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_83),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_141),
.B(n_150),
.Y(n_193)
);

INVx2_ASAP7_75t_R g142 ( 
.A(n_123),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_142),
.B(n_171),
.Y(n_198)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_102),
.A2(n_66),
.B1(n_71),
.B2(n_77),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_144),
.A2(n_152),
.B1(n_155),
.B2(n_127),
.Y(n_182)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_147),
.Y(n_190)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_149),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_93),
.B(n_24),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_111),
.A2(n_61),
.B(n_81),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_129),
.C(n_114),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_130),
.A2(n_76),
.B1(n_86),
.B2(n_84),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_104),
.A2(n_48),
.B1(n_46),
.B2(n_70),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_153),
.A2(n_158),
.B1(n_160),
.B2(n_164),
.Y(n_191)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_52),
.B1(n_64),
.B2(n_57),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_104),
.A2(n_75),
.B1(n_72),
.B2(n_67),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_96),
.A2(n_75),
.B1(n_72),
.B2(n_50),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_41),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_162),
.B(n_165),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_47),
.B1(n_39),
.B2(n_35),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_163),
.A2(n_137),
.B1(n_135),
.B2(n_127),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_110),
.A2(n_41),
.B1(n_35),
.B2(n_63),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_116),
.B(n_27),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_99),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_166),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_114),
.A2(n_19),
.B1(n_39),
.B2(n_27),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_SL g183 ( 
.A1(n_167),
.A2(n_172),
.B(n_174),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_168),
.Y(n_199)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_125),
.B(n_22),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_173),
.B(n_175),
.Y(n_188)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_95),
.B(n_22),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_177),
.Y(n_215)
);

AND2x4_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_30),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

AO21x2_ASAP7_75t_L g179 ( 
.A1(n_151),
.A2(n_137),
.B(n_138),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_179),
.A2(n_182),
.B1(n_186),
.B2(n_109),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_166),
.B(n_25),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_165),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_157),
.A2(n_91),
.B1(n_108),
.B2(n_120),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_144),
.A2(n_155),
.B1(n_171),
.B2(n_139),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_189),
.A2(n_196),
.B1(n_202),
.B2(n_126),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_142),
.A2(n_120),
.B1(n_108),
.B2(n_117),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_139),
.A2(n_91),
.B1(n_109),
.B2(n_129),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_203),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_212),
.Y(n_235)
);

OAI22x1_ASAP7_75t_SL g207 ( 
.A1(n_179),
.A2(n_142),
.B1(n_140),
.B2(n_162),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_207),
.A2(n_211),
.B1(n_179),
.B2(n_176),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_150),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_214),
.Y(n_240)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_209),
.Y(n_241)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_210),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_178),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_156),
.Y(n_214)
);

AND2x6_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_140),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_218),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_156),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_221),
.Y(n_242)
);

AND2x6_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_175),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_219),
.Y(n_237)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_220),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_177),
.B(n_192),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_222),
.B(n_145),
.Y(n_254)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_223),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_189),
.A2(n_161),
.B1(n_159),
.B2(n_146),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_224),
.A2(n_225),
.B1(n_204),
.B2(n_221),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_182),
.A2(n_161),
.B1(n_169),
.B2(n_172),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_191),
.A2(n_183),
.B1(n_179),
.B2(n_197),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_226),
.A2(n_198),
.B(n_199),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_198),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_227),
.Y(n_244)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_180),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_228),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_230),
.A2(n_233),
.B(n_251),
.Y(n_261)
);

OAI32xp33_ASAP7_75t_L g231 ( 
.A1(n_214),
.A2(n_198),
.A3(n_177),
.B1(n_170),
.B2(n_173),
.Y(n_231)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_231),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_232),
.B(n_247),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_207),
.A2(n_185),
.B1(n_154),
.B2(n_147),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_234),
.A2(n_219),
.B1(n_195),
.B2(n_172),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_188),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_243),
.C(n_225),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_188),
.C(n_181),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_211),
.A2(n_180),
.B1(n_201),
.B2(n_148),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_245),
.A2(n_204),
.B1(n_185),
.B2(n_195),
.Y(n_267)
);

AO22x1_ASAP7_75t_L g247 ( 
.A1(n_227),
.A2(n_197),
.B1(n_201),
.B2(n_200),
.Y(n_247)
);

AOI21xp33_ASAP7_75t_SL g249 ( 
.A1(n_215),
.A2(n_197),
.B(n_30),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_L g264 ( 
.A1(n_249),
.A2(n_209),
.B(n_220),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_222),
.B(n_143),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_213),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_217),
.A2(n_199),
.B(n_200),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_254),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_235),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_255),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_235),
.B(n_206),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_257),
.B(n_239),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_208),
.Y(n_258)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_258),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_224),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_259),
.B(n_274),
.Y(n_301)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_237),
.Y(n_262)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_205),
.Y(n_263)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_263),
.Y(n_290)
);

OAI21xp33_ASAP7_75t_L g288 ( 
.A1(n_264),
.A2(n_242),
.B(n_254),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_247),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_271),
.Y(n_295)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_266),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_267),
.A2(n_280),
.B1(n_234),
.B2(n_236),
.Y(n_300)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_229),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_270),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_260),
.C(n_274),
.Y(n_292)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_246),
.Y(n_270)
);

INVx13_ASAP7_75t_L g271 ( 
.A(n_247),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_229),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_276),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_244),
.B(n_223),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_275),
.B(n_278),
.Y(n_309)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_241),
.Y(n_276)
);

NOR2x1_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_244),
.Y(n_277)
);

NOR2x1_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_273),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_241),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_242),
.B(n_210),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_279),
.B(n_282),
.Y(n_310)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_283),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_231),
.B(n_228),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_232),
.A2(n_218),
.B1(n_216),
.B2(n_190),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_253),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_284),
.B(n_147),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_292),
.Y(n_313)
);

OAI221xp5_ASAP7_75t_L g289 ( 
.A1(n_257),
.A2(n_251),
.B1(n_238),
.B2(n_250),
.C(n_243),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_289),
.B(n_303),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_265),
.A2(n_233),
.B1(n_252),
.B2(n_232),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_256),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_260),
.C(n_261),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_296),
.B(n_302),
.C(n_311),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_255),
.B(n_239),
.Y(n_297)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_297),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_298),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_299),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_300),
.A2(n_304),
.B1(n_307),
.B2(n_306),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_261),
.B(n_246),
.C(n_236),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_263),
.B(n_258),
.Y(n_303)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_305),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_273),
.B(n_148),
.Y(n_306)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_306),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_273),
.B(n_154),
.Y(n_307)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_307),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_283),
.B(n_168),
.C(n_149),
.Y(n_311)
);

NOR3xp33_ASAP7_75t_L g312 ( 
.A(n_277),
.B(n_107),
.C(n_174),
.Y(n_312)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_312),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_315),
.B(n_299),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_256),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_317),
.B(n_303),
.Y(n_352)
);

INVx3_ASAP7_75t_SL g320 ( 
.A(n_308),
.Y(n_320)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_320),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_295),
.A2(n_271),
.B(n_281),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_321),
.A2(n_320),
.B(n_297),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_322),
.Y(n_350)
);

AO22x1_ASAP7_75t_L g323 ( 
.A1(n_298),
.A2(n_280),
.B1(n_284),
.B2(n_276),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_323),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_304),
.A2(n_272),
.B1(n_268),
.B2(n_270),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_325),
.A2(n_329),
.B1(n_332),
.B2(n_300),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_292),
.B(n_266),
.C(n_262),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_326),
.B(n_293),
.C(n_287),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_290),
.A2(n_118),
.B1(n_126),
.B2(n_128),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_296),
.B(n_138),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_330),
.B(n_302),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_290),
.A2(n_118),
.B1(n_106),
.B2(n_105),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_301),
.B(n_105),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_334),
.B(n_305),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_291),
.B(n_106),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_335),
.B(n_287),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_336),
.B(n_338),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_337),
.B(n_340),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_318),
.B(n_309),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_339),
.B(n_342),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_333),
.B(n_310),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_313),
.B(n_330),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_334),
.B(n_311),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_343),
.B(n_344),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_313),
.B(n_293),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_345),
.B(n_348),
.C(n_351),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_346),
.A2(n_335),
.B1(n_321),
.B2(n_325),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_349),
.A2(n_354),
.B1(n_327),
.B2(n_328),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_324),
.B(n_289),
.Y(n_351)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_352),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_324),
.B(n_326),
.C(n_314),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_353),
.B(n_355),
.Y(n_358)
);

INVxp33_ASAP7_75t_SL g354 ( 
.A(n_323),
.Y(n_354)
);

INVxp33_ASAP7_75t_L g372 ( 
.A(n_354),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_315),
.B(n_285),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_331),
.B(n_285),
.C(n_294),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_356),
.B(n_357),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_335),
.B(n_294),
.C(n_286),
.Y(n_357)
);

BUFx24_ASAP7_75t_SL g359 ( 
.A(n_351),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_359),
.B(n_370),
.Y(n_387)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_363),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_341),
.B(n_316),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_365),
.B(n_369),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_367),
.Y(n_379)
);

NOR3xp33_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_298),
.C(n_316),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_345),
.B(n_332),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_355),
.B(n_286),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_373),
.A2(n_342),
.B(n_14),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_349),
.B(n_319),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_374),
.B(n_375),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_357),
.B(n_329),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_361),
.A2(n_350),
.B1(n_347),
.B2(n_348),
.Y(n_376)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_376),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_377),
.B(n_383),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_368),
.A2(n_14),
.B(n_17),
.Y(n_378)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_378),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_362),
.B(n_107),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_380),
.B(n_382),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_362),
.B(n_363),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_360),
.A2(n_13),
.B1(n_17),
.B2(n_16),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_79),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_384),
.B(n_388),
.C(n_375),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_366),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_386),
.B(n_374),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_371),
.B(n_74),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_385),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_391),
.B(n_392),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_387),
.B(n_358),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_393),
.B(n_397),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_389),
.B(n_367),
.Y(n_394)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_394),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_382),
.B(n_372),
.C(n_56),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_399),
.B(n_400),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_379),
.B(n_381),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_380),
.B(n_372),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_401),
.B(n_384),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_395),
.B(n_376),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_402),
.B(n_403),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_398),
.B(n_388),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_404),
.B(n_408),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_396),
.A2(n_9),
.B(n_16),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_405),
.A2(n_397),
.B(n_7),
.Y(n_415)
);

OAI21x1_ASAP7_75t_L g408 ( 
.A1(n_390),
.A2(n_9),
.B(n_16),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_396),
.B(n_8),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_410),
.B(n_6),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_399),
.A2(n_19),
.B(n_7),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_411),
.A2(n_12),
.B(n_15),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_415),
.B(n_416),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_406),
.B(n_6),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_417),
.B(n_418),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_409),
.B(n_12),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_412),
.B(n_12),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_419),
.A2(n_15),
.B(n_407),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_420),
.B(n_407),
.C(n_13),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_421),
.B(n_424),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_414),
.B(n_15),
.C(n_37),
.Y(n_425)
);

OAI21x1_ASAP7_75t_L g428 ( 
.A1(n_425),
.A2(n_0),
.B(n_1),
.Y(n_428)
);

AOI322xp5_ASAP7_75t_L g427 ( 
.A1(n_423),
.A2(n_413),
.A3(n_422),
.B1(n_37),
.B2(n_5),
.C1(n_3),
.C2(n_0),
.Y(n_427)
);

AOI21x1_ASAP7_75t_L g429 ( 
.A1(n_427),
.A2(n_428),
.B(n_426),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_429),
.B(n_0),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_430),
.A2(n_1),
.B(n_3),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_431),
.B(n_37),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_432),
.A2(n_37),
.B(n_197),
.Y(n_433)
);


endmodule