module fake_ariane_1912_n_1762 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1762);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1762;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1252;
wire n_1129;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_11),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_110),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_24),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_13),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_39),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_31),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_32),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_24),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_136),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_64),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_5),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_58),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_91),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_99),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_132),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_52),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_29),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_42),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_32),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_9),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_97),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_9),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_42),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_33),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_96),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_94),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_6),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_18),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_35),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_38),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_65),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_45),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_162),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_43),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_118),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_78),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_16),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_155),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_14),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_62),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_124),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_77),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_148),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_47),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_125),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_2),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_82),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_139),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_30),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_109),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_105),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_128),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_69),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_135),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_86),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_156),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_152),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g225 ( 
.A(n_27),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_39),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_76),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_121),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_2),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_123),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_153),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_101),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_154),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_74),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_88),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_67),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_137),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_119),
.Y(n_238)
);

BUFx5_ASAP7_75t_L g239 ( 
.A(n_55),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_83),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_35),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_51),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_71),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_16),
.Y(n_244)
);

BUFx8_ASAP7_75t_SL g245 ( 
.A(n_100),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_98),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_149),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_53),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_93),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_140),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_56),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_54),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_147),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_8),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_60),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_108),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_7),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_150),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_28),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_46),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_73),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_133),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_30),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_115),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_31),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_111),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_85),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_90),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_61),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_84),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_43),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_46),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_81),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_144),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_122),
.Y(n_275)
);

BUFx8_ASAP7_75t_SL g276 ( 
.A(n_113),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_6),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_23),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_54),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_116),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_75),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_37),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_87),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_33),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_3),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_63),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_59),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_141),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_129),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_72),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_18),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_10),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_57),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_95),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g295 ( 
.A(n_5),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_8),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_0),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_45),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_112),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_104),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_47),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_7),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_51),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_138),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_26),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_70),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_163),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_80),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_103),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_157),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_102),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_106),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_56),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_92),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_23),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_151),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_127),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_29),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_68),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_53),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_114),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_107),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_48),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_145),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_14),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_34),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_130),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_66),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_131),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_44),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_44),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_4),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_17),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_225),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_225),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_225),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_225),
.Y(n_337)
);

NOR2xp67_ASAP7_75t_L g338 ( 
.A(n_182),
.B(n_0),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_245),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_320),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_225),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_193),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_225),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_225),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_225),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_214),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_228),
.B(n_1),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_239),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_276),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_239),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_239),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_164),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_310),
.B(n_1),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_222),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_185),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_224),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_264),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_R g358 ( 
.A(n_205),
.B(n_120),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_311),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_169),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_164),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_204),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_239),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_182),
.B(n_3),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_211),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_213),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_226),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_284),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_239),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_279),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_185),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_239),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_166),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_239),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_241),
.Y(n_375)
);

NAND2xp33_ASAP7_75t_R g376 ( 
.A(n_165),
.B(n_117),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_254),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_209),
.Y(n_378)
);

NOR2xp67_ASAP7_75t_L g379 ( 
.A(n_284),
.B(n_4),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_239),
.B(n_10),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_257),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_257),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_210),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_257),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_176),
.B(n_12),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_257),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_260),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_217),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_166),
.Y(n_389)
);

INVxp33_ASAP7_75t_SL g390 ( 
.A(n_167),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_304),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_304),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_304),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_167),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_257),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_265),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_259),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_220),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_259),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_259),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_259),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_277),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g403 ( 
.A(n_244),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_220),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_278),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_282),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_243),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_259),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_170),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_243),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_170),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_246),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_186),
.Y(n_413)
);

NOR2xp67_ASAP7_75t_L g414 ( 
.A(n_252),
.B(n_12),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_168),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_168),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_305),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_186),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_336),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_334),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_334),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_360),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_335),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_356),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_409),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_381),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_381),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_R g428 ( 
.A(n_339),
.B(n_202),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_349),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_336),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_335),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_411),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_398),
.B(n_244),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_337),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_342),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_337),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_341),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_352),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_382),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_346),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_378),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_R g442 ( 
.A(n_362),
.B(n_207),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_341),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_354),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_357),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_382),
.Y(n_446)
);

BUFx10_ASAP7_75t_L g447 ( 
.A(n_365),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_343),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_343),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_344),
.Y(n_450)
);

AND2x6_ASAP7_75t_L g451 ( 
.A(n_344),
.B(n_177),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_384),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_398),
.B(n_180),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_361),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_345),
.Y(n_455)
);

AND2x4_ASAP7_75t_SL g456 ( 
.A(n_404),
.B(n_295),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_410),
.B(n_165),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_359),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_345),
.Y(n_459)
);

INVx6_ASAP7_75t_L g460 ( 
.A(n_410),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_370),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_348),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_348),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_373),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_384),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_366),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_350),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_386),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_350),
.Y(n_469)
);

OA21x2_ASAP7_75t_L g470 ( 
.A1(n_380),
.A2(n_183),
.B(n_181),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_355),
.B(n_188),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_367),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_351),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_351),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_371),
.B(n_198),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_403),
.B(n_271),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_386),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_368),
.B(n_203),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_363),
.B(n_208),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_395),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_338),
.B(n_271),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_363),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_388),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_395),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_369),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_375),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_369),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_377),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_379),
.B(n_305),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_397),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_397),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_383),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_372),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_372),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_419),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_419),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_430),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_459),
.B(n_387),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_430),
.Y(n_499)
);

AND2x6_ASAP7_75t_L g500 ( 
.A(n_433),
.B(n_177),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_430),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_459),
.B(n_396),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_419),
.Y(n_503)
);

NAND2xp33_ASAP7_75t_SL g504 ( 
.A(n_466),
.B(n_358),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_446),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_446),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_433),
.B(n_413),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_419),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_446),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_L g510 ( 
.A1(n_470),
.A2(n_364),
.B1(n_347),
.B2(n_353),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_453),
.B(n_390),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_481),
.B(n_402),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_460),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_460),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_441),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_471),
.B(n_405),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_481),
.B(n_406),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_446),
.Y(n_518)
);

NOR2x1p5_ASAP7_75t_L g519 ( 
.A(n_472),
.B(n_418),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_459),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_459),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_420),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_420),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_475),
.B(n_385),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_446),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_421),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_421),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_423),
.B(n_389),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_423),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_470),
.A2(n_414),
.B1(n_330),
.B2(n_195),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_447),
.B(n_227),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_431),
.B(n_394),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_431),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_460),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_434),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_486),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_434),
.Y(n_537)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_492),
.B(n_340),
.Y(n_538)
);

AO21x2_ASAP7_75t_L g539 ( 
.A1(n_457),
.A2(n_238),
.B(n_237),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_436),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_447),
.B(n_240),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_481),
.B(n_489),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_436),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_460),
.B(n_407),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_437),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_437),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_438),
.B(n_454),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_447),
.B(n_249),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_446),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_443),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_443),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_470),
.A2(n_451),
.B1(n_489),
.B2(n_476),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_448),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_447),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_481),
.B(n_412),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_470),
.A2(n_285),
.B1(n_292),
.B2(n_302),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_448),
.B(n_374),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_449),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_452),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_449),
.Y(n_560)
);

NAND3xp33_ASAP7_75t_L g561 ( 
.A(n_488),
.B(n_376),
.C(n_190),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_442),
.B(n_256),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_452),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_452),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_450),
.Y(n_565)
);

BUFx10_ASAP7_75t_L g566 ( 
.A(n_429),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_450),
.B(n_374),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_455),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_455),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_462),
.B(n_399),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_492),
.B(n_174),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_462),
.B(n_399),
.Y(n_572)
);

OR2x6_ASAP7_75t_L g573 ( 
.A(n_432),
.B(n_425),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_L g574 ( 
.A(n_463),
.B(n_467),
.Y(n_574)
);

INVxp33_ASAP7_75t_L g575 ( 
.A(n_432),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_463),
.B(n_415),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_424),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_451),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_452),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_464),
.B(n_391),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_467),
.B(n_469),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_469),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_473),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_473),
.B(n_400),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_474),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_474),
.B(n_400),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_482),
.B(n_415),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_489),
.B(n_416),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_452),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_422),
.Y(n_590)
);

AND3x2_ASAP7_75t_L g591 ( 
.A(n_476),
.B(n_184),
.C(n_171),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_489),
.B(n_416),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_452),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_482),
.B(n_261),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_478),
.B(n_417),
.Y(n_595)
);

BUFx10_ASAP7_75t_L g596 ( 
.A(n_456),
.Y(n_596)
);

NOR3xp33_ASAP7_75t_L g597 ( 
.A(n_435),
.B(n_263),
.C(n_206),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_485),
.B(n_401),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g599 ( 
.A(n_440),
.Y(n_599)
);

INVxp33_ASAP7_75t_L g600 ( 
.A(n_428),
.Y(n_600)
);

INVx6_ASAP7_75t_L g601 ( 
.A(n_484),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_487),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_487),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_444),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_493),
.B(n_401),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_493),
.B(n_408),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_494),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_451),
.A2(n_323),
.B1(n_296),
.B2(n_189),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_456),
.B(n_187),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_494),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_456),
.B(n_187),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_484),
.Y(n_612)
);

AND2x6_ASAP7_75t_L g613 ( 
.A(n_426),
.B(n_234),
.Y(n_613)
);

INVx4_ASAP7_75t_L g614 ( 
.A(n_451),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_479),
.B(n_417),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_451),
.B(n_408),
.Y(n_616)
);

BUFx4f_ASAP7_75t_L g617 ( 
.A(n_451),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_445),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_426),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_484),
.B(n_266),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_451),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_427),
.B(n_268),
.Y(n_622)
);

NOR2x1p5_ASAP7_75t_L g623 ( 
.A(n_458),
.B(n_190),
.Y(n_623)
);

INVx8_ASAP7_75t_L g624 ( 
.A(n_483),
.Y(n_624)
);

NAND3xp33_ASAP7_75t_L g625 ( 
.A(n_427),
.B(n_201),
.C(n_196),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_491),
.A2(n_301),
.B1(n_194),
.B2(n_332),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_439),
.B(n_274),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_439),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_465),
.B(n_230),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_465),
.B(n_275),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_468),
.B(n_197),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_468),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_477),
.B(n_199),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_484),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_477),
.B(n_191),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_480),
.B(n_231),
.Y(n_636)
);

NOR2x1p5_ASAP7_75t_L g637 ( 
.A(n_461),
.B(n_191),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_480),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_484),
.B(n_281),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_491),
.Y(n_640)
);

NAND3xp33_ASAP7_75t_L g641 ( 
.A(n_484),
.B(n_301),
.C(n_196),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_490),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_490),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_490),
.B(n_250),
.Y(n_644)
);

INVx4_ASAP7_75t_L g645 ( 
.A(n_490),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_497),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_524),
.B(n_392),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_514),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_556),
.A2(n_530),
.B1(n_500),
.B2(n_552),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_524),
.B(n_393),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_546),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_514),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_542),
.B(n_295),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_554),
.B(n_172),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_534),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_511),
.B(n_194),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_554),
.B(n_172),
.Y(n_657)
);

O2A1O1Ixp33_ASAP7_75t_L g658 ( 
.A1(n_581),
.A2(n_574),
.B(n_502),
.C(n_498),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_614),
.B(n_173),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_546),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_497),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_511),
.B(n_201),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_542),
.B(n_295),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_516),
.B(n_294),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_516),
.A2(n_319),
.B1(n_200),
.B2(n_192),
.Y(n_665)
);

OAI22xp33_ASAP7_75t_L g666 ( 
.A1(n_575),
.A2(n_313),
.B1(n_298),
.B2(n_332),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_551),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_510),
.A2(n_313),
.B1(n_298),
.B2(n_331),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_614),
.B(n_173),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_590),
.B(n_297),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_615),
.B(n_317),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_574),
.A2(n_319),
.B(n_327),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_615),
.B(n_528),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_SL g674 ( 
.A(n_577),
.B(n_297),
.Y(n_674)
);

NOR2x1p5_ASAP7_75t_L g675 ( 
.A(n_609),
.B(n_318),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_542),
.B(n_216),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_615),
.B(n_321),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_614),
.B(n_520),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_520),
.B(n_175),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_528),
.B(n_532),
.Y(n_680)
);

O2A1O1Ixp33_ASAP7_75t_L g681 ( 
.A1(n_498),
.A2(n_303),
.B(n_333),
.C(n_272),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_547),
.B(n_318),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_558),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_532),
.B(n_175),
.Y(n_684)
);

NOR2x1p5_ASAP7_75t_L g685 ( 
.A(n_611),
.B(n_325),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_595),
.B(n_178),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_595),
.B(n_500),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_499),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_600),
.B(n_325),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_595),
.B(n_178),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_499),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_521),
.B(n_179),
.Y(n_692)
);

NOR3xp33_ASAP7_75t_L g693 ( 
.A(n_536),
.B(n_229),
.C(n_242),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_515),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_521),
.B(n_578),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_500),
.B(n_192),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_500),
.B(n_200),
.Y(n_697)
);

NAND3xp33_ASAP7_75t_L g698 ( 
.A(n_510),
.B(n_331),
.C(n_309),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_500),
.B(n_235),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_600),
.B(n_235),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_575),
.B(n_290),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_555),
.B(n_290),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_604),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_607),
.B(n_293),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_578),
.B(n_293),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_527),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_501),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_588),
.B(n_299),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_534),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_501),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_533),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_502),
.B(n_299),
.Y(n_712)
);

OAI21xp5_ASAP7_75t_L g713 ( 
.A1(n_567),
.A2(n_307),
.B(n_308),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_540),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_621),
.B(n_300),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_588),
.B(n_300),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_531),
.B(n_309),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_531),
.A2(n_312),
.B1(n_329),
.B2(n_328),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_588),
.B(n_312),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_592),
.B(n_314),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_543),
.Y(n_721)
);

NOR2xp67_ASAP7_75t_L g722 ( 
.A(n_599),
.B(n_314),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_522),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_561),
.B(n_617),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_557),
.A2(n_322),
.B(n_324),
.Y(n_725)
);

OAI21xp5_ASAP7_75t_L g726 ( 
.A1(n_567),
.A2(n_234),
.B(n_269),
.Y(n_726)
);

OAI22xp33_ASAP7_75t_L g727 ( 
.A1(n_573),
.A2(n_291),
.B1(n_248),
.B2(n_315),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_522),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_SL g729 ( 
.A1(n_580),
.A2(n_326),
.B1(n_251),
.B2(n_328),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_592),
.B(n_329),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_617),
.B(n_255),
.Y(n_731)
);

NAND2xp33_ASAP7_75t_L g732 ( 
.A(n_523),
.B(n_221),
.Y(n_732)
);

NAND2xp33_ASAP7_75t_SL g733 ( 
.A(n_519),
.B(n_255),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_544),
.B(n_507),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_541),
.A2(n_548),
.B1(n_504),
.B2(n_512),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_541),
.A2(n_262),
.B1(n_215),
.B2(n_218),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_538),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_517),
.B(n_316),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_523),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_548),
.A2(n_267),
.B1(n_219),
.B2(n_223),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_508),
.B(n_270),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_513),
.B(n_232),
.Y(n_742)
);

OAI221xp5_ASAP7_75t_L g743 ( 
.A1(n_626),
.A2(n_273),
.B1(n_316),
.B2(n_269),
.C(n_289),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_556),
.A2(n_530),
.B1(n_552),
.B2(n_608),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_571),
.B(n_212),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_545),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_508),
.B(n_233),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_573),
.Y(n_748)
);

NAND2xp33_ASAP7_75t_L g749 ( 
.A(n_526),
.B(n_221),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_562),
.B(n_236),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_562),
.B(n_247),
.Y(n_751)
);

AND2x4_ASAP7_75t_SL g752 ( 
.A(n_596),
.B(n_490),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_553),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_560),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_565),
.B(n_283),
.Y(n_755)
);

INVxp67_ASAP7_75t_L g756 ( 
.A(n_573),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_526),
.B(n_273),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_596),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_504),
.B(n_253),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_568),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_569),
.B(n_286),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_582),
.B(n_288),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_583),
.B(n_287),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_585),
.B(n_280),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_539),
.B(n_258),
.Y(n_765)
);

INVx1_ASAP7_75t_SL g766 ( 
.A(n_618),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_566),
.B(n_13),
.Y(n_767)
);

OR2x2_ASAP7_75t_L g768 ( 
.A(n_624),
.B(n_15),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_529),
.B(n_306),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_535),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_535),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_539),
.B(n_15),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_602),
.B(n_289),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_603),
.B(n_246),
.Y(n_774)
);

NOR2xp67_ASAP7_75t_L g775 ( 
.A(n_641),
.B(n_126),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_537),
.B(n_306),
.Y(n_776)
);

INVx1_ASAP7_75t_SL g777 ( 
.A(n_624),
.Y(n_777)
);

OR2x2_ASAP7_75t_SL g778 ( 
.A(n_624),
.B(n_596),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_610),
.B(n_17),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_537),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_576),
.B(n_19),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_550),
.A2(n_306),
.B1(n_221),
.B2(n_21),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_550),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_566),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_505),
.B(n_306),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_566),
.B(n_19),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_576),
.B(n_20),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_645),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_594),
.A2(n_306),
.B1(n_221),
.B2(n_22),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_587),
.B(n_20),
.Y(n_790)
);

OAI21xp5_ASAP7_75t_L g791 ( 
.A1(n_495),
.A2(n_221),
.B(n_161),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_587),
.B(n_21),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_601),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_638),
.B(n_22),
.Y(n_794)
);

NAND3xp33_ASAP7_75t_L g795 ( 
.A(n_625),
.B(n_25),
.C(n_26),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_629),
.B(n_25),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_505),
.B(n_27),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_635),
.B(n_28),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_496),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_636),
.B(n_34),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_503),
.Y(n_801)
);

OAI21xp5_ASAP7_75t_L g802 ( 
.A1(n_594),
.A2(n_642),
.B(n_570),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_601),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_619),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_631),
.B(n_36),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_628),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_631),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_505),
.B(n_40),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_505),
.B(n_40),
.Y(n_809)
);

BUFx8_ASAP7_75t_L g810 ( 
.A(n_784),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_703),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_678),
.A2(n_695),
.B(n_658),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_648),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_647),
.B(n_645),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_680),
.B(n_633),
.Y(n_815)
);

AOI21x1_ASAP7_75t_L g816 ( 
.A1(n_695),
.A2(n_644),
.B(n_632),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_650),
.B(n_645),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_646),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_678),
.A2(n_642),
.B(n_598),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_648),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_656),
.A2(n_623),
.B1(n_643),
.B2(n_633),
.Y(n_821)
);

OAI21xp5_ASAP7_75t_L g822 ( 
.A1(n_802),
.A2(n_572),
.B(n_584),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_659),
.A2(n_589),
.B(n_579),
.Y(n_823)
);

O2A1O1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_662),
.A2(n_586),
.B(n_605),
.C(n_606),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_664),
.B(n_631),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_659),
.A2(n_669),
.B(n_705),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_673),
.B(n_633),
.Y(n_827)
);

OA21x2_ASAP7_75t_L g828 ( 
.A1(n_791),
.A2(n_616),
.B(n_640),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_669),
.A2(n_593),
.B(n_634),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_717),
.A2(n_627),
.B1(n_630),
.B2(n_622),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_684),
.B(n_608),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_705),
.A2(n_593),
.B(n_634),
.Y(n_832)
);

O2A1O1Ixp33_ASAP7_75t_SL g833 ( 
.A1(n_781),
.A2(n_639),
.B(n_620),
.C(n_627),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_L g834 ( 
.A1(n_649),
.A2(n_579),
.B1(n_564),
.B2(n_589),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_712),
.A2(n_630),
.B1(n_622),
.B2(n_637),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_715),
.A2(n_612),
.B(n_639),
.Y(n_836)
);

AOI21x1_ASAP7_75t_L g837 ( 
.A1(n_731),
.A2(n_620),
.B(n_601),
.Y(n_837)
);

AOI21x1_ASAP7_75t_L g838 ( 
.A1(n_731),
.A2(n_549),
.B(n_509),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_671),
.B(n_591),
.Y(n_839)
);

OR2x2_ASAP7_75t_SL g840 ( 
.A(n_768),
.B(n_597),
.Y(n_840)
);

OR2x2_ASAP7_75t_L g841 ( 
.A(n_737),
.B(n_563),
.Y(n_841)
);

O2A1O1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_668),
.A2(n_41),
.B(n_48),
.C(n_49),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_741),
.A2(n_525),
.B(n_563),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_747),
.A2(n_559),
.B(n_549),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_744),
.A2(n_559),
.B1(n_509),
.B2(n_518),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_801),
.A2(n_559),
.B(n_549),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_734),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_735),
.B(n_559),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_677),
.B(n_525),
.Y(n_849)
);

CKINVDCx10_ASAP7_75t_R g850 ( 
.A(n_703),
.Y(n_850)
);

O2A1O1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_787),
.A2(n_41),
.B(n_49),
.C(n_50),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_801),
.A2(n_518),
.B(n_509),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_651),
.B(n_655),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_723),
.A2(n_518),
.B(n_506),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_723),
.A2(n_518),
.B(n_506),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_702),
.B(n_660),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_700),
.B(n_506),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_728),
.A2(n_506),
.B(n_613),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_652),
.Y(n_859)
);

A2O1A1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_713),
.A2(n_798),
.B(n_698),
.C(n_772),
.Y(n_860)
);

O2A1O1Ixp5_ASAP7_75t_L g861 ( 
.A1(n_790),
.A2(n_613),
.B(n_52),
.C(n_55),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_745),
.B(n_613),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_652),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_793),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_667),
.B(n_50),
.Y(n_865)
);

BUFx4f_ASAP7_75t_L g866 ( 
.A(n_758),
.Y(n_866)
);

A2O1A1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_807),
.A2(n_726),
.B(n_665),
.C(n_792),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_739),
.A2(n_79),
.B(n_89),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_784),
.Y(n_869)
);

OR2x2_ASAP7_75t_L g870 ( 
.A(n_670),
.B(n_142),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_711),
.B(n_143),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_682),
.B(n_160),
.Y(n_872)
);

INVx4_ASAP7_75t_L g873 ( 
.A(n_651),
.Y(n_873)
);

O2A1O1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_797),
.A2(n_809),
.B(n_808),
.C(n_666),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_770),
.A2(n_771),
.B(n_783),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_661),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_766),
.B(n_694),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_714),
.B(n_721),
.Y(n_878)
);

AOI21x1_ASAP7_75t_L g879 ( 
.A1(n_724),
.A2(n_757),
.B(n_769),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_770),
.A2(n_771),
.B(n_783),
.Y(n_880)
);

BUFx8_ASAP7_75t_L g881 ( 
.A(n_767),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_746),
.B(n_753),
.Y(n_882)
);

OR2x2_ASAP7_75t_L g883 ( 
.A(n_748),
.B(n_756),
.Y(n_883)
);

AOI21xp33_ASAP7_75t_L g884 ( 
.A1(n_701),
.A2(n_750),
.B(n_751),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_780),
.A2(n_704),
.B(n_799),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_754),
.B(n_760),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_674),
.B(n_653),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_759),
.B(n_689),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_793),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_780),
.A2(n_764),
.B(n_755),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_676),
.B(n_686),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_676),
.B(n_690),
.Y(n_892)
);

O2A1O1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_797),
.A2(n_809),
.B(n_808),
.C(n_654),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_672),
.A2(n_681),
.B(n_789),
.C(n_729),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_777),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_796),
.A2(n_800),
.B(n_804),
.Y(n_896)
);

NOR3xp33_ASAP7_75t_L g897 ( 
.A(n_733),
.B(n_693),
.C(n_795),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_806),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_806),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_786),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_683),
.B(n_653),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_663),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_724),
.A2(n_725),
.B(n_692),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_761),
.A2(n_763),
.B(n_762),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_663),
.B(n_655),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_709),
.B(n_742),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_687),
.A2(n_709),
.B1(n_654),
.B2(n_657),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_661),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_803),
.A2(n_738),
.B(n_657),
.Y(n_909)
);

AOI21x1_ASAP7_75t_L g910 ( 
.A1(n_757),
.A2(n_776),
.B(n_769),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_758),
.B(n_716),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_679),
.A2(n_692),
.B(n_707),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_708),
.B(n_719),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_720),
.B(n_730),
.Y(n_914)
);

INVx1_ASAP7_75t_SL g915 ( 
.A(n_733),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_722),
.B(n_805),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_688),
.A2(n_710),
.B(n_691),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_778),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_688),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_779),
.A2(n_718),
.B1(n_696),
.B2(n_697),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_691),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_675),
.B(n_685),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_L g923 ( 
.A1(n_765),
.A2(n_743),
.B1(n_707),
.B2(n_710),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_699),
.A2(n_773),
.B(n_774),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_732),
.A2(n_749),
.B(n_794),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_727),
.B(n_775),
.Y(n_926)
);

AOI21x1_ASAP7_75t_L g927 ( 
.A1(n_785),
.A2(n_782),
.B(n_749),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_752),
.B(n_736),
.Y(n_928)
);

BUFx12f_ASAP7_75t_L g929 ( 
.A(n_740),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_706),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_735),
.B(n_651),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_680),
.B(n_664),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_703),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_706),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_735),
.B(n_651),
.Y(n_935)
);

O2A1O1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_680),
.A2(n_662),
.B(n_656),
.C(n_668),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_680),
.B(n_664),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_680),
.B(n_664),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_706),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_735),
.B(n_651),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_680),
.B(n_664),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_678),
.A2(n_695),
.B(n_574),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_682),
.B(n_547),
.Y(n_943)
);

BUFx2_ASAP7_75t_L g944 ( 
.A(n_703),
.Y(n_944)
);

CKINVDCx20_ASAP7_75t_R g945 ( 
.A(n_703),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_678),
.A2(n_695),
.B(n_574),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_735),
.B(n_651),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_680),
.B(n_664),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_646),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_735),
.B(n_651),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_682),
.B(n_547),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_735),
.B(n_651),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_680),
.A2(n_713),
.B(n_656),
.C(n_662),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_680),
.B(n_664),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_680),
.B(n_664),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_682),
.B(n_547),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_680),
.B(n_664),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_647),
.B(n_650),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_678),
.A2(n_695),
.B(n_802),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_678),
.A2(n_695),
.B(n_802),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_680),
.A2(n_662),
.B(n_656),
.C(n_668),
.Y(n_961)
);

OAI21x1_ASAP7_75t_L g962 ( 
.A1(n_802),
.A2(n_661),
.B(n_646),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_678),
.A2(n_695),
.B(n_574),
.Y(n_963)
);

AO21x1_ASAP7_75t_L g964 ( 
.A1(n_791),
.A2(n_726),
.B(n_772),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_680),
.A2(n_662),
.B(n_656),
.C(n_668),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_678),
.A2(n_695),
.B(n_574),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_678),
.A2(n_695),
.B(n_574),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_680),
.B(n_664),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_706),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_646),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_706),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_647),
.B(n_650),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_678),
.A2(n_695),
.B(n_574),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_735),
.B(n_651),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_646),
.Y(n_975)
);

AO21x1_ASAP7_75t_L g976 ( 
.A1(n_791),
.A2(n_726),
.B(n_772),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_678),
.A2(n_695),
.B(n_574),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_818),
.Y(n_978)
);

O2A1O1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_953),
.A2(n_936),
.B(n_961),
.C(n_965),
.Y(n_979)
);

NOR2x1_ASAP7_75t_SL g980 ( 
.A(n_931),
.B(n_935),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_932),
.B(n_937),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_810),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_930),
.Y(n_983)
);

INVxp33_ASAP7_75t_L g984 ( 
.A(n_877),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_953),
.A2(n_860),
.B(n_972),
.C(n_958),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_938),
.B(n_941),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_820),
.Y(n_987)
);

OAI21xp33_ASAP7_75t_L g988 ( 
.A1(n_958),
.A2(n_972),
.B(n_954),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_810),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_948),
.B(n_955),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_962),
.A2(n_812),
.B(n_838),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_SL g992 ( 
.A1(n_860),
.A2(n_867),
.B(n_815),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_904),
.A2(n_976),
.B(n_964),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_884),
.A2(n_867),
.B(n_968),
.C(n_957),
.Y(n_994)
);

OA22x2_ASAP7_75t_L g995 ( 
.A1(n_835),
.A2(n_821),
.B1(n_902),
.B2(n_887),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_888),
.B(n_913),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_L g997 ( 
.A1(n_827),
.A2(n_892),
.B1(n_891),
.B2(n_831),
.Y(n_997)
);

AO21x1_ASAP7_75t_L g998 ( 
.A1(n_893),
.A2(n_947),
.B(n_940),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_873),
.Y(n_999)
);

OAI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_830),
.A2(n_946),
.B(n_942),
.Y(n_1000)
);

AO31x2_ASAP7_75t_L g1001 ( 
.A1(n_845),
.A2(n_920),
.A3(n_890),
.B(n_924),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_L g1002 ( 
.A1(n_879),
.A2(n_816),
.B(n_917),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_L g1003 ( 
.A1(n_875),
.A2(n_880),
.B(n_837),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_943),
.B(n_951),
.Y(n_1004)
);

OAI21x1_ASAP7_75t_L g1005 ( 
.A1(n_959),
.A2(n_960),
.B(n_844),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_811),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_820),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_963),
.A2(n_977),
.B(n_966),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_967),
.A2(n_973),
.B(n_885),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_940),
.A2(n_952),
.B(n_950),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_926),
.A2(n_825),
.B1(n_897),
.B2(n_929),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_956),
.B(n_847),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_869),
.B(n_918),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_847),
.B(n_856),
.Y(n_1014)
);

INVx2_ASAP7_75t_SL g1015 ( 
.A(n_850),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_843),
.A2(n_910),
.B(n_858),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_934),
.Y(n_1017)
);

NAND2x1p5_ASAP7_75t_L g1018 ( 
.A(n_859),
.B(n_820),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_939),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_933),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_820),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_947),
.A2(n_952),
.B(n_974),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_863),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_950),
.A2(n_974),
.B(n_814),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_SL g1025 ( 
.A1(n_868),
.A2(n_862),
.B(n_926),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_876),
.Y(n_1026)
);

INVxp67_ASAP7_75t_L g1027 ( 
.A(n_841),
.Y(n_1027)
);

INVxp67_ASAP7_75t_L g1028 ( 
.A(n_865),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_856),
.B(n_814),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_817),
.B(n_914),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_921),
.Y(n_1031)
);

AOI21x1_ASAP7_75t_L g1032 ( 
.A1(n_848),
.A2(n_826),
.B(n_925),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_817),
.A2(n_906),
.B(n_833),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_854),
.A2(n_855),
.B(n_846),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_944),
.B(n_900),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_895),
.A2(n_897),
.B1(n_915),
.B2(n_872),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_969),
.Y(n_1037)
);

INVx8_ASAP7_75t_L g1038 ( 
.A(n_864),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_883),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_874),
.A2(n_842),
.B(n_894),
.C(n_861),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_852),
.A2(n_912),
.B(n_819),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_833),
.A2(n_857),
.B(n_896),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_834),
.A2(n_903),
.B(n_824),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_907),
.B(n_873),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_971),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_878),
.B(n_882),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_822),
.A2(n_848),
.B(n_916),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_823),
.A2(n_829),
.B(n_927),
.Y(n_1048)
);

NAND2x1p5_ASAP7_75t_L g1049 ( 
.A(n_859),
.B(n_863),
.Y(n_1049)
);

NOR2xp67_ASAP7_75t_SL g1050 ( 
.A(n_918),
.B(n_922),
.Y(n_1050)
);

NAND3xp33_ASAP7_75t_L g1051 ( 
.A(n_894),
.B(n_851),
.C(n_865),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_836),
.A2(n_909),
.B(n_832),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_863),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_853),
.A2(n_871),
.B(n_886),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_901),
.B(n_839),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_864),
.Y(n_1056)
);

NAND2x1p5_ASAP7_75t_L g1057 ( 
.A(n_813),
.B(n_864),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_928),
.B(n_919),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_905),
.B(n_911),
.Y(n_1059)
);

AO31x2_ASAP7_75t_L g1060 ( 
.A1(n_898),
.A2(n_899),
.A3(n_908),
.B(n_949),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_881),
.Y(n_1061)
);

INVx5_ASAP7_75t_L g1062 ( 
.A(n_864),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_828),
.A2(n_849),
.B(n_975),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_919),
.B(n_923),
.Y(n_1064)
);

OAI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_861),
.A2(n_923),
.B(n_970),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_SL g1066 ( 
.A1(n_870),
.A2(n_828),
.B(n_866),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_889),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_919),
.A2(n_840),
.B(n_881),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_962),
.A2(n_812),
.B(n_838),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_953),
.B(n_860),
.Y(n_1070)
);

NAND2x1p5_ASAP7_75t_L g1071 ( 
.A(n_859),
.B(n_648),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_SL g1072 ( 
.A1(n_874),
.A2(n_893),
.B(n_961),
.Y(n_1072)
);

NAND2x1_ASAP7_75t_L g1073 ( 
.A(n_873),
.B(n_788),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_936),
.A2(n_961),
.B(n_965),
.C(n_953),
.Y(n_1074)
);

AO21x1_ASAP7_75t_L g1075 ( 
.A1(n_888),
.A2(n_961),
.B(n_936),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_930),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_SL g1077 ( 
.A1(n_874),
.A2(n_893),
.B(n_961),
.Y(n_1077)
);

INVx8_ASAP7_75t_L g1078 ( 
.A(n_945),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_943),
.B(n_951),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_962),
.A2(n_812),
.B(n_838),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_820),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_818),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_932),
.B(n_937),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_953),
.A2(n_904),
.B(n_964),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_932),
.B(n_937),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_932),
.B(n_937),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_818),
.Y(n_1087)
);

OR2x6_ASAP7_75t_L g1088 ( 
.A(n_877),
.B(n_624),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_850),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_818),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_930),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_953),
.A2(n_961),
.B(n_936),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_930),
.Y(n_1093)
);

AOI21xp33_ASAP7_75t_L g1094 ( 
.A1(n_936),
.A2(n_662),
.B(n_656),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_818),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_953),
.A2(n_961),
.B(n_936),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_953),
.A2(n_904),
.B(n_964),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_877),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_810),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_953),
.A2(n_936),
.B1(n_965),
.B2(n_961),
.Y(n_1100)
);

AOI21xp33_ASAP7_75t_L g1101 ( 
.A1(n_936),
.A2(n_662),
.B(n_656),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_932),
.B(n_937),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_932),
.B(n_937),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_953),
.A2(n_904),
.B(n_964),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_962),
.A2(n_812),
.B(n_838),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_953),
.A2(n_904),
.B(n_964),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_932),
.B(n_937),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_953),
.A2(n_904),
.B(n_964),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_869),
.B(n_918),
.Y(n_1109)
);

AOI21x1_ASAP7_75t_L g1110 ( 
.A1(n_848),
.A2(n_838),
.B(n_964),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_930),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_818),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_958),
.B(n_647),
.Y(n_1113)
);

OAI22x1_ASAP7_75t_L g1114 ( 
.A1(n_835),
.A2(n_972),
.B1(n_958),
.B2(n_435),
.Y(n_1114)
);

INVx1_ASAP7_75t_SL g1115 ( 
.A(n_877),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_943),
.B(n_951),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_869),
.B(n_918),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_930),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_932),
.B(n_937),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_988),
.B(n_1029),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_987),
.Y(n_1121)
);

BUFx10_ASAP7_75t_L g1122 ( 
.A(n_1089),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_983),
.Y(n_1123)
);

O2A1O1Ixp5_ASAP7_75t_SL g1124 ( 
.A1(n_1070),
.A2(n_1100),
.B(n_1101),
.C(n_1094),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_1061),
.Y(n_1125)
);

BUFx10_ASAP7_75t_L g1126 ( 
.A(n_1015),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1127)
);

AOI21xp33_ASAP7_75t_L g1128 ( 
.A1(n_1051),
.A2(n_1113),
.B(n_979),
.Y(n_1128)
);

OR2x2_ASAP7_75t_SL g1129 ( 
.A(n_1014),
.B(n_1039),
.Y(n_1129)
);

O2A1O1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_985),
.A2(n_1113),
.B(n_994),
.C(n_1074),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1004),
.B(n_1079),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_996),
.B(n_981),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_R g1133 ( 
.A(n_1078),
.B(n_982),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1134)
);

AOI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1114),
.A2(n_996),
.B1(n_1028),
.B2(n_985),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_1062),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1017),
.Y(n_1137)
);

O2A1O1Ixp5_ASAP7_75t_SL g1138 ( 
.A1(n_1070),
.A2(n_1096),
.B(n_1092),
.C(n_1058),
.Y(n_1138)
);

OR2x6_ASAP7_75t_L g1139 ( 
.A(n_1088),
.B(n_1038),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1078),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_1117),
.B(n_1068),
.Y(n_1141)
);

O2A1O1Ixp5_ASAP7_75t_L g1142 ( 
.A1(n_1075),
.A2(n_1074),
.B(n_1097),
.C(n_1104),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1019),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_1062),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1037),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_1115),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1045),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_986),
.B(n_990),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1083),
.B(n_1085),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1028),
.A2(n_994),
.B1(n_1107),
.B2(n_1103),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1116),
.B(n_1012),
.Y(n_1151)
);

INVxp67_ASAP7_75t_SL g1152 ( 
.A(n_1046),
.Y(n_1152)
);

INVx4_ASAP7_75t_SL g1153 ( 
.A(n_982),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_1036),
.B(n_1030),
.Y(n_1154)
);

INVx4_ASAP7_75t_L g1155 ( 
.A(n_1078),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1086),
.B(n_1102),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1119),
.B(n_1098),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_995),
.A2(n_984),
.B1(n_1011),
.B2(n_1055),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1039),
.B(n_997),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1011),
.A2(n_995),
.B1(n_997),
.B2(n_1088),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1117),
.B(n_1062),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_992),
.B(n_980),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1059),
.B(n_984),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_979),
.A2(n_1043),
.B(n_1025),
.Y(n_1164)
);

OAI21xp33_ASAP7_75t_L g1165 ( 
.A1(n_1040),
.A2(n_1108),
.B(n_1106),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_SL g1166 ( 
.A(n_1050),
.B(n_989),
.Y(n_1166)
);

AOI21xp33_ASAP7_75t_L g1167 ( 
.A1(n_1072),
.A2(n_1077),
.B(n_1040),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1076),
.Y(n_1168)
);

OR2x6_ASAP7_75t_L g1169 ( 
.A(n_1088),
.B(n_1038),
.Y(n_1169)
);

NAND2x1p5_ASAP7_75t_L g1170 ( 
.A(n_1062),
.B(n_989),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_987),
.Y(n_1171)
);

INVx1_ASAP7_75t_SL g1172 ( 
.A(n_1035),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_1026),
.A2(n_1082),
.B1(n_1112),
.B2(n_1031),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_1099),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_1099),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_1006),
.B(n_1020),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_SL g1177 ( 
.A1(n_1084),
.A2(n_1108),
.B(n_1106),
.C(n_1097),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1038),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_1027),
.B(n_1091),
.Y(n_1179)
);

NAND2xp33_ASAP7_75t_L g1180 ( 
.A(n_999),
.B(n_1000),
.Y(n_1180)
);

OR2x2_ASAP7_75t_L g1181 ( 
.A(n_1027),
.B(n_1093),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1111),
.B(n_1118),
.Y(n_1182)
);

OR2x6_ASAP7_75t_L g1183 ( 
.A(n_1018),
.B(n_1049),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1024),
.A2(n_1104),
.B(n_1084),
.C(n_1010),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1087),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_987),
.Y(n_1186)
);

OAI21xp33_ASAP7_75t_L g1187 ( 
.A1(n_1033),
.A2(n_1024),
.B(n_993),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_991),
.A2(n_1080),
.B(n_1105),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1044),
.A2(n_1033),
.B(n_1009),
.Y(n_1189)
);

INVx5_ASAP7_75t_L g1190 ( 
.A(n_987),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1067),
.B(n_1071),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1090),
.A2(n_1095),
.B1(n_1058),
.B2(n_1064),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1053),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1010),
.A2(n_1022),
.B1(n_1044),
.B2(n_993),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1022),
.B(n_1053),
.Y(n_1195)
);

NAND3xp33_ASAP7_75t_L g1196 ( 
.A(n_1047),
.B(n_1042),
.C(n_1008),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1069),
.A2(n_1002),
.B(n_1016),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1042),
.A2(n_998),
.B(n_1066),
.C(n_1054),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1056),
.B(n_1081),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_1056),
.B(n_1060),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1007),
.B(n_1081),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_1007),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1064),
.B(n_999),
.Y(n_1203)
);

O2A1O1Ixp5_ASAP7_75t_L g1204 ( 
.A1(n_1052),
.A2(n_1065),
.B(n_1032),
.C(n_1110),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_1021),
.Y(n_1205)
);

OR2x6_ASAP7_75t_L g1206 ( 
.A(n_1057),
.B(n_1021),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1060),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_1021),
.Y(n_1208)
);

NAND2x1_ASAP7_75t_L g1209 ( 
.A(n_1021),
.B(n_1081),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_1023),
.Y(n_1210)
);

INVx3_ASAP7_75t_SL g1211 ( 
.A(n_1023),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1063),
.A2(n_1005),
.B(n_1041),
.C(n_1003),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1073),
.A2(n_1001),
.B1(n_1048),
.B2(n_1034),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_1001),
.Y(n_1214)
);

BUFx2_ASAP7_75t_L g1215 ( 
.A(n_1001),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1001),
.B(n_1004),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_983),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1092),
.A2(n_1096),
.B(n_953),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1113),
.B(n_988),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1092),
.A2(n_1096),
.B(n_953),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_983),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_991),
.A2(n_1080),
.B(n_1069),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1224)
);

INVx4_ASAP7_75t_L g1225 ( 
.A(n_1078),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1039),
.Y(n_1226)
);

OR2x6_ASAP7_75t_L g1227 ( 
.A(n_1088),
.B(n_1038),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1004),
.B(n_1079),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_983),
.Y(n_1229)
);

OAI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_985),
.A2(n_953),
.B(n_1074),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1113),
.B(n_647),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1092),
.A2(n_1096),
.B(n_953),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_987),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_978),
.Y(n_1234)
);

OAI21xp33_ASAP7_75t_L g1235 ( 
.A1(n_1113),
.A2(n_953),
.B(n_1094),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1115),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_983),
.Y(n_1237)
);

OR2x2_ASAP7_75t_L g1238 ( 
.A(n_1115),
.B(n_1014),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_978),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1092),
.A2(n_1096),
.B(n_953),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_1078),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1092),
.A2(n_1096),
.B(n_953),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1113),
.A2(n_936),
.B(n_965),
.C(n_961),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_985),
.A2(n_953),
.B1(n_680),
.B2(n_1029),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_978),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_991),
.A2(n_1080),
.B(n_1069),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_987),
.Y(n_1247)
);

AND2x2_ASAP7_75t_SL g1248 ( 
.A(n_1011),
.B(n_456),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1113),
.B(n_988),
.Y(n_1250)
);

AO21x2_ASAP7_75t_L g1251 ( 
.A1(n_993),
.A2(n_976),
.B(n_964),
.Y(n_1251)
);

BUFx12f_ASAP7_75t_L g1252 ( 
.A(n_1089),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1013),
.B(n_1109),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_978),
.Y(n_1254)
);

AOI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1113),
.A2(n_662),
.B1(n_656),
.B2(n_953),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_1062),
.Y(n_1256)
);

A2O1A1Ixp33_ASAP7_75t_SL g1257 ( 
.A1(n_1092),
.A2(n_1096),
.B(n_1101),
.C(n_1094),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1115),
.B(n_1014),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_SL g1259 ( 
.A1(n_1092),
.A2(n_1096),
.B(n_1101),
.C(n_1094),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1078),
.Y(n_1260)
);

OR2x6_ASAP7_75t_L g1261 ( 
.A(n_1088),
.B(n_1038),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1248),
.A2(n_1231),
.B1(n_1230),
.B2(n_1150),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1255),
.A2(n_1154),
.B1(n_1235),
.B2(n_1128),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1132),
.B(n_1148),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_1161),
.Y(n_1265)
);

BUFx4f_ASAP7_75t_SL g1266 ( 
.A(n_1252),
.Y(n_1266)
);

BUFx8_ASAP7_75t_L g1267 ( 
.A(n_1131),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1123),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_SL g1269 ( 
.A1(n_1130),
.A2(n_1221),
.B(n_1218),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1141),
.B(n_1183),
.Y(n_1270)
);

INVx1_ASAP7_75t_SL g1271 ( 
.A(n_1228),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1137),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1143),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1145),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1147),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1149),
.B(n_1156),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1168),
.Y(n_1277)
);

INVx2_ASAP7_75t_SL g1278 ( 
.A(n_1127),
.Y(n_1278)
);

INVxp67_ASAP7_75t_L g1279 ( 
.A(n_1176),
.Y(n_1279)
);

CKINVDCx11_ASAP7_75t_R g1280 ( 
.A(n_1122),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1255),
.B(n_1128),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1235),
.A2(n_1158),
.B1(n_1160),
.B2(n_1135),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1160),
.A2(n_1135),
.B1(n_1150),
.B2(n_1152),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1210),
.Y(n_1284)
);

AOI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1166),
.A2(n_1159),
.B1(n_1250),
.B2(n_1220),
.Y(n_1285)
);

BUFx2_ASAP7_75t_R g1286 ( 
.A(n_1174),
.Y(n_1286)
);

OAI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1166),
.A2(n_1157),
.B1(n_1230),
.B2(n_1240),
.Y(n_1287)
);

OA21x2_ASAP7_75t_L g1288 ( 
.A1(n_1187),
.A2(n_1189),
.B(n_1212),
.Y(n_1288)
);

AO21x1_ASAP7_75t_L g1289 ( 
.A1(n_1232),
.A2(n_1242),
.B(n_1244),
.Y(n_1289)
);

AO21x1_ASAP7_75t_L g1290 ( 
.A1(n_1244),
.A2(n_1164),
.B(n_1167),
.Y(n_1290)
);

INVx4_ASAP7_75t_SL g1291 ( 
.A(n_1211),
.Y(n_1291)
);

HB1xp67_ASAP7_75t_L g1292 ( 
.A(n_1226),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1216),
.A2(n_1172),
.B1(n_1163),
.B2(n_1258),
.Y(n_1293)
);

OR2x6_ASAP7_75t_L g1294 ( 
.A(n_1141),
.B(n_1139),
.Y(n_1294)
);

BUFx2_ASAP7_75t_R g1295 ( 
.A(n_1125),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1217),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1222),
.Y(n_1297)
);

INVx1_ASAP7_75t_SL g1298 ( 
.A(n_1127),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1229),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1237),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1179),
.Y(n_1301)
);

INVx2_ASAP7_75t_SL g1302 ( 
.A(n_1134),
.Y(n_1302)
);

INVxp33_ASAP7_75t_L g1303 ( 
.A(n_1134),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_SL g1304 ( 
.A1(n_1162),
.A2(n_1146),
.B1(n_1236),
.B2(n_1238),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_SL g1305 ( 
.A1(n_1162),
.A2(n_1146),
.B1(n_1236),
.B2(n_1215),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1207),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1120),
.B(n_1181),
.Y(n_1307)
);

CKINVDCx6p67_ASAP7_75t_R g1308 ( 
.A(n_1122),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_1121),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1219),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1243),
.A2(n_1129),
.B1(n_1165),
.B2(n_1260),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1188),
.A2(n_1223),
.B(n_1246),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1165),
.A2(n_1249),
.B1(n_1253),
.B2(n_1224),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1249),
.A2(n_1253),
.B1(n_1254),
.B2(n_1185),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1200),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1193),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1153),
.B(n_1241),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1234),
.A2(n_1245),
.B1(n_1239),
.B2(n_1251),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1124),
.A2(n_1259),
.B(n_1257),
.Y(n_1319)
);

OA21x2_ASAP7_75t_L g1320 ( 
.A1(n_1187),
.A2(n_1204),
.B(n_1142),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1251),
.A2(n_1192),
.B1(n_1173),
.B2(n_1194),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1184),
.A2(n_1140),
.B1(n_1225),
.B2(n_1155),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1195),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1194),
.A2(n_1261),
.B1(n_1227),
.B2(n_1169),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1139),
.A2(n_1261),
.B1(n_1227),
.B2(n_1169),
.Y(n_1325)
);

INVx3_ASAP7_75t_SL g1326 ( 
.A(n_1153),
.Y(n_1326)
);

CKINVDCx12_ASAP7_75t_R g1327 ( 
.A(n_1139),
.Y(n_1327)
);

CKINVDCx20_ASAP7_75t_R g1328 ( 
.A(n_1133),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1155),
.B(n_1225),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1214),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1197),
.A2(n_1213),
.B(n_1198),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1138),
.B(n_1191),
.Y(n_1332)
);

INVx4_ASAP7_75t_L g1333 ( 
.A(n_1190),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1126),
.Y(n_1334)
);

BUFx6f_ASAP7_75t_L g1335 ( 
.A(n_1190),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_1175),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1203),
.Y(n_1337)
);

AOI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1261),
.A2(n_1170),
.B1(n_1180),
.B2(n_1183),
.Y(n_1338)
);

BUFx2_ASAP7_75t_R g1339 ( 
.A(n_1178),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1199),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1196),
.A2(n_1209),
.B(n_1201),
.Y(n_1341)
);

AOI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1206),
.A2(n_1205),
.B(n_1202),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1208),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_SL g1344 ( 
.A(n_1126),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1121),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_SL g1346 ( 
.A1(n_1177),
.A2(n_1206),
.B(n_1144),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1171),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1171),
.Y(n_1348)
);

OA21x2_ASAP7_75t_L g1349 ( 
.A1(n_1186),
.A2(n_1233),
.B(n_1247),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1233),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1247),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1247),
.A2(n_1136),
.B1(n_1144),
.B2(n_1256),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_SL g1353 ( 
.A1(n_1231),
.A2(n_1113),
.B1(n_1114),
.B2(n_662),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1125),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1226),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1231),
.A2(n_1113),
.B1(n_1248),
.B2(n_1255),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1231),
.A2(n_1113),
.B1(n_1248),
.B2(n_1255),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1210),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1226),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_1125),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1231),
.A2(n_1113),
.B1(n_1248),
.B2(n_1255),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1231),
.A2(n_1113),
.B1(n_1248),
.B2(n_1255),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1151),
.B(n_1131),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1255),
.A2(n_953),
.B1(n_1231),
.B2(n_1135),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1182),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_1210),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1231),
.A2(n_1113),
.B1(n_1248),
.B2(n_1255),
.Y(n_1367)
);

INVx2_ASAP7_75t_SL g1368 ( 
.A(n_1127),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_L g1369 ( 
.A(n_1335),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1323),
.B(n_1281),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1337),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1306),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1281),
.B(n_1268),
.Y(n_1373)
);

AND2x4_ASAP7_75t_SL g1374 ( 
.A(n_1294),
.B(n_1324),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1272),
.B(n_1273),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1285),
.B(n_1263),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1274),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1341),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1320),
.Y(n_1379)
);

OAI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1364),
.A2(n_1357),
.B(n_1356),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1275),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1320),
.Y(n_1382)
);

INVx3_ASAP7_75t_L g1383 ( 
.A(n_1341),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1279),
.B(n_1354),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1277),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1349),
.Y(n_1386)
);

BUFx4f_ASAP7_75t_SL g1387 ( 
.A(n_1328),
.Y(n_1387)
);

AO21x2_ASAP7_75t_L g1388 ( 
.A1(n_1332),
.A2(n_1319),
.B(n_1289),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1296),
.B(n_1297),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1299),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1300),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1315),
.B(n_1363),
.Y(n_1392)
);

OA21x2_ASAP7_75t_L g1393 ( 
.A1(n_1331),
.A2(n_1312),
.B(n_1290),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1320),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1288),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1292),
.B(n_1355),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1330),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1316),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1262),
.B(n_1359),
.Y(n_1399)
);

INVxp67_ASAP7_75t_L g1400 ( 
.A(n_1311),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_SL g1401 ( 
.A1(n_1287),
.A2(n_1294),
.B(n_1338),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1282),
.A2(n_1353),
.B1(n_1357),
.B2(n_1367),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1269),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1288),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1301),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1271),
.B(n_1263),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1321),
.A2(n_1283),
.B(n_1318),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1340),
.Y(n_1408)
);

AO21x1_ASAP7_75t_SL g1409 ( 
.A1(n_1283),
.A2(n_1282),
.B(n_1324),
.Y(n_1409)
);

AO21x2_ASAP7_75t_L g1410 ( 
.A1(n_1365),
.A2(n_1342),
.B(n_1346),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1307),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1321),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1270),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1356),
.B(n_1361),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1350),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1361),
.B(n_1367),
.Y(n_1416)
);

CKINVDCx14_ASAP7_75t_R g1417 ( 
.A(n_1328),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1345),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1347),
.Y(n_1419)
);

INVxp67_ASAP7_75t_SL g1420 ( 
.A(n_1362),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1348),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1309),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1293),
.B(n_1362),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1305),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1309),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1325),
.A2(n_1322),
.B(n_1313),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1276),
.B(n_1264),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1284),
.B(n_1366),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1291),
.B(n_1351),
.Y(n_1429)
);

INVxp67_ASAP7_75t_L g1430 ( 
.A(n_1343),
.Y(n_1430)
);

INVx4_ASAP7_75t_L g1431 ( 
.A(n_1369),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1370),
.B(n_1358),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1398),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1373),
.B(n_1304),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1373),
.B(n_1343),
.Y(n_1435)
);

INVx2_ASAP7_75t_R g1436 ( 
.A(n_1386),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1402),
.A2(n_1327),
.B1(n_1314),
.B2(n_1267),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1398),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1408),
.B(n_1352),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1396),
.B(n_1405),
.Y(n_1440)
);

INVxp67_ASAP7_75t_SL g1441 ( 
.A(n_1379),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1379),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1377),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1408),
.B(n_1267),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1381),
.Y(n_1445)
);

INVx5_ASAP7_75t_L g1446 ( 
.A(n_1395),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1397),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1381),
.Y(n_1448)
);

INVxp67_ASAP7_75t_SL g1449 ( 
.A(n_1382),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1382),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1385),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1387),
.B(n_1334),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1385),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1409),
.A2(n_1298),
.B1(n_1303),
.B2(n_1267),
.Y(n_1454)
);

INVxp67_ASAP7_75t_L g1455 ( 
.A(n_1410),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1404),
.B(n_1291),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1395),
.B(n_1291),
.Y(n_1457)
);

AOI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1414),
.A2(n_1368),
.B1(n_1302),
.B2(n_1278),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1395),
.B(n_1310),
.Y(n_1459)
);

BUFx2_ASAP7_75t_L g1460 ( 
.A(n_1422),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1422),
.Y(n_1461)
);

NAND3xp33_ASAP7_75t_L g1462 ( 
.A(n_1400),
.B(n_1334),
.C(n_1280),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1415),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1372),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1394),
.B(n_1329),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1393),
.B(n_1303),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1415),
.Y(n_1467)
);

BUFx2_ASAP7_75t_SL g1468 ( 
.A(n_1429),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1396),
.B(n_1336),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1371),
.B(n_1333),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1405),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1392),
.B(n_1317),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1375),
.B(n_1265),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_SL g1474 ( 
.A1(n_1434),
.A2(n_1420),
.B1(n_1414),
.B2(n_1416),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1465),
.B(n_1378),
.Y(n_1475)
);

OAI221xp5_ASAP7_75t_SL g1476 ( 
.A1(n_1437),
.A2(n_1400),
.B1(n_1420),
.B2(n_1376),
.C(n_1416),
.Y(n_1476)
);

NAND3xp33_ASAP7_75t_L g1477 ( 
.A(n_1455),
.B(n_1380),
.C(n_1376),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1433),
.B(n_1411),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1464),
.Y(n_1479)
);

NOR3xp33_ASAP7_75t_L g1480 ( 
.A(n_1462),
.B(n_1380),
.C(n_1403),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1433),
.B(n_1399),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1438),
.B(n_1399),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1438),
.B(n_1440),
.Y(n_1483)
);

OAI21xp33_ASAP7_75t_L g1484 ( 
.A1(n_1434),
.A2(n_1423),
.B(n_1424),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1437),
.A2(n_1423),
.B1(n_1417),
.B2(n_1430),
.Y(n_1485)
);

OAI221xp5_ASAP7_75t_SL g1486 ( 
.A1(n_1455),
.A2(n_1424),
.B1(n_1406),
.B2(n_1412),
.C(n_1401),
.Y(n_1486)
);

AOI21xp33_ASAP7_75t_L g1487 ( 
.A1(n_1439),
.A2(n_1388),
.B(n_1412),
.Y(n_1487)
);

NAND3xp33_ASAP7_75t_L g1488 ( 
.A(n_1439),
.B(n_1418),
.C(n_1371),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_SL g1489 ( 
.A(n_1444),
.B(n_1430),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1471),
.B(n_1389),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1471),
.B(n_1435),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1435),
.B(n_1389),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1465),
.B(n_1378),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1465),
.B(n_1388),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1432),
.B(n_1469),
.Y(n_1495)
);

NAND3xp33_ASAP7_75t_L g1496 ( 
.A(n_1442),
.B(n_1418),
.C(n_1419),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1432),
.B(n_1388),
.Y(n_1497)
);

NAND4xp25_ASAP7_75t_L g1498 ( 
.A(n_1462),
.B(n_1384),
.C(n_1428),
.D(n_1425),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1459),
.B(n_1383),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1444),
.A2(n_1428),
.B1(n_1401),
.B2(n_1374),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1469),
.B(n_1473),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1456),
.B(n_1383),
.Y(n_1502)
);

OAI21xp5_ASAP7_75t_SL g1503 ( 
.A1(n_1456),
.A2(n_1406),
.B(n_1429),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1473),
.B(n_1388),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1454),
.A2(n_1458),
.B1(n_1468),
.B2(n_1470),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1443),
.B(n_1427),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1463),
.B(n_1413),
.Y(n_1507)
);

NAND3xp33_ASAP7_75t_L g1508 ( 
.A(n_1442),
.B(n_1419),
.C(n_1421),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1443),
.B(n_1427),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1463),
.B(n_1413),
.Y(n_1510)
);

NAND4xp25_ASAP7_75t_L g1511 ( 
.A(n_1460),
.B(n_1425),
.C(n_1391),
.D(n_1390),
.Y(n_1511)
);

AOI211xp5_ASAP7_75t_L g1512 ( 
.A1(n_1441),
.A2(n_1426),
.B(n_1326),
.C(n_1391),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_SL g1513 ( 
.A1(n_1452),
.A2(n_1457),
.B(n_1458),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1472),
.B(n_1280),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_SL g1515 ( 
.A(n_1431),
.B(n_1295),
.Y(n_1515)
);

NOR3xp33_ASAP7_75t_SL g1516 ( 
.A(n_1470),
.B(n_1360),
.C(n_1354),
.Y(n_1516)
);

NAND3xp33_ASAP7_75t_L g1517 ( 
.A(n_1477),
.B(n_1450),
.C(n_1449),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1497),
.B(n_1450),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1475),
.B(n_1493),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1494),
.B(n_1441),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1475),
.B(n_1493),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1479),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1483),
.B(n_1449),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1508),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1490),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1504),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1496),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1478),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1477),
.B(n_1445),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_1499),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1502),
.B(n_1446),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1506),
.B(n_1445),
.Y(n_1532)
);

OA21x2_ASAP7_75t_L g1533 ( 
.A1(n_1487),
.A2(n_1466),
.B(n_1447),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1488),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1507),
.B(n_1436),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1509),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1489),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1512),
.B(n_1467),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1481),
.B(n_1460),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1510),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1491),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1495),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1482),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1498),
.B(n_1344),
.Y(n_1544)
);

AND2x4_ASAP7_75t_SL g1545 ( 
.A(n_1516),
.B(n_1457),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1492),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1503),
.B(n_1436),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1523),
.B(n_1501),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1524),
.B(n_1448),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1529),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1524),
.B(n_1448),
.Y(n_1551)
);

INVx2_ASAP7_75t_SL g1552 ( 
.A(n_1547),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1529),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1547),
.B(n_1514),
.Y(n_1554)
);

INVx1_ASAP7_75t_SL g1555 ( 
.A(n_1534),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1545),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1547),
.B(n_1446),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1534),
.B(n_1451),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1531),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1530),
.B(n_1489),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1522),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1530),
.B(n_1513),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1527),
.B(n_1451),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1522),
.Y(n_1564)
);

OR2x6_ASAP7_75t_L g1565 ( 
.A(n_1517),
.B(n_1426),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1519),
.B(n_1436),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1522),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1531),
.B(n_1446),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1519),
.B(n_1467),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1537),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1519),
.B(n_1521),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1523),
.B(n_1511),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1523),
.B(n_1461),
.Y(n_1573)
);

INVxp67_ASAP7_75t_L g1574 ( 
.A(n_1527),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1522),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1532),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1528),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1540),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1546),
.B(n_1453),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1536),
.B(n_1453),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1555),
.B(n_1528),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1570),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1555),
.B(n_1537),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1556),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1574),
.B(n_1536),
.Y(n_1585)
);

INVxp67_ASAP7_75t_SL g1586 ( 
.A(n_1574),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1549),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1571),
.B(n_1562),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1549),
.Y(n_1589)
);

OAI21xp33_ASAP7_75t_L g1590 ( 
.A1(n_1565),
.A2(n_1517),
.B(n_1538),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1571),
.B(n_1531),
.Y(n_1591)
);

AOI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1550),
.A2(n_1484),
.B1(n_1520),
.B2(n_1526),
.C(n_1544),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1562),
.B(n_1556),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1565),
.A2(n_1484),
.B1(n_1474),
.B2(n_1533),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1580),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1556),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1551),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1570),
.B(n_1542),
.Y(n_1598)
);

INVxp67_ASAP7_75t_SL g1599 ( 
.A(n_1577),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1580),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1561),
.Y(n_1601)
);

AOI31xp33_ASAP7_75t_L g1602 ( 
.A1(n_1577),
.A2(n_1544),
.A3(n_1538),
.B(n_1512),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1551),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1550),
.B(n_1542),
.Y(n_1604)
);

NAND4xp75_ASAP7_75t_L g1605 ( 
.A(n_1552),
.B(n_1533),
.C(n_1407),
.D(n_1535),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1548),
.B(n_1518),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1563),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1560),
.B(n_1531),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1563),
.Y(n_1609)
);

INVx3_ASAP7_75t_L g1610 ( 
.A(n_1568),
.Y(n_1610)
);

NAND4xp25_ASAP7_75t_L g1611 ( 
.A(n_1572),
.B(n_1480),
.C(n_1515),
.D(n_1539),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1554),
.B(n_1266),
.Y(n_1612)
);

NAND4xp25_ASAP7_75t_L g1613 ( 
.A(n_1572),
.B(n_1539),
.C(n_1541),
.D(n_1525),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1560),
.B(n_1531),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1553),
.B(n_1541),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1565),
.A2(n_1486),
.B(n_1476),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1548),
.B(n_1518),
.Y(n_1617)
);

INVx4_ASAP7_75t_L g1618 ( 
.A(n_1565),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1553),
.B(n_1543),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1558),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1558),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1559),
.B(n_1545),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1579),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1605),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1623),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1588),
.B(n_1554),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1586),
.Y(n_1627)
);

INVx1_ASAP7_75t_SL g1628 ( 
.A(n_1593),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1588),
.B(n_1559),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1623),
.Y(n_1630)
);

NOR2x1_ASAP7_75t_L g1631 ( 
.A(n_1618),
.B(n_1605),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1593),
.Y(n_1632)
);

INVx1_ASAP7_75t_SL g1633 ( 
.A(n_1582),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1618),
.B(n_1565),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1606),
.B(n_1576),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1606),
.B(n_1617),
.Y(n_1636)
);

OAI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1602),
.A2(n_1565),
.B1(n_1552),
.B2(n_1545),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1612),
.B(n_1266),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1604),
.Y(n_1639)
);

OAI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1594),
.A2(n_1618),
.B1(n_1616),
.B2(n_1590),
.Y(n_1640)
);

INVx2_ASAP7_75t_SL g1641 ( 
.A(n_1584),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1601),
.Y(n_1642)
);

INVx3_ASAP7_75t_L g1643 ( 
.A(n_1622),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1601),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1583),
.B(n_1581),
.Y(n_1645)
);

OR2x6_ASAP7_75t_L g1646 ( 
.A(n_1596),
.B(n_1552),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1592),
.A2(n_1533),
.B1(n_1407),
.B2(n_1485),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1617),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1619),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1584),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1615),
.Y(n_1651)
);

AOI22x1_ASAP7_75t_L g1652 ( 
.A1(n_1599),
.A2(n_1559),
.B1(n_1360),
.B2(n_1557),
.Y(n_1652)
);

INVxp67_ASAP7_75t_L g1653 ( 
.A(n_1596),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1622),
.B(n_1559),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1585),
.B(n_1576),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1595),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1598),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1595),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1622),
.B(n_1566),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1628),
.B(n_1620),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1624),
.A2(n_1611),
.B1(n_1613),
.B2(n_1533),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1632),
.B(n_1621),
.Y(n_1662)
);

OAI22xp5_ASAP7_75t_SL g1663 ( 
.A1(n_1627),
.A2(n_1584),
.B1(n_1326),
.B2(n_1557),
.Y(n_1663)
);

INVx4_ASAP7_75t_L g1664 ( 
.A(n_1627),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1636),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1648),
.B(n_1587),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1636),
.Y(n_1667)
);

OAI21xp33_ASAP7_75t_SL g1668 ( 
.A1(n_1631),
.A2(n_1614),
.B(n_1608),
.Y(n_1668)
);

AOI221x1_ASAP7_75t_L g1669 ( 
.A1(n_1640),
.A2(n_1610),
.B1(n_1589),
.B2(n_1603),
.C(n_1609),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1624),
.A2(n_1610),
.B1(n_1591),
.B2(n_1614),
.Y(n_1670)
);

INVxp67_ASAP7_75t_L g1671 ( 
.A(n_1650),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1648),
.B(n_1597),
.Y(n_1672)
);

AND2x4_ASAP7_75t_SL g1673 ( 
.A(n_1638),
.B(n_1308),
.Y(n_1673)
);

AOI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1624),
.A2(n_1533),
.B1(n_1607),
.B2(n_1500),
.Y(n_1674)
);

AOI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1631),
.A2(n_1533),
.B1(n_1600),
.B2(n_1566),
.Y(n_1675)
);

INVxp67_ASAP7_75t_SL g1676 ( 
.A(n_1653),
.Y(n_1676)
);

OAI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1637),
.A2(n_1610),
.B1(n_1520),
.B2(n_1505),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1648),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1633),
.B(n_1600),
.Y(n_1679)
);

AOI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1647),
.A2(n_1566),
.B1(n_1557),
.B2(n_1535),
.Y(n_1680)
);

BUFx3_ASAP7_75t_L g1681 ( 
.A(n_1650),
.Y(n_1681)
);

AOI21xp33_ASAP7_75t_SL g1682 ( 
.A1(n_1652),
.A2(n_1557),
.B(n_1608),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1625),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1625),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1630),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1664),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1664),
.B(n_1676),
.Y(n_1687)
);

NOR2x1_ASAP7_75t_L g1688 ( 
.A(n_1681),
.B(n_1643),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1665),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1667),
.B(n_1626),
.Y(n_1690)
);

INVx2_ASAP7_75t_SL g1691 ( 
.A(n_1673),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1670),
.B(n_1626),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1668),
.B(n_1643),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1678),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1671),
.B(n_1657),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1669),
.B(n_1639),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1683),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1666),
.B(n_1639),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1684),
.Y(n_1699)
);

INVx1_ASAP7_75t_SL g1700 ( 
.A(n_1679),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1668),
.B(n_1643),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1661),
.B(n_1643),
.Y(n_1702)
);

NOR2x1_ASAP7_75t_L g1703 ( 
.A(n_1685),
.B(n_1646),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_L g1704 ( 
.A(n_1660),
.B(n_1641),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1672),
.B(n_1649),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_SL g1706 ( 
.A(n_1693),
.B(n_1675),
.Y(n_1706)
);

NAND3xp33_ASAP7_75t_L g1707 ( 
.A(n_1696),
.B(n_1701),
.C(n_1693),
.Y(n_1707)
);

AOI211xp5_ASAP7_75t_L g1708 ( 
.A1(n_1701),
.A2(n_1677),
.B(n_1663),
.C(n_1634),
.Y(n_1708)
);

AOI211xp5_ASAP7_75t_SL g1709 ( 
.A1(n_1687),
.A2(n_1662),
.B(n_1634),
.C(n_1680),
.Y(n_1709)
);

OAI21xp33_ASAP7_75t_L g1710 ( 
.A1(n_1702),
.A2(n_1645),
.B(n_1674),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_SL g1711 ( 
.A1(n_1702),
.A2(n_1634),
.B1(n_1652),
.B2(n_1651),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_L g1712 ( 
.A(n_1691),
.B(n_1700),
.Y(n_1712)
);

AOI221xp5_ASAP7_75t_L g1713 ( 
.A1(n_1694),
.A2(n_1634),
.B1(n_1649),
.B2(n_1651),
.C(n_1630),
.Y(n_1713)
);

AOI221xp5_ASAP7_75t_L g1714 ( 
.A1(n_1705),
.A2(n_1658),
.B1(n_1656),
.B2(n_1655),
.C(n_1642),
.Y(n_1714)
);

AOI222xp33_ASAP7_75t_L g1715 ( 
.A1(n_1689),
.A2(n_1642),
.B1(n_1644),
.B2(n_1658),
.C1(n_1656),
.C2(n_1641),
.Y(n_1715)
);

AOI222xp33_ASAP7_75t_L g1716 ( 
.A1(n_1698),
.A2(n_1642),
.B1(n_1644),
.B2(n_1629),
.C1(n_1659),
.C2(n_1564),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1690),
.A2(n_1682),
.B1(n_1646),
.B2(n_1635),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1712),
.Y(n_1718)
);

AOI211xp5_ASAP7_75t_L g1719 ( 
.A1(n_1706),
.A2(n_1704),
.B(n_1692),
.C(n_1695),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1715),
.Y(n_1720)
);

AOI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1710),
.A2(n_1704),
.B1(n_1703),
.B2(n_1688),
.Y(n_1721)
);

NOR2x1_ASAP7_75t_L g1722 ( 
.A(n_1707),
.B(n_1686),
.Y(n_1722)
);

NOR2x1_ASAP7_75t_L g1723 ( 
.A(n_1717),
.B(n_1686),
.Y(n_1723)
);

NOR3x1_ASAP7_75t_L g1724 ( 
.A(n_1709),
.B(n_1691),
.C(n_1697),
.Y(n_1724)
);

NAND5xp2_ASAP7_75t_L g1725 ( 
.A(n_1708),
.B(n_1711),
.C(n_1716),
.D(n_1713),
.E(n_1714),
.Y(n_1725)
);

NAND4xp75_ASAP7_75t_L g1726 ( 
.A(n_1706),
.B(n_1699),
.C(n_1659),
.D(n_1629),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1712),
.Y(n_1727)
);

XNOR2x1_ASAP7_75t_SL g1728 ( 
.A(n_1712),
.B(n_1654),
.Y(n_1728)
);

NOR2x1_ASAP7_75t_L g1729 ( 
.A(n_1707),
.B(n_1699),
.Y(n_1729)
);

NOR3xp33_ASAP7_75t_L g1730 ( 
.A(n_1718),
.B(n_1635),
.C(n_1654),
.Y(n_1730)
);

O2A1O1Ixp33_ASAP7_75t_SL g1731 ( 
.A1(n_1725),
.A2(n_1573),
.B(n_1646),
.C(n_1286),
.Y(n_1731)
);

AOI211xp5_ASAP7_75t_L g1732 ( 
.A1(n_1720),
.A2(n_1568),
.B(n_1591),
.C(n_1646),
.Y(n_1732)
);

NOR3xp33_ASAP7_75t_SL g1733 ( 
.A(n_1726),
.B(n_1344),
.C(n_1646),
.Y(n_1733)
);

AOI22xp5_ASAP7_75t_L g1734 ( 
.A1(n_1729),
.A2(n_1564),
.B1(n_1561),
.B2(n_1578),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1727),
.B(n_1721),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1728),
.B(n_1569),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1735),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1736),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1730),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1734),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1732),
.Y(n_1741)
);

AOI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1731),
.A2(n_1722),
.B1(n_1719),
.B2(n_1723),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1737),
.Y(n_1743)
);

BUFx2_ASAP7_75t_L g1744 ( 
.A(n_1738),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1740),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1739),
.Y(n_1746)
);

NAND3xp33_ASAP7_75t_L g1747 ( 
.A(n_1742),
.B(n_1733),
.C(n_1724),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1743),
.Y(n_1748)
);

XNOR2x1_ASAP7_75t_L g1749 ( 
.A(n_1745),
.B(n_1742),
.Y(n_1749)
);

AND2x2_ASAP7_75t_SL g1750 ( 
.A(n_1744),
.B(n_1741),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1750),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1751),
.Y(n_1752)
);

OAI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1752),
.A2(n_1748),
.B1(n_1747),
.B2(n_1749),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1752),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1754),
.Y(n_1755)
);

XNOR2xp5_ASAP7_75t_L g1756 ( 
.A(n_1753),
.B(n_1747),
.Y(n_1756)
);

INVxp67_ASAP7_75t_SL g1757 ( 
.A(n_1756),
.Y(n_1757)
);

OAI21xp5_ASAP7_75t_SL g1758 ( 
.A1(n_1755),
.A2(n_1748),
.B(n_1746),
.Y(n_1758)
);

OAI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1758),
.A2(n_1578),
.B(n_1564),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1759),
.Y(n_1760)
);

AOI221xp5_ASAP7_75t_L g1761 ( 
.A1(n_1760),
.A2(n_1757),
.B1(n_1561),
.B2(n_1567),
.C(n_1575),
.Y(n_1761)
);

AOI211xp5_ASAP7_75t_L g1762 ( 
.A1(n_1761),
.A2(n_1339),
.B(n_1568),
.C(n_1575),
.Y(n_1762)
);


endmodule