module fake_jpeg_16135_n_272 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_31;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_40),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_38),
.Y(n_60)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_47),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_30),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_30),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_22),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_30),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_48),
.A2(n_54),
.B(n_47),
.C(n_49),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_22),
.Y(n_49)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_28),
.Y(n_54)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_16),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_21),
.B1(n_18),
.B2(n_25),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_19),
.B1(n_23),
.B2(n_28),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_45),
.A2(n_21),
.B1(n_25),
.B2(n_18),
.Y(n_63)
);

OAI32xp33_ASAP7_75t_L g100 ( 
.A1(n_63),
.A2(n_74),
.A3(n_80),
.B1(n_83),
.B2(n_27),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_68),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_21),
.B1(n_25),
.B2(n_18),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_65),
.B(n_71),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_18),
.B1(n_60),
.B2(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_73),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_43),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_44),
.A2(n_42),
.B1(n_38),
.B2(n_34),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_42),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_87),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_38),
.B1(n_34),
.B2(n_23),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_50),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_56),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_67),
.C(n_71),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_33),
.B1(n_32),
.B2(n_17),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_51),
.A2(n_23),
.B1(n_19),
.B2(n_28),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_82),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_60),
.A2(n_33),
.B1(n_32),
.B2(n_17),
.Y(n_83)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_81),
.Y(n_89)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_46),
.C(n_56),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_104),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_101),
.Y(n_128)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_27),
.B1(n_20),
.B2(n_29),
.Y(n_136)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_105),
.Y(n_131)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_77),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_110),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_64),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_108),
.A2(n_86),
.B1(n_87),
.B2(n_48),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_48),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_111),
.Y(n_113)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_73),
.C(n_86),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_103),
.B(n_84),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_120),
.B(n_124),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_100),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_117),
.A2(n_75),
.B(n_13),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_63),
.B1(n_50),
.B2(n_51),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_50),
.B1(n_51),
.B2(n_66),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_122),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_66),
.B1(n_65),
.B2(n_57),
.Y(n_123)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_66),
.B1(n_57),
.B2(n_52),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_102),
.Y(n_125)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_53),
.B1(n_79),
.B2(n_15),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_127),
.A2(n_133),
.B(n_106),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_101),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_132),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_90),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_53),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_95),
.A2(n_14),
.B1(n_11),
.B2(n_13),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_134),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_137),
.Y(n_146)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_56),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_138),
.B(n_16),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_111),
.B(n_104),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_139),
.A2(n_162),
.B1(n_137),
.B2(n_119),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_118),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_153),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_92),
.C(n_109),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_145),
.C(n_147),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_143),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_155),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_93),
.C(n_108),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_108),
.C(n_56),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_88),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_158),
.Y(n_168)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_77),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_134),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_156),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_75),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_77),
.Y(n_156)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_75),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_163),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_130),
.A2(n_89),
.B1(n_26),
.B2(n_29),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_129),
.B(n_0),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_134),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_99),
.Y(n_183)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_148),
.A2(n_115),
.B1(n_113),
.B2(n_135),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_173),
.B1(n_186),
.B2(n_189),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_159),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_170),
.B(n_179),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_171),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_115),
.Y(n_172)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_113),
.B1(n_120),
.B2(n_123),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_114),
.Y(n_174)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_165),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_184),
.Y(n_201)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_160),
.A2(n_114),
.B1(n_124),
.B2(n_127),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_143),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_187),
.B(n_140),
.Y(n_194)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_141),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_162),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_146),
.A2(n_133),
.B1(n_89),
.B2(n_134),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_188),
.A2(n_141),
.B(n_155),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_192),
.A2(n_206),
.B(n_184),
.Y(n_218)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_142),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_169),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_167),
.A2(n_144),
.B1(n_145),
.B2(n_152),
.Y(n_196)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

XNOR2x1_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_158),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_198),
.B(n_189),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_147),
.C(n_139),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_204),
.C(n_205),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_L g202 ( 
.A1(n_167),
.A2(n_161),
.B(n_163),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_202),
.A2(n_207),
.B(n_175),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_164),
.C(n_154),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_150),
.C(n_61),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_174),
.A2(n_150),
.B(n_11),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_61),
.C(n_37),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_209),
.C(n_170),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_31),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_210),
.A2(n_218),
.B1(n_200),
.B2(n_191),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_180),
.Y(n_213)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_220),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_172),
.C(n_169),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_217),
.C(n_219),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_177),
.Y(n_216)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_173),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_182),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_181),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_222),
.C(n_223),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_177),
.C(n_186),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_196),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_192),
.C(n_206),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_229),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_203),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_232),
.C(n_234),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_197),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_236),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_224),
.A2(n_190),
.B1(n_191),
.B2(n_176),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_214),
.B(n_201),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_29),
.C(n_26),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_233),
.A2(n_231),
.B1(n_190),
.B2(n_201),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_238),
.A2(n_243),
.B1(n_244),
.B2(n_9),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_232),
.A2(n_176),
.B(n_211),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_240),
.A2(n_1),
.B(n_2),
.Y(n_252)
);

NOR3xp33_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_211),
.C(n_209),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_247),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_223),
.B1(n_219),
.B2(n_221),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_217),
.B1(n_10),
.B2(n_12),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_246),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_26),
.C(n_31),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_248),
.A2(n_249),
.B(n_252),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_226),
.B(n_228),
.Y(n_249)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_239),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_255),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_8),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_253),
.Y(n_261)
);

AOI221xp5_ASAP7_75t_L g257 ( 
.A1(n_254),
.A2(n_238),
.B1(n_9),
.B2(n_10),
.C(n_5),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_9),
.Y(n_255)
);

INVx11_ASAP7_75t_L g256 ( 
.A(n_251),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_260),
.Y(n_263)
);

AOI31xp67_ASAP7_75t_L g264 ( 
.A1(n_257),
.A2(n_7),
.A3(n_14),
.B(n_12),
.Y(n_264)
);

AOI322xp5_ASAP7_75t_L g260 ( 
.A1(n_248),
.A2(n_7),
.A3(n_14),
.B1(n_12),
.B2(n_6),
.C1(n_31),
.C2(n_24),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_7),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_259),
.C(n_24),
.Y(n_267)
);

NOR3xp33_ASAP7_75t_L g266 ( 
.A(n_264),
.B(n_260),
.C(n_2),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_6),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_1),
.Y(n_268)
);

AOI321xp33_ASAP7_75t_L g269 ( 
.A1(n_266),
.A2(n_267),
.A3(n_268),
.B1(n_1),
.B2(n_2),
.C(n_3),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_269),
.B(n_263),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_2),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_3),
.Y(n_272)
);


endmodule