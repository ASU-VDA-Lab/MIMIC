module fake_jpeg_4261_n_71 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_71);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_71;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_24;
wire n_26;
wire n_38;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_43;
wire n_37;
wire n_50;
wire n_29;
wire n_32;
wire n_70;
wire n_66;

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_5),
.B(n_18),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_11),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

AO22x1_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_21),
.B1(n_16),
.B2(n_14),
.Y(n_40)
);

A2O1A1O1Ixp25_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_49),
.B(n_51),
.C(n_26),
.D(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_42),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_28),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_1),
.C(n_2),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_47),
.C(n_50),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_2),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_52),
.B1(n_26),
.B2(n_36),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_24),
.A2(n_9),
.B(n_12),
.C(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_32),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_39),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_33),
.A2(n_38),
.B1(n_37),
.B2(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_55),
.Y(n_61)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_40),
.B1(n_44),
.B2(n_51),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_62),
.A2(n_57),
.B1(n_40),
.B2(n_59),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_58),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

BUFx4f_ASAP7_75t_SL g67 ( 
.A(n_66),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_68),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_60),
.C(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_69),
.B(n_65),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_53),
.B(n_46),
.Y(n_71)
);


endmodule