module fake_jpeg_31141_n_554 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_554);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_554;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

INVx11_ASAP7_75t_SL g39 ( 
.A(n_6),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_54),
.Y(n_139)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

NOR3xp33_ASAP7_75t_L g56 ( 
.A(n_23),
.B(n_10),
.C(n_16),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_56),
.A2(n_25),
.B1(n_42),
.B2(n_31),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_57),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_58),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_59),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

BUFx24_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVxp67_ASAP7_75t_SL g144 ( 
.A(n_61),
.Y(n_144)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g131 ( 
.A(n_63),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_64),
.Y(n_172)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_67),
.Y(n_162)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_69),
.Y(n_149)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_70),
.Y(n_111)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_73),
.Y(n_159)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_18),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_77),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_81),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_18),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_100),
.Y(n_127)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_88),
.Y(n_152)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_91),
.Y(n_160)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_23),
.B(n_38),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_107),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_94),
.Y(n_161)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_95),
.Y(n_157)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_96),
.Y(n_168)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_97),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_98),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_99),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_39),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_101),
.Y(n_177)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

CKINVDCx6p67_ASAP7_75t_R g118 ( 
.A(n_103),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_24),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_105),
.Y(n_135)
);

BUFx8_ASAP7_75t_L g105 ( 
.A(n_24),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_106),
.B(n_108),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_24),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_109),
.B(n_110),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_28),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_67),
.A2(n_24),
.B1(n_45),
.B2(n_49),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_115),
.A2(n_163),
.B1(n_167),
.B2(n_82),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_38),
.B1(n_50),
.B2(n_26),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_124),
.A2(n_130),
.B1(n_155),
.B2(n_156),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_126),
.B(n_145),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_84),
.A2(n_20),
.B1(n_49),
.B2(n_25),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_56),
.B(n_50),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_140),
.B(n_146),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_55),
.A2(n_26),
.B1(n_51),
.B2(n_44),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_77),
.B(n_31),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_53),
.A2(n_20),
.B1(n_49),
.B2(n_45),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_147),
.A2(n_64),
.B1(n_66),
.B2(n_73),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_86),
.A2(n_94),
.B1(n_99),
.B2(n_58),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_54),
.A2(n_51),
.B1(n_32),
.B2(n_44),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_59),
.A2(n_45),
.B1(n_20),
.B2(n_42),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_60),
.A2(n_43),
.B1(n_36),
.B2(n_32),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_165),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_63),
.A2(n_45),
.B1(n_43),
.B2(n_36),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_81),
.B(n_45),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_170),
.B(n_13),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_76),
.B(n_37),
.C(n_10),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_107),
.C(n_103),
.Y(n_187)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_172),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_178),
.Y(n_282)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_179),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_180),
.B(n_187),
.Y(n_258)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_181),
.Y(n_251)
);

BUFx12f_ASAP7_75t_L g182 ( 
.A(n_118),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g243 ( 
.A(n_182),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_184),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_127),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_185),
.B(n_186),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_128),
.B(n_79),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_121),
.B(n_105),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_188),
.Y(n_252)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_189),
.Y(n_245)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_190),
.Y(n_248)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_191),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_192),
.Y(n_253)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_193),
.Y(n_274)
);

BUFx8_ASAP7_75t_L g194 ( 
.A(n_112),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_194),
.Y(n_254)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_195),
.Y(n_247)
);

AND2x2_ASAP7_75t_SL g196 ( 
.A(n_113),
.B(n_101),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_196),
.B(n_221),
.C(n_3),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_118),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_197),
.B(n_213),
.Y(n_260)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_122),
.Y(n_198)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_198),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_135),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_199),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_200),
.A2(n_238),
.B1(n_143),
.B2(n_144),
.Y(n_269)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_129),
.Y(n_201)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_201),
.Y(n_285)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_132),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_202),
.Y(n_281)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_203),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_157),
.B(n_37),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_204),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_136),
.A2(n_80),
.B1(n_78),
.B2(n_61),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_206),
.A2(n_211),
.B1(n_224),
.B2(n_227),
.Y(n_262)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_151),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_207),
.B(n_209),
.Y(n_279)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_208),
.Y(n_263)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_151),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_126),
.A2(n_10),
.B(n_17),
.C(n_16),
.Y(n_210)
);

NAND4xp25_ASAP7_75t_L g273 ( 
.A(n_210),
.B(n_219),
.C(n_228),
.D(n_239),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_167),
.A2(n_37),
.B1(n_9),
.B2(n_11),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_158),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_212),
.Y(n_286)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_166),
.B(n_37),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_214),
.B(n_218),
.Y(n_255)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_215),
.B(n_216),
.Y(n_267)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_138),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

BUFx12_ASAP7_75t_L g259 ( 
.A(n_217),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_126),
.B(n_37),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_133),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_168),
.B(n_0),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_222),
.A2(n_223),
.B1(n_225),
.B2(n_226),
.Y(n_272)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_161),
.Y(n_223)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_134),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_119),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_131),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_227)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_133),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_163),
.A2(n_6),
.B1(n_14),
.B2(n_13),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_229),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_277)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_123),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_234),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_130),
.B(n_6),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_131),
.A2(n_6),
.B1(n_13),
.B2(n_12),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_125),
.B(n_5),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_125),
.B(n_5),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_138),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_235),
.B(n_237),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_155),
.A2(n_17),
.B1(n_5),
.B2(n_11),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_236),
.A2(n_115),
.B1(n_169),
.B2(n_154),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_111),
.B(n_11),
.Y(n_237)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_117),
.Y(n_239)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_117),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_159),
.B1(n_114),
.B2(n_172),
.Y(n_246)
);

AND2x2_ASAP7_75t_SL g244 ( 
.A(n_205),
.B(n_173),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_244),
.B(n_256),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_246),
.Y(n_320)
);

OA22x2_ASAP7_75t_L g249 ( 
.A1(n_183),
.A2(n_116),
.B1(n_119),
.B2(n_148),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_249),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_220),
.A2(n_111),
.B(n_112),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_250),
.A2(n_182),
.B(n_194),
.Y(n_317)
);

AND2x2_ASAP7_75t_SL g256 ( 
.A(n_221),
.B(n_149),
.Y(n_256)
);

OA22x2_ASAP7_75t_L g257 ( 
.A1(n_183),
.A2(n_116),
.B1(n_148),
.B2(n_147),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_257),
.A2(n_278),
.B1(n_182),
.B2(n_192),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_266),
.A2(n_268),
.B1(n_271),
.B2(n_275),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_217),
.A2(n_153),
.B1(n_141),
.B2(n_169),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_269),
.A2(n_196),
.B1(n_197),
.B2(n_213),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_236),
.A2(n_154),
.B1(n_139),
.B2(n_2),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_224),
.A2(n_139),
.B1(n_1),
.B2(n_3),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_180),
.A2(n_144),
.B1(n_11),
.B2(n_12),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_280),
.B(n_221),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_220),
.A2(n_0),
.B1(n_1),
.B2(n_187),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_287),
.A2(n_201),
.B1(n_202),
.B2(n_184),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_289),
.B(n_323),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_199),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_291),
.Y(n_333)
);

BUFx24_ASAP7_75t_SL g292 ( 
.A(n_252),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_292),
.B(n_295),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_220),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_293),
.B(n_294),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_198),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_281),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_241),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_296),
.B(n_298),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_241),
.B(n_189),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_299),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_270),
.A2(n_240),
.B1(n_239),
.B2(n_228),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_300),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_270),
.A2(n_178),
.B1(n_216),
.B2(n_179),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_301),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_276),
.B(n_210),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_302),
.B(n_303),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_191),
.Y(n_303)
);

INVx3_ASAP7_75t_SL g304 ( 
.A(n_282),
.Y(n_304)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_304),
.Y(n_340)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_285),
.Y(n_305)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_305),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_276),
.B(n_196),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_306),
.B(n_309),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_307),
.A2(n_321),
.B1(n_328),
.B2(n_266),
.Y(n_334)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_248),
.Y(n_308)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_308),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_252),
.B(n_279),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_310),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_258),
.B(n_244),
.C(n_264),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_311),
.B(n_319),
.C(n_256),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_281),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_312),
.B(n_314),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_288),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_248),
.Y(n_315)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_315),
.Y(n_349)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_274),
.Y(n_316)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_316),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_317),
.A2(n_260),
.B(n_267),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_258),
.B(n_193),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_318),
.B(n_322),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_258),
.B(n_244),
.C(n_255),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_280),
.B(n_225),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_255),
.B(n_223),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_257),
.A2(n_249),
.B1(n_262),
.B2(n_250),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_324),
.A2(n_249),
.B1(n_257),
.B2(n_273),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_273),
.A2(n_181),
.B1(n_226),
.B2(n_195),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_325),
.A2(n_272),
.B1(n_254),
.B2(n_260),
.Y(n_352)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_263),
.Y(n_326)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_326),
.Y(n_353)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_274),
.Y(n_327)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_327),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_269),
.A2(n_203),
.B1(n_194),
.B2(n_1),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_331),
.A2(n_320),
.B1(n_257),
.B2(n_275),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_334),
.A2(n_324),
.B1(n_290),
.B2(n_297),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_335),
.B(n_339),
.C(n_360),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_336),
.A2(n_347),
.B(n_361),
.Y(n_383)
);

NAND3xp33_ASAP7_75t_L g337 ( 
.A(n_302),
.B(n_310),
.C(n_306),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_337),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_277),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_317),
.A2(n_260),
.B(n_279),
.Y(n_347)
);

NAND2x1p5_ASAP7_75t_L g348 ( 
.A(n_313),
.B(n_256),
.Y(n_348)
);

AO22x1_ASAP7_75t_L g370 ( 
.A1(n_348),
.A2(n_313),
.B1(n_289),
.B2(n_322),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_304),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_351),
.B(n_253),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_352),
.A2(n_297),
.B1(n_321),
.B2(n_271),
.Y(n_365)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_308),
.Y(n_357)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_357),
.Y(n_376)
);

MAJx2_ASAP7_75t_L g359 ( 
.A(n_319),
.B(n_267),
.C(n_259),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_359),
.B(n_259),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_311),
.B(n_267),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_307),
.A2(n_328),
.B(n_318),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_293),
.A2(n_286),
.B(n_249),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_363),
.A2(n_305),
.B(n_251),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_364),
.A2(n_366),
.B1(n_368),
.B2(n_242),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_365),
.A2(n_374),
.B1(n_382),
.B2(n_395),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_334),
.A2(n_290),
.B1(n_363),
.B2(n_358),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_329),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_367),
.B(n_372),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_358),
.A2(n_296),
.B1(n_298),
.B2(n_303),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_370),
.B(n_353),
.Y(n_414)
);

CKINVDCx14_ASAP7_75t_R g371 ( 
.A(n_329),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_371),
.B(n_386),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_347),
.Y(n_372)
);

XNOR2x2_ASAP7_75t_SL g373 ( 
.A(n_346),
.B(n_323),
.Y(n_373)
);

AO22x1_ASAP7_75t_L g402 ( 
.A1(n_373),
.A2(n_362),
.B1(n_348),
.B2(n_360),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_331),
.A2(n_325),
.B1(n_304),
.B2(n_315),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_375),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_351),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_377),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_342),
.B(n_294),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_379),
.Y(n_428)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_380),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_342),
.B(n_286),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_381),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_361),
.A2(n_352),
.B1(n_333),
.B2(n_354),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_345),
.B(n_291),
.Y(n_384)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_384),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_335),
.B(n_309),
.C(n_299),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_385),
.B(n_348),
.C(n_330),
.Y(n_403)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_344),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_344),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_387),
.B(n_392),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_343),
.B(n_332),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_388),
.B(n_391),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_389),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_390),
.B(n_327),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_332),
.B(n_259),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_349),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_350),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_393),
.B(n_243),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_336),
.A2(n_346),
.B(n_354),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_394),
.A2(n_245),
.B(n_261),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_338),
.A2(n_300),
.B1(n_295),
.B2(n_312),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_356),
.A2(n_301),
.B(n_251),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_396),
.A2(n_340),
.B(n_355),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_382),
.A2(n_345),
.B1(n_339),
.B2(n_359),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_398),
.B(n_399),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_365),
.A2(n_359),
.B1(n_362),
.B2(n_357),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_374),
.A2(n_349),
.B1(n_330),
.B2(n_341),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_401),
.B(n_407),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_402),
.B(n_410),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_403),
.B(n_418),
.C(n_385),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_375),
.A2(n_341),
.B1(n_340),
.B2(n_351),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_408),
.A2(n_422),
.B(n_395),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_383),
.A2(n_355),
.B1(n_350),
.B2(n_353),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_412),
.B(n_414),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_371),
.A2(n_314),
.B1(n_282),
.B2(n_242),
.Y(n_415)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_415),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_416),
.B(n_421),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_381),
.B(n_254),
.Y(n_417)
);

CKINVDCx14_ASAP7_75t_R g435 ( 
.A(n_417),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_378),
.B(n_316),
.C(n_247),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_378),
.B(n_390),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_419),
.B(n_383),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_367),
.A2(n_253),
.B1(n_326),
.B2(n_247),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_420),
.Y(n_441)
);

NAND3xp33_ASAP7_75t_L g421 ( 
.A(n_369),
.B(n_261),
.C(n_284),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_396),
.A2(n_243),
.B(n_284),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_423),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_427),
.B(n_379),
.Y(n_447)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_425),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_430),
.B(n_438),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_431),
.B(n_434),
.C(n_436),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_433),
.B(n_447),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_370),
.C(n_394),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_419),
.B(n_370),
.C(n_391),
.Y(n_436)
);

BUFx12f_ASAP7_75t_SL g437 ( 
.A(n_417),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_437),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_409),
.B(n_388),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_409),
.B(n_411),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_439),
.B(n_445),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_403),
.B(n_370),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_442),
.B(n_448),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_405),
.B(n_389),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_446),
.B(n_454),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_398),
.B(n_384),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_412),
.B(n_399),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_449),
.B(n_451),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_426),
.A2(n_396),
.B(n_373),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_450),
.B(n_452),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_414),
.B(n_366),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_405),
.B(n_364),
.Y(n_452)
);

INVx13_ASAP7_75t_L g454 ( 
.A(n_423),
.Y(n_454)
);

MAJx2_ASAP7_75t_L g455 ( 
.A(n_402),
.B(n_373),
.C(n_368),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_455),
.B(n_402),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_432),
.A2(n_416),
.B1(n_404),
.B2(n_424),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_457),
.B(n_479),
.Y(n_490)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_437),
.Y(n_462)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_462),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_452),
.A2(n_397),
.B1(n_407),
.B2(n_410),
.Y(n_463)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_463),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_466),
.B(n_458),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_433),
.B(n_397),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_467),
.B(n_470),
.C(n_472),
.Y(n_482)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_447),
.Y(n_468)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_468),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_431),
.B(n_427),
.C(n_428),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_452),
.A2(n_401),
.B1(n_428),
.B2(n_411),
.Y(n_471)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_471),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_434),
.B(n_406),
.C(n_400),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_445),
.A2(n_441),
.B1(n_443),
.B2(n_435),
.Y(n_473)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_473),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_449),
.B(n_406),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_474),
.B(n_475),
.C(n_477),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_436),
.B(n_424),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_442),
.B(n_400),
.C(n_408),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_453),
.B(n_393),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_467),
.A2(n_441),
.B1(n_451),
.B2(n_446),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_481),
.A2(n_487),
.B1(n_425),
.B2(n_455),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_476),
.B(n_460),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_483),
.B(n_486),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_460),
.B(n_444),
.C(n_448),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_485),
.B(n_464),
.C(n_472),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_461),
.B(n_444),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_469),
.A2(n_445),
.B1(n_430),
.B2(n_415),
.Y(n_487)
);

AO21x1_ASAP7_75t_L g488 ( 
.A1(n_478),
.A2(n_450),
.B(n_422),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_488),
.B(n_497),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_473),
.A2(n_456),
.B(n_440),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_489),
.A2(n_463),
.B(n_477),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_459),
.B(n_413),
.Y(n_491)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_491),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_493),
.B(n_465),
.Y(n_511)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_471),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_498),
.B(n_503),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_482),
.B(n_485),
.C(n_484),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_499),
.B(n_506),
.C(n_513),
.Y(n_516)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_502),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_490),
.B(n_470),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_492),
.A2(n_430),
.B1(n_474),
.B2(n_458),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_504),
.A2(n_496),
.B1(n_489),
.B2(n_488),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_505),
.A2(n_429),
.B1(n_377),
.B2(n_380),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_482),
.B(n_484),
.C(n_475),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_495),
.A2(n_425),
.B(n_413),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_507),
.B(n_487),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_490),
.B(n_420),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_509),
.A2(n_510),
.B1(n_512),
.B2(n_387),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_480),
.B(n_454),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_511),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_480),
.B(n_392),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_481),
.B(n_465),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_508),
.A2(n_497),
.B(n_495),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_514),
.B(n_519),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_515),
.B(n_521),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_499),
.B(n_492),
.C(n_496),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_517),
.B(n_523),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_506),
.B(n_494),
.C(n_491),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_501),
.A2(n_494),
.B1(n_376),
.B2(n_386),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_524),
.A2(n_526),
.B1(n_377),
.B2(n_243),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_498),
.B(n_429),
.C(n_376),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_525),
.B(n_513),
.C(n_504),
.Y(n_531)
);

A2O1A1Ixp33_ASAP7_75t_SL g527 ( 
.A1(n_515),
.A2(n_507),
.B(n_508),
.C(n_505),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_527),
.B(n_529),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_520),
.B(n_511),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_SL g530 ( 
.A(n_518),
.B(n_502),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_530),
.B(n_531),
.C(n_523),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_516),
.B(n_500),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_533),
.B(n_536),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_516),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_534),
.B(n_525),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_538),
.B(n_542),
.C(n_527),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_528),
.B(n_517),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_539),
.A2(n_541),
.B(n_535),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_532),
.B(n_522),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_SL g547 ( 
.A1(n_543),
.A2(n_544),
.B(n_545),
.Y(n_547)
);

NOR3xp33_ASAP7_75t_L g544 ( 
.A(n_540),
.B(n_535),
.C(n_539),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_537),
.A2(n_527),
.B(n_526),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_SL g548 ( 
.A(n_546),
.B(n_377),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_548),
.B(n_243),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_549),
.B(n_547),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_550),
.B(n_263),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_245),
.C(n_288),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_552),
.A2(n_0),
.B1(n_1),
.B2(n_539),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_553),
.B(n_0),
.Y(n_554)
);


endmodule