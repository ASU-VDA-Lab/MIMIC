module real_aes_6602_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g113 ( .A(n_0), .Y(n_113) );
INVx1_ASAP7_75t_L g483 ( .A(n_1), .Y(n_483) );
INVx1_ASAP7_75t_L g196 ( .A(n_2), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_3), .A2(n_35), .B1(n_152), .B2(n_499), .Y(n_509) );
AOI21xp33_ASAP7_75t_L g176 ( .A1(n_4), .A2(n_133), .B(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_5), .B(n_126), .Y(n_474) );
AND2x6_ASAP7_75t_L g138 ( .A(n_6), .B(n_139), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_7), .A2(n_235), .B(n_236), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_8), .B(n_36), .Y(n_114) );
INVx1_ASAP7_75t_L g744 ( .A(n_8), .Y(n_744) );
INVx1_ASAP7_75t_L g183 ( .A(n_9), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_10), .B(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g131 ( .A(n_11), .Y(n_131) );
INVx1_ASAP7_75t_L g478 ( .A(n_12), .Y(n_478) );
INVx1_ASAP7_75t_L g241 ( .A(n_13), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_14), .B(n_164), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_15), .B(n_127), .Y(n_455) );
AO32x2_ASAP7_75t_L g507 ( .A1(n_16), .A2(n_126), .A3(n_161), .B1(n_461), .B2(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_17), .B(n_152), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_18), .B(n_147), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_19), .B(n_127), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_20), .A2(n_50), .B1(n_152), .B2(n_499), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_21), .B(n_133), .Y(n_207) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_22), .A2(n_74), .B1(n_152), .B2(n_164), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_23), .B(n_152), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_24), .B(n_155), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_25), .A2(n_239), .B(n_240), .C(n_242), .Y(n_238) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_26), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_27), .B(n_185), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_28), .B(n_181), .Y(n_198) );
INVx1_ASAP7_75t_L g170 ( .A(n_29), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_30), .B(n_185), .Y(n_522) );
INVx2_ASAP7_75t_L g136 ( .A(n_31), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_32), .B(n_152), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_33), .B(n_185), .Y(n_500) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_34), .A2(n_138), .B(n_142), .C(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_36), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g168 ( .A(n_37), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_38), .B(n_181), .Y(n_251) );
AOI222xp33_ASAP7_75t_L g115 ( .A1(n_39), .A2(n_43), .B1(n_116), .B2(n_725), .C1(n_730), .C2(n_731), .Y(n_115) );
CKINVDCx14_ASAP7_75t_R g730 ( .A(n_39), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_40), .B(n_152), .Y(n_468) );
AOI22xp33_ASAP7_75t_SL g99 ( .A1(n_41), .A2(n_100), .B1(n_739), .B2(n_749), .Y(n_99) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_42), .A2(n_85), .B1(n_214), .B2(n_499), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_44), .B(n_152), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_45), .B(n_152), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_46), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g171 ( .A(n_47), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_48), .B(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_49), .B(n_133), .Y(n_229) );
AOI22xp33_ASAP7_75t_SL g460 ( .A1(n_51), .A2(n_60), .B1(n_152), .B2(n_164), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g163 ( .A1(n_52), .A2(n_142), .B1(n_164), .B2(n_166), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g217 ( .A(n_53), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_54), .B(n_152), .Y(n_493) );
CKINVDCx16_ASAP7_75t_R g193 ( .A(n_55), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_56), .B(n_152), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_57), .A2(n_151), .B(n_180), .C(n_182), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g255 ( .A(n_58), .Y(n_255) );
INVx1_ASAP7_75t_L g178 ( .A(n_59), .Y(n_178) );
INVx1_ASAP7_75t_L g139 ( .A(n_61), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_62), .B(n_152), .Y(n_484) );
INVx1_ASAP7_75t_L g130 ( .A(n_63), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_64), .Y(n_105) );
AO32x2_ASAP7_75t_L g502 ( .A1(n_65), .A2(n_126), .A3(n_221), .B1(n_461), .B2(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g541 ( .A(n_66), .Y(n_541) );
INVx1_ASAP7_75t_L g517 ( .A(n_67), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_SL g146 ( .A1(n_68), .A2(n_147), .B(n_148), .C(n_151), .Y(n_146) );
INVxp67_ASAP7_75t_L g149 ( .A(n_69), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_70), .B(n_164), .Y(n_518) );
INVx1_ASAP7_75t_L g748 ( .A(n_71), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_72), .Y(n_174) );
INVx1_ASAP7_75t_L g248 ( .A(n_73), .Y(n_248) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_75), .A2(n_138), .B(n_142), .C(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_76), .B(n_499), .Y(n_498) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_77), .A2(n_117), .B1(n_118), .B2(n_735), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_77), .Y(n_735) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_78), .B(n_164), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_79), .B(n_197), .Y(n_210) );
INVx2_ASAP7_75t_L g128 ( .A(n_80), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_81), .B(n_147), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_82), .B(n_164), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_83), .A2(n_138), .B(n_142), .C(n_195), .Y(n_194) );
OR2x2_ASAP7_75t_L g110 ( .A(n_84), .B(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g445 ( .A(n_84), .B(n_112), .Y(n_445) );
INVx2_ASAP7_75t_L g447 ( .A(n_84), .Y(n_447) );
NAND3xp33_ASAP7_75t_SL g745 ( .A(n_84), .B(n_113), .C(n_746), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_86), .A2(n_98), .B1(n_164), .B2(n_165), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_87), .B(n_185), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_88), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_89), .A2(n_138), .B(n_142), .C(n_224), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_90), .Y(n_231) );
INVx1_ASAP7_75t_L g145 ( .A(n_91), .Y(n_145) );
CKINVDCx16_ASAP7_75t_R g237 ( .A(n_92), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_93), .B(n_197), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_94), .B(n_164), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_95), .B(n_126), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g132 ( .A1(n_96), .A2(n_133), .B(n_140), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_97), .B(n_748), .Y(n_747) );
AOI22x1_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_115), .B1(n_732), .B2(n_733), .Y(n_100) );
NOR2xp33_ASAP7_75t_L g101 ( .A(n_102), .B(n_106), .Y(n_101) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
BUFx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_SL g732 ( .A(n_104), .Y(n_732) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g733 ( .A1(n_106), .A2(n_734), .B(n_736), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_110), .Y(n_738) );
NOR2x2_ASAP7_75t_L g731 ( .A(n_111), .B(n_447), .Y(n_731) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g446 ( .A(n_112), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OAI22x1_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_443), .B1(n_446), .B2(n_448), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_118), .A2(n_726), .B1(n_727), .B2(n_729), .Y(n_725) );
AND2x2_ASAP7_75t_SL g118 ( .A(n_119), .B(n_380), .Y(n_118) );
NOR4xp25_ASAP7_75t_L g119 ( .A(n_120), .B(n_310), .C(n_341), .D(n_360), .Y(n_119) );
NAND4xp25_ASAP7_75t_L g120 ( .A(n_121), .B(n_268), .C(n_283), .D(n_301), .Y(n_120) );
AOI222xp33_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_203), .B1(n_244), .B2(n_256), .C1(n_261), .C2(n_263), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_186), .Y(n_122) );
INVx1_ASAP7_75t_L g324 ( .A(n_123), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_157), .Y(n_123) );
AND2x2_ASAP7_75t_L g187 ( .A(n_124), .B(n_175), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_124), .B(n_190), .Y(n_353) );
INVx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g260 ( .A(n_125), .B(n_159), .Y(n_260) );
AND2x2_ASAP7_75t_L g269 ( .A(n_125), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g295 ( .A(n_125), .Y(n_295) );
AND2x2_ASAP7_75t_L g316 ( .A(n_125), .B(n_159), .Y(n_316) );
BUFx2_ASAP7_75t_L g339 ( .A(n_125), .Y(n_339) );
AND2x2_ASAP7_75t_L g363 ( .A(n_125), .B(n_160), .Y(n_363) );
AND2x2_ASAP7_75t_L g427 ( .A(n_125), .B(n_175), .Y(n_427) );
OA21x2_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_132), .B(n_154), .Y(n_125) );
INVx4_ASAP7_75t_L g156 ( .A(n_126), .Y(n_156) );
OA21x2_ASAP7_75t_L g465 ( .A1(n_126), .A2(n_466), .B(n_474), .Y(n_465) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g161 ( .A(n_127), .Y(n_161) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
AND2x2_ASAP7_75t_SL g185 ( .A(n_128), .B(n_129), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
BUFx2_ASAP7_75t_L g235 ( .A(n_133), .Y(n_235) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_138), .Y(n_133) );
NAND2x1p5_ASAP7_75t_L g172 ( .A(n_134), .B(n_138), .Y(n_172) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx1_ASAP7_75t_L g473 ( .A(n_135), .Y(n_473) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g143 ( .A(n_136), .Y(n_143) );
INVx1_ASAP7_75t_L g165 ( .A(n_136), .Y(n_165) );
INVx1_ASAP7_75t_L g144 ( .A(n_137), .Y(n_144) );
INVx1_ASAP7_75t_L g147 ( .A(n_137), .Y(n_147) );
INVx3_ASAP7_75t_L g150 ( .A(n_137), .Y(n_150) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_137), .Y(n_167) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_137), .Y(n_181) );
INVx4_ASAP7_75t_SL g153 ( .A(n_138), .Y(n_153) );
BUFx3_ASAP7_75t_L g461 ( .A(n_138), .Y(n_461) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_138), .A2(n_467), .B(n_470), .Y(n_466) );
OAI21xp5_ASAP7_75t_L g476 ( .A1(n_138), .A2(n_477), .B(n_481), .Y(n_476) );
OAI21xp5_ASAP7_75t_L g491 ( .A1(n_138), .A2(n_492), .B(n_496), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_138), .A2(n_516), .B(n_519), .Y(n_515) );
O2A1O1Ixp33_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_145), .B(n_146), .C(n_153), .Y(n_140) );
O2A1O1Ixp33_ASAP7_75t_L g177 ( .A1(n_141), .A2(n_153), .B(n_178), .C(n_179), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_141), .A2(n_153), .B(n_237), .C(n_238), .Y(n_236) );
INVx5_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x6_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_143), .Y(n_152) );
BUFx3_ASAP7_75t_L g214 ( .A(n_143), .Y(n_214) );
INVx1_ASAP7_75t_L g499 ( .A(n_143), .Y(n_499) );
INVx1_ASAP7_75t_L g495 ( .A(n_147), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_150), .B(n_183), .Y(n_182) );
INVx5_ASAP7_75t_L g197 ( .A(n_150), .Y(n_197) );
OAI22xp5_ASAP7_75t_SL g503 ( .A1(n_150), .A2(n_181), .B1(n_504), .B2(n_505), .Y(n_503) );
O2A1O1Ixp5_ASAP7_75t_SL g516 ( .A1(n_151), .A2(n_197), .B(n_517), .C(n_518), .Y(n_516) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_152), .Y(n_228) );
OAI22xp33_ASAP7_75t_L g162 ( .A1(n_153), .A2(n_163), .B1(n_171), .B2(n_172), .Y(n_162) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_155), .A2(n_176), .B(n_184), .Y(n_175) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_SL g216 ( .A(n_156), .B(n_217), .Y(n_216) );
NAND3xp33_ASAP7_75t_L g456 ( .A(n_156), .B(n_457), .C(n_461), .Y(n_456) );
AO21x1_ASAP7_75t_L g549 ( .A1(n_156), .A2(n_457), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g328 ( .A(n_157), .B(n_259), .Y(n_328) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_158), .B(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g158 ( .A(n_159), .B(n_175), .Y(n_158) );
OR2x2_ASAP7_75t_L g288 ( .A(n_159), .B(n_191), .Y(n_288) );
AND2x2_ASAP7_75t_L g300 ( .A(n_159), .B(n_259), .Y(n_300) );
BUFx2_ASAP7_75t_L g432 ( .A(n_159), .Y(n_432) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
OR2x2_ASAP7_75t_L g189 ( .A(n_160), .B(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g282 ( .A(n_160), .B(n_191), .Y(n_282) );
AND2x2_ASAP7_75t_L g335 ( .A(n_160), .B(n_175), .Y(n_335) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_160), .Y(n_371) );
AO21x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_173), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_161), .B(n_174), .Y(n_173) );
AO21x2_ASAP7_75t_L g191 ( .A1(n_161), .A2(n_192), .B(n_200), .Y(n_191) );
INVx2_ASAP7_75t_L g215 ( .A(n_161), .Y(n_215) );
INVx2_ASAP7_75t_L g199 ( .A(n_164), .Y(n_199) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
OAI22xp5_ASAP7_75t_SL g166 ( .A1(n_167), .A2(n_168), .B1(n_169), .B2(n_170), .Y(n_166) );
INVx2_ASAP7_75t_L g169 ( .A(n_167), .Y(n_169) );
INVx4_ASAP7_75t_L g239 ( .A(n_167), .Y(n_239) );
OAI21xp5_ASAP7_75t_L g192 ( .A1(n_172), .A2(n_193), .B(n_194), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g247 ( .A1(n_172), .A2(n_248), .B(n_249), .Y(n_247) );
AND2x2_ASAP7_75t_L g258 ( .A(n_175), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_SL g270 ( .A(n_175), .Y(n_270) );
INVx2_ASAP7_75t_L g281 ( .A(n_175), .Y(n_281) );
BUFx2_ASAP7_75t_L g305 ( .A(n_175), .Y(n_305) );
AND2x2_ASAP7_75t_SL g362 ( .A(n_175), .B(n_363), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_180), .A2(n_497), .B(n_498), .Y(n_496) );
O2A1O1Ixp5_ASAP7_75t_L g540 ( .A1(n_180), .A2(n_482), .B(n_541), .C(n_542), .Y(n_540) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx4_ASAP7_75t_L g227 ( .A(n_181), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_181), .A2(n_458), .B1(n_459), .B2(n_460), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_181), .A2(n_459), .B1(n_509), .B2(n_510), .Y(n_508) );
INVx1_ASAP7_75t_L g202 ( .A(n_185), .Y(n_202) );
INVx2_ASAP7_75t_L g221 ( .A(n_185), .Y(n_221) );
OA21x2_ASAP7_75t_L g233 ( .A1(n_185), .A2(n_234), .B(n_243), .Y(n_233) );
OA21x2_ASAP7_75t_L g490 ( .A1(n_185), .A2(n_491), .B(n_500), .Y(n_490) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_185), .A2(n_515), .B(n_522), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_188), .Y(n_186) );
AOI332xp33_ASAP7_75t_L g283 ( .A1(n_187), .A2(n_284), .A3(n_288), .B1(n_289), .B2(n_293), .B3(n_296), .C1(n_297), .C2(n_299), .Y(n_283) );
NAND2x1_ASAP7_75t_L g368 ( .A(n_187), .B(n_259), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_187), .B(n_273), .Y(n_419) );
A2O1A1Ixp33_ASAP7_75t_SL g301 ( .A1(n_188), .A2(n_302), .B(n_305), .C(n_306), .Y(n_301) );
AND2x2_ASAP7_75t_L g440 ( .A(n_188), .B(n_281), .Y(n_440) );
INVx3_ASAP7_75t_SL g188 ( .A(n_189), .Y(n_188) );
OR2x2_ASAP7_75t_L g337 ( .A(n_189), .B(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g342 ( .A(n_189), .B(n_339), .Y(n_342) );
INVx1_ASAP7_75t_L g273 ( .A(n_190), .Y(n_273) );
AND2x2_ASAP7_75t_L g376 ( .A(n_190), .B(n_335), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_190), .B(n_316), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_190), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_190), .B(n_294), .Y(n_402) );
INVx3_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx3_ASAP7_75t_L g259 ( .A(n_191), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_198), .C(n_199), .Y(n_195) );
INVx2_ASAP7_75t_L g459 ( .A(n_197), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_197), .A2(n_468), .B(n_469), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_197), .A2(n_538), .B(n_539), .Y(n_537) );
O2A1O1Ixp33_ASAP7_75t_L g477 ( .A1(n_199), .A2(n_478), .B(n_479), .C(n_480), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_202), .B(n_231), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_202), .B(n_255), .Y(n_254) );
OAI31xp33_ASAP7_75t_L g441 ( .A1(n_203), .A2(n_362), .A3(n_369), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_218), .Y(n_203) );
AND2x2_ASAP7_75t_L g244 ( .A(n_204), .B(n_245), .Y(n_244) );
NAND2x1_ASAP7_75t_SL g264 ( .A(n_204), .B(n_265), .Y(n_264) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_204), .Y(n_351) );
AND2x2_ASAP7_75t_L g356 ( .A(n_204), .B(n_267), .Y(n_356) );
INVx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_205), .A2(n_269), .B(n_271), .C(n_274), .Y(n_268) );
OR2x2_ASAP7_75t_L g285 ( .A(n_205), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g298 ( .A(n_205), .Y(n_298) );
AND2x2_ASAP7_75t_L g304 ( .A(n_205), .B(n_246), .Y(n_304) );
INVx2_ASAP7_75t_L g322 ( .A(n_205), .Y(n_322) );
AND2x2_ASAP7_75t_L g333 ( .A(n_205), .B(n_287), .Y(n_333) );
AND2x2_ASAP7_75t_L g365 ( .A(n_205), .B(n_323), .Y(n_365) );
AND2x2_ASAP7_75t_L g369 ( .A(n_205), .B(n_292), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_205), .B(n_218), .Y(n_374) );
AND2x2_ASAP7_75t_L g408 ( .A(n_205), .B(n_409), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_205), .B(n_311), .Y(n_442) );
OR2x6_ASAP7_75t_L g205 ( .A(n_206), .B(n_216), .Y(n_205) );
AOI21xp5_ASAP7_75t_SL g206 ( .A1(n_207), .A2(n_208), .B(n_215), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_212), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_212), .A2(n_251), .B(n_252), .Y(n_250) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g242 ( .A(n_214), .Y(n_242) );
INVx1_ASAP7_75t_L g253 ( .A(n_215), .Y(n_253) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_215), .A2(n_476), .B(n_485), .Y(n_475) );
OA21x2_ASAP7_75t_L g535 ( .A1(n_215), .A2(n_536), .B(n_543), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_218), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g350 ( .A(n_218), .Y(n_350) );
AND2x2_ASAP7_75t_L g412 ( .A(n_218), .B(n_333), .Y(n_412) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_232), .Y(n_218) );
OR2x2_ASAP7_75t_L g266 ( .A(n_219), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g276 ( .A(n_219), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_219), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g384 ( .A(n_219), .Y(n_384) );
AND2x2_ASAP7_75t_L g401 ( .A(n_219), .B(n_246), .Y(n_401) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g292 ( .A(n_220), .B(n_232), .Y(n_292) );
AND2x2_ASAP7_75t_L g321 ( .A(n_220), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g332 ( .A(n_220), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_220), .B(n_287), .Y(n_423) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_230), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_229), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_228), .Y(n_224) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g245 ( .A(n_233), .B(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g267 ( .A(n_233), .Y(n_267) );
AND2x2_ASAP7_75t_L g323 ( .A(n_233), .B(n_287), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_239), .B(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g480 ( .A(n_239), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_239), .A2(n_520), .B(n_521), .Y(n_519) );
INVx1_ASAP7_75t_L g425 ( .A(n_244), .Y(n_425) );
INVx1_ASAP7_75t_L g429 ( .A(n_245), .Y(n_429) );
INVx2_ASAP7_75t_L g287 ( .A(n_246), .Y(n_287) );
AO21x2_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_253), .B(n_254), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_257), .B(n_260), .Y(n_256) );
INVx1_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_258), .B(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_258), .B(n_363), .Y(n_421) );
OR2x2_ASAP7_75t_L g262 ( .A(n_259), .B(n_260), .Y(n_262) );
INVx1_ASAP7_75t_SL g314 ( .A(n_259), .Y(n_314) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AOI221xp5_ASAP7_75t_L g317 ( .A1(n_265), .A2(n_318), .B1(n_320), .B2(n_324), .C(n_325), .Y(n_317) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g345 ( .A(n_266), .B(n_309), .Y(n_345) );
INVx2_ASAP7_75t_L g277 ( .A(n_267), .Y(n_277) );
INVx1_ASAP7_75t_L g303 ( .A(n_267), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_267), .B(n_287), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_267), .B(n_290), .Y(n_397) );
INVx1_ASAP7_75t_L g405 ( .A(n_267), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_269), .B(n_273), .Y(n_319) );
AND2x4_ASAP7_75t_L g294 ( .A(n_270), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g407 ( .A(n_273), .B(n_363), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_275), .B(n_278), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_276), .B(n_308), .Y(n_307) );
INVxp67_ASAP7_75t_L g415 ( .A(n_277), .Y(n_415) );
INVxp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
INVx1_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g315 ( .A(n_281), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g387 ( .A(n_281), .B(n_363), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_281), .B(n_300), .Y(n_393) );
AOI322xp5_ASAP7_75t_L g347 ( .A1(n_282), .A2(n_316), .A3(n_323), .B1(n_348), .B2(n_351), .C1(n_352), .C2(n_354), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_282), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g413 ( .A(n_285), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g359 ( .A(n_286), .Y(n_359) );
INVx2_ASAP7_75t_L g290 ( .A(n_287), .Y(n_290) );
INVx1_ASAP7_75t_L g349 ( .A(n_287), .Y(n_349) );
CKINVDCx16_ASAP7_75t_R g296 ( .A(n_288), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
AND2x2_ASAP7_75t_L g385 ( .A(n_290), .B(n_298), .Y(n_385) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g297 ( .A(n_292), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g340 ( .A(n_292), .B(n_333), .Y(n_340) );
AND2x2_ASAP7_75t_L g344 ( .A(n_292), .B(n_304), .Y(n_344) );
OAI21xp33_ASAP7_75t_SL g354 ( .A1(n_293), .A2(n_355), .B(n_357), .Y(n_354) );
OAI22xp33_ASAP7_75t_L g424 ( .A1(n_293), .A2(n_425), .B1(n_426), .B2(n_428), .Y(n_424) );
INVx3_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g299 ( .A(n_294), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_294), .B(n_314), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_296), .B(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_L g436 ( .A(n_303), .Y(n_436) );
INVx4_ASAP7_75t_L g309 ( .A(n_304), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_304), .B(n_331), .Y(n_379) );
INVx1_ASAP7_75t_SL g391 ( .A(n_305), .Y(n_391) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NOR2xp67_ASAP7_75t_L g404 ( .A(n_309), .B(n_405), .Y(n_404) );
OAI211xp5_ASAP7_75t_SL g310 ( .A1(n_311), .A2(n_312), .B(n_317), .C(n_334), .Y(n_310) );
OAI221xp5_ASAP7_75t_SL g430 ( .A1(n_312), .A2(n_350), .B1(n_429), .B2(n_431), .C(n_433), .Y(n_430) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_314), .B(n_427), .Y(n_426) );
OAI31xp33_ASAP7_75t_L g406 ( .A1(n_315), .A2(n_392), .A3(n_407), .B(n_408), .Y(n_406) );
INVx1_ASAP7_75t_L g346 ( .A(n_316), .Y(n_346) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
INVx1_ASAP7_75t_L g396 ( .A(n_321), .Y(n_396) );
AND2x2_ASAP7_75t_L g409 ( .A(n_323), .B(n_332), .Y(n_409) );
AOI21xp33_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_327), .B(n_329), .Y(n_325) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVxp67_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_333), .B(n_436), .Y(n_435) );
OAI21xp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_336), .B(n_340), .Y(n_334) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OAI221xp5_ASAP7_75t_SL g341 ( .A1(n_342), .A2(n_343), .B1(n_345), .B2(n_346), .C(n_347), .Y(n_341) );
A2O1A1Ixp33_ASAP7_75t_L g410 ( .A1(n_342), .A2(n_411), .B(n_413), .C(n_416), .Y(n_410) );
CKINVDCx16_ASAP7_75t_R g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_345), .B(n_395), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx1_ASAP7_75t_L g372 ( .A(n_353), .Y(n_372) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g358 ( .A(n_356), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g400 ( .A(n_356), .B(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI211xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_364), .B(n_366), .C(n_375), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI221xp5_ASAP7_75t_L g437 ( .A1(n_364), .A2(n_374), .B1(n_438), .B2(n_439), .C(n_441), .Y(n_437) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_369), .B1(n_370), .B2(n_373), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OAI21xp5_ASAP7_75t_SL g375 ( .A1(n_376), .A2(n_377), .B(n_378), .Y(n_375) );
INVx1_ASAP7_75t_SL g438 ( .A(n_377), .Y(n_438) );
INVxp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NOR4xp25_ASAP7_75t_L g380 ( .A(n_381), .B(n_410), .C(n_430), .D(n_437), .Y(n_380) );
OAI211xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_386), .B(n_388), .C(n_406), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
INVxp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
O2A1O1Ixp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_392), .B(n_394), .C(n_398), .Y(n_388) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_SL g417 ( .A(n_395), .Y(n_417) );
OR2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
OR2x2_ASAP7_75t_L g428 ( .A(n_396), .B(n_429), .Y(n_428) );
OAI21xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_402), .B(n_403), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B1(n_420), .B2(n_422), .C(n_424), .Y(n_416) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVxp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_427), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g726 ( .A(n_444), .Y(n_726) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g728 ( .A(n_446), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_448), .Y(n_729) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_SL g449 ( .A(n_450), .B(n_659), .Y(n_449) );
NOR5xp2_ASAP7_75t_L g450 ( .A(n_451), .B(n_572), .C(n_618), .D(n_631), .E(n_643), .Y(n_450) );
OAI211xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_486), .B(n_526), .C(n_553), .Y(n_451) );
INVx1_ASAP7_75t_SL g654 ( .A(n_452), .Y(n_654) );
OR2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_462), .Y(n_452) );
AND2x2_ASAP7_75t_L g578 ( .A(n_453), .B(n_463), .Y(n_578) );
AND2x2_ASAP7_75t_L g606 ( .A(n_453), .B(n_552), .Y(n_606) );
AND2x2_ASAP7_75t_L g614 ( .A(n_453), .B(n_557), .Y(n_614) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g544 ( .A(n_454), .B(n_464), .Y(n_544) );
INVx2_ASAP7_75t_L g556 ( .A(n_454), .Y(n_556) );
AND2x2_ASAP7_75t_L g681 ( .A(n_454), .B(n_623), .Y(n_681) );
OR2x2_ASAP7_75t_L g683 ( .A(n_454), .B(n_684), .Y(n_683) );
AND2x4_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
INVx1_ASAP7_75t_L g550 ( .A(n_455), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_459), .A2(n_471), .B(n_472), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_459), .A2(n_482), .B(n_483), .C(n_484), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g536 ( .A1(n_461), .A2(n_537), .B(n_540), .Y(n_536) );
INVx2_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g594 ( .A(n_463), .B(n_566), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_463), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g708 ( .A(n_463), .B(n_548), .Y(n_708) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_475), .Y(n_463) );
AND2x2_ASAP7_75t_L g551 ( .A(n_464), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g598 ( .A(n_464), .Y(n_598) );
AND2x2_ASAP7_75t_L g623 ( .A(n_464), .B(n_535), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_464), .B(n_656), .Y(n_693) );
INVx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g557 ( .A(n_465), .B(n_535), .Y(n_557) );
AND2x2_ASAP7_75t_L g571 ( .A(n_465), .B(n_534), .Y(n_571) );
AND2x2_ASAP7_75t_L g588 ( .A(n_465), .B(n_475), .Y(n_588) );
AND2x2_ASAP7_75t_L g645 ( .A(n_465), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_465), .B(n_552), .Y(n_658) );
AND2x2_ASAP7_75t_L g710 ( .A(n_465), .B(n_635), .Y(n_710) );
INVx2_ASAP7_75t_L g482 ( .A(n_473), .Y(n_482) );
AND2x2_ASAP7_75t_L g533 ( .A(n_475), .B(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g552 ( .A(n_475), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_475), .B(n_535), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_511), .B(n_523), .Y(n_486) );
INVx1_ASAP7_75t_SL g642 ( .A(n_487), .Y(n_642) );
AND2x4_ASAP7_75t_L g487 ( .A(n_488), .B(n_501), .Y(n_487) );
BUFx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_SL g530 ( .A(n_489), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g525 ( .A(n_490), .Y(n_525) );
INVx1_ASAP7_75t_L g562 ( .A(n_490), .Y(n_562) );
AND2x2_ASAP7_75t_L g583 ( .A(n_490), .B(n_506), .Y(n_583) );
AND2x2_ASAP7_75t_L g617 ( .A(n_490), .B(n_507), .Y(n_617) );
OR2x2_ASAP7_75t_L g636 ( .A(n_490), .B(n_513), .Y(n_636) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_490), .Y(n_650) );
AND2x2_ASAP7_75t_L g663 ( .A(n_490), .B(n_664), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_494), .B(n_495), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_501), .A2(n_585), .B1(n_586), .B2(n_595), .Y(n_584) );
AND2x2_ASAP7_75t_L g668 ( .A(n_501), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_506), .Y(n_501) );
INVx1_ASAP7_75t_L g529 ( .A(n_502), .Y(n_529) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_502), .Y(n_566) );
INVx1_ASAP7_75t_L g577 ( .A(n_502), .Y(n_577) );
AND2x2_ASAP7_75t_L g592 ( .A(n_502), .B(n_507), .Y(n_592) );
OR2x2_ASAP7_75t_L g546 ( .A(n_506), .B(n_531), .Y(n_546) );
AND2x2_ASAP7_75t_L g576 ( .A(n_506), .B(n_577), .Y(n_576) );
NOR2xp67_ASAP7_75t_L g664 ( .A(n_506), .B(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g524 ( .A(n_507), .B(n_525), .Y(n_524) );
BUFx2_ASAP7_75t_L g633 ( .A(n_507), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_511), .B(n_649), .Y(n_648) );
BUFx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g611 ( .A(n_512), .B(n_577), .Y(n_611) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g523 ( .A(n_513), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g582 ( .A(n_513), .Y(n_582) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g531 ( .A(n_514), .Y(n_531) );
OR2x2_ASAP7_75t_L g561 ( .A(n_514), .B(n_562), .Y(n_561) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_514), .Y(n_616) );
AOI32xp33_ASAP7_75t_L g653 ( .A1(n_523), .A2(n_583), .A3(n_654), .B1(n_655), .B2(n_657), .Y(n_653) );
AND2x2_ASAP7_75t_L g579 ( .A(n_524), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_524), .B(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_524), .B(n_611), .Y(n_697) );
INVx1_ASAP7_75t_L g702 ( .A(n_524), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_532), .B1(n_545), .B2(n_547), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_530), .Y(n_527) );
AND2x2_ASAP7_75t_L g632 ( .A(n_528), .B(n_633), .Y(n_632) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_529), .B(n_531), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_530), .A2(n_554), .B1(n_558), .B2(n_568), .Y(n_553) );
AND2x2_ASAP7_75t_L g575 ( .A(n_530), .B(n_576), .Y(n_575) );
A2O1A1Ixp33_ASAP7_75t_L g626 ( .A1(n_530), .A2(n_544), .B(n_592), .C(n_627), .Y(n_626) );
OAI332xp33_ASAP7_75t_L g631 ( .A1(n_530), .A2(n_632), .A3(n_634), .B1(n_636), .B2(n_637), .B3(n_639), .C1(n_640), .C2(n_642), .Y(n_631) );
INVx2_ASAP7_75t_L g672 ( .A(n_530), .Y(n_672) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_531), .Y(n_590) );
INVx1_ASAP7_75t_L g665 ( .A(n_531), .Y(n_665) );
AND2x2_ASAP7_75t_L g719 ( .A(n_531), .B(n_583), .Y(n_719) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_544), .Y(n_532) );
AND2x2_ASAP7_75t_L g599 ( .A(n_534), .B(n_549), .Y(n_599) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g548 ( .A(n_535), .B(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g647 ( .A(n_535), .B(n_549), .Y(n_647) );
INVx1_ASAP7_75t_L g656 ( .A(n_535), .Y(n_656) );
INVx1_ASAP7_75t_L g630 ( .A(n_544), .Y(n_630) );
INVxp67_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g714 ( .A(n_546), .B(n_566), .Y(n_714) );
INVx1_ASAP7_75t_SL g625 ( .A(n_547), .Y(n_625) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_551), .Y(n_547) );
AND2x2_ASAP7_75t_L g652 ( .A(n_548), .B(n_610), .Y(n_652) );
INVx1_ASAP7_75t_L g671 ( .A(n_548), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_548), .B(n_638), .Y(n_673) );
INVx1_ASAP7_75t_L g570 ( .A(n_549), .Y(n_570) );
AND2x2_ASAP7_75t_L g574 ( .A(n_551), .B(n_555), .Y(n_574) );
AND2x2_ASAP7_75t_L g641 ( .A(n_551), .B(n_599), .Y(n_641) );
INVx2_ASAP7_75t_L g684 ( .A(n_551), .Y(n_684) );
INVx2_ASAP7_75t_L g567 ( .A(n_552), .Y(n_567) );
AND2x2_ASAP7_75t_L g569 ( .A(n_552), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_557), .Y(n_554) );
INVx1_ASAP7_75t_L g585 ( .A(n_555), .Y(n_585) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_556), .B(n_629), .Y(n_635) );
OR2x2_ASAP7_75t_L g699 ( .A(n_556), .B(n_658), .Y(n_699) );
INVx1_ASAP7_75t_L g723 ( .A(n_556), .Y(n_723) );
INVx1_ASAP7_75t_L g679 ( .A(n_557), .Y(n_679) );
AND2x2_ASAP7_75t_L g724 ( .A(n_557), .B(n_567), .Y(n_724) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_561), .A2(n_587), .B1(n_589), .B2(n_593), .Y(n_586) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OAI322xp33_ASAP7_75t_SL g670 ( .A1(n_564), .A2(n_671), .A3(n_672), .B1(n_673), .B2(n_674), .C1(n_677), .C2(n_679), .Y(n_670) );
OR2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .Y(n_564) );
AND2x2_ASAP7_75t_L g667 ( .A(n_565), .B(n_583), .Y(n_667) );
OR2x2_ASAP7_75t_L g701 ( .A(n_565), .B(n_702), .Y(n_701) );
OR2x2_ASAP7_75t_L g704 ( .A(n_565), .B(n_636), .Y(n_704) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g649 ( .A(n_566), .B(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g705 ( .A(n_566), .B(n_636), .Y(n_705) );
INVx3_ASAP7_75t_L g638 ( .A(n_567), .Y(n_638) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
INVx1_ASAP7_75t_L g694 ( .A(n_569), .Y(n_694) );
AOI222xp33_ASAP7_75t_L g573 ( .A1(n_571), .A2(n_574), .B1(n_575), .B2(n_578), .C1(n_579), .C2(n_581), .Y(n_573) );
INVx1_ASAP7_75t_L g604 ( .A(n_571), .Y(n_604) );
NAND3xp33_ASAP7_75t_SL g572 ( .A(n_573), .B(n_584), .C(n_601), .Y(n_572) );
AND2x2_ASAP7_75t_L g689 ( .A(n_576), .B(n_590), .Y(n_689) );
BUFx2_ASAP7_75t_L g580 ( .A(n_577), .Y(n_580) );
INVx1_ASAP7_75t_L g621 ( .A(n_577), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_578), .A2(n_614), .B1(n_667), .B2(n_668), .C(n_670), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_580), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_583), .Y(n_607) );
AND2x2_ASAP7_75t_L g620 ( .A(n_583), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_588), .B(n_599), .Y(n_600) );
OR2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
OAI21xp33_ASAP7_75t_L g595 ( .A1(n_590), .A2(n_596), .B(n_600), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_590), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g687 ( .A(n_592), .B(n_669), .Y(n_687) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
INVx1_ASAP7_75t_L g610 ( .A(n_598), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_599), .B(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g716 ( .A(n_599), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_607), .B1(n_608), .B2(n_611), .C(n_612), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_603), .B(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g712 ( .A(n_611), .B(n_617), .Y(n_712) );
INVxp67_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
OAI31xp33_ASAP7_75t_SL g680 ( .A1(n_615), .A2(n_654), .A3(n_681), .B(n_682), .Y(n_680) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVx1_ASAP7_75t_L g669 ( .A(n_616), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g720 ( .A(n_617), .B(n_621), .Y(n_720) );
OAI221xp5_ASAP7_75t_SL g618 ( .A1(n_619), .A2(n_622), .B1(n_624), .B2(n_625), .C(n_626), .Y(n_618) );
INVx1_ASAP7_75t_L g624 ( .A(n_620), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_623), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx1_ASAP7_75t_L g639 ( .A(n_632), .Y(n_639) );
INVx2_ASAP7_75t_L g675 ( .A(n_633), .Y(n_675) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g661 ( .A(n_638), .B(n_647), .Y(n_661) );
A2O1A1Ixp33_ASAP7_75t_L g711 ( .A1(n_638), .A2(n_655), .B(n_712), .C(n_713), .Y(n_711) );
OAI221xp5_ASAP7_75t_SL g643 ( .A1(n_639), .A2(n_644), .B1(n_648), .B2(n_651), .C(n_653), .Y(n_643) );
INVx1_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
A2O1A1Ixp33_ASAP7_75t_L g706 ( .A1(n_642), .A2(n_707), .B(n_709), .C(n_711), .Y(n_706) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_645), .A2(n_696), .B1(n_698), .B2(n_700), .C(n_703), .Y(n_695) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
NOR4xp25_ASAP7_75t_L g659 ( .A(n_660), .B(n_685), .C(n_706), .D(n_717), .Y(n_659) );
OAI211xp5_ASAP7_75t_SL g660 ( .A1(n_661), .A2(n_662), .B(n_666), .C(n_680), .Y(n_660) );
INVx1_ASAP7_75t_SL g715 ( .A(n_667), .Y(n_715) );
OR2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
INVx1_ASAP7_75t_SL g678 ( .A(n_676), .Y(n_678) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_683), .A2(n_692), .B1(n_704), .B2(n_705), .Y(n_703) );
A2O1A1Ixp33_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_688), .B(n_690), .C(n_695), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AOI31xp33_ASAP7_75t_L g717 ( .A1(n_688), .A2(n_718), .A3(n_720), .B(n_721), .Y(n_717) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVxp67_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
OR2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B(n_716), .Y(n_713) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_724), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_740), .Y(n_739) );
INVx5_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
CKINVDCx9p33_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_742), .Y(n_750) );
OR2x4_ASAP7_75t_L g742 ( .A(n_743), .B(n_745), .Y(n_742) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
endmodule