module fake_jpeg_16447_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

AND2x4_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_0),
.Y(n_34)
);

OR2x2_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_38),
.Y(n_49)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_18),
.B1(n_25),
.B2(n_30),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_45),
.B1(n_15),
.B2(n_23),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_18),
.B1(n_25),
.B2(n_30),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_18),
.B1(n_30),
.B2(n_25),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_46),
.A2(n_50),
.B1(n_51),
.B2(n_35),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_18),
.B1(n_30),
.B2(n_25),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_25),
.B1(n_26),
.B2(n_23),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_58),
.B(n_74),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_50),
.A2(n_34),
.B1(n_40),
.B2(n_26),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_59),
.A2(n_62),
.B1(n_69),
.B2(n_70),
.Y(n_94)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_60),
.A2(n_84),
.B1(n_87),
.B2(n_16),
.Y(n_106)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_36),
.B1(n_23),
.B2(n_26),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_63),
.B(n_73),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_32),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_64),
.B(n_78),
.Y(n_111)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_76),
.Y(n_100)
);

AO22x1_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_40),
.B1(n_32),
.B2(n_41),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_67),
.A2(n_68),
.B1(n_72),
.B2(n_81),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_36),
.B1(n_23),
.B2(n_26),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_23),
.B1(n_26),
.B2(n_15),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_40),
.B1(n_15),
.B2(n_35),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_54),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_42),
.B(n_33),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_49),
.B(n_40),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_77),
.A2(n_24),
.B(n_22),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_32),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_32),
.C(n_37),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_32),
.C(n_77),
.Y(n_107)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_47),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_52),
.A2(n_40),
.B1(n_35),
.B2(n_20),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_85),
.B1(n_88),
.B2(n_24),
.Y(n_113)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_43),
.A2(n_20),
.B1(n_29),
.B2(n_28),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_43),
.A2(n_41),
.B1(n_19),
.B2(n_27),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_43),
.A2(n_20),
.B1(n_29),
.B2(n_28),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_43),
.A2(n_19),
.B1(n_29),
.B2(n_28),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_77),
.A2(n_64),
.B(n_78),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_89),
.A2(n_31),
.B(n_19),
.C(n_80),
.Y(n_131)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_57),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_91),
.B(n_92),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_79),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_93),
.Y(n_126)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_38),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_107),
.C(n_115),
.Y(n_120)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_58),
.B(n_17),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_104),
.B(n_105),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_74),
.B(n_16),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_113),
.B1(n_22),
.B2(n_71),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_67),
.A2(n_41),
.B1(n_37),
.B2(n_47),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_76),
.B1(n_83),
.B2(n_86),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_37),
.C(n_53),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_53),
.C(n_19),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_80),
.C(n_76),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_67),
.A2(n_24),
.B1(n_22),
.B2(n_16),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_0),
.B(n_2),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_117),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_128),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_122),
.B(n_110),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_112),
.A2(n_67),
.B1(n_63),
.B2(n_60),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_136),
.B1(n_137),
.B2(n_141),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_85),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_125),
.A2(n_131),
.B(n_103),
.Y(n_176)
);

INVxp33_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_73),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_147),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_144),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_93),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_134),
.B(n_145),
.Y(n_157)
);

NAND3xp33_ASAP7_75t_SL g135 ( 
.A(n_113),
.B(n_71),
.C(n_10),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_135),
.B(n_141),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_66),
.B1(n_17),
.B2(n_31),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_114),
.A2(n_98),
.B1(n_119),
.B2(n_94),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_139),
.B(n_114),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_66),
.B1(n_8),
.B2(n_9),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_143),
.B(n_146),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_89),
.B(n_17),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_90),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_17),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_2),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_148),
.Y(n_188)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

INVxp33_ASAP7_75t_L g210 ( 
.A(n_152),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_153),
.A2(n_176),
.B(n_178),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_147),
.B(n_98),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_163),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_157),
.Y(n_196)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_158),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_124),
.A2(n_121),
.B1(n_127),
.B2(n_136),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_159),
.A2(n_168),
.B1(n_131),
.B2(n_108),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_161),
.B(n_162),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_97),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_115),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_99),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_165),
.Y(n_185)
);

NOR3xp33_ASAP7_75t_SL g165 ( 
.A(n_140),
.B(n_127),
.C(n_143),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_166),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_169),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_120),
.A2(n_114),
.B1(n_99),
.B2(n_96),
.Y(n_168)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_110),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_171),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_120),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_103),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_172),
.B(n_179),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_173),
.A2(n_132),
.B1(n_131),
.B2(n_137),
.Y(n_181)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_174),
.Y(n_190)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_131),
.Y(n_177)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_109),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_187),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_160),
.C(n_163),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_198),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_151),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_153),
.A2(n_108),
.B1(n_109),
.B2(n_118),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_189),
.A2(n_195),
.B1(n_205),
.B2(n_161),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_173),
.A2(n_118),
.B1(n_17),
.B2(n_31),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_175),
.A2(n_31),
.B1(n_17),
.B2(n_4),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_197),
.A2(n_200),
.B1(n_201),
.B2(n_177),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_31),
.C(n_17),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_158),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_169),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_178),
.A2(n_13),
.B1(n_10),
.B2(n_9),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_178),
.A2(n_13),
.B1(n_10),
.B2(n_9),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_154),
.B(n_31),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_206),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_177),
.A2(n_8),
.B1(n_3),
.B2(n_4),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_154),
.B(n_164),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_8),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_209),
.B(n_156),
.Y(n_224)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_211),
.Y(n_250)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_213),
.B(n_214),
.Y(n_241)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_186),
.A2(n_165),
.B1(n_159),
.B2(n_150),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_218),
.A2(n_219),
.B(n_227),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_208),
.A2(n_185),
.B(n_206),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_231),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_221),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_155),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_223),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_230),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_170),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_226),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_168),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_185),
.A2(n_176),
.B(n_150),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_196),
.A2(n_183),
.B1(n_191),
.B2(n_180),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_228),
.A2(n_234),
.B1(n_210),
.B2(n_3),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_208),
.A2(n_148),
.B(n_174),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_229),
.A2(n_233),
.B(n_201),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_156),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_180),
.B(n_166),
.Y(n_231)
);

XNOR2x1_ASAP7_75t_L g232 ( 
.A(n_182),
.B(n_167),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_232),
.A2(n_203),
.B1(n_194),
.B2(n_198),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_184),
.A2(n_7),
.B(n_3),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_193),
.Y(n_234)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_227),
.A2(n_200),
.B(n_187),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_238),
.A2(n_240),
.B1(n_245),
.B2(n_229),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_217),
.A2(n_203),
.B1(n_191),
.B2(n_192),
.Y(n_240)
);

FAx1_ASAP7_75t_SL g243 ( 
.A(n_225),
.B(n_202),
.CI(n_192),
.CON(n_243),
.SN(n_243)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_243),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_249),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_226),
.A2(n_232),
.B1(n_231),
.B2(n_220),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_209),
.C(n_197),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_224),
.C(n_222),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_233),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_210),
.Y(n_249)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_253),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_268),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_219),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_257),
.C(n_259),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_222),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_251),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_218),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_260),
.A2(n_264),
.B1(n_236),
.B2(n_240),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_250),
.A2(n_211),
.B(n_215),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_261),
.A2(n_237),
.B(n_6),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_230),
.C(n_212),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_263),
.C(n_243),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_223),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_238),
.A2(n_213),
.B1(n_3),
.B2(n_5),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_242),
.B(n_246),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_244),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_241),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_239),
.B(n_2),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_269),
.Y(n_283)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_265),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_279),
.C(n_280),
.Y(n_294)
);

INVxp33_ASAP7_75t_L g277 ( 
.A(n_264),
.Y(n_277)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_262),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_284),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_250),
.C(n_243),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_253),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_281),
.B(n_272),
.Y(n_289)
);

AOI21x1_ASAP7_75t_L g282 ( 
.A1(n_259),
.A2(n_247),
.B(n_252),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_282),
.A2(n_270),
.B(n_257),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_281),
.Y(n_285)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_265),
.Y(n_286)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_274),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_279),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_295),
.Y(n_301)
);

OAI21xp33_ASAP7_75t_L g296 ( 
.A1(n_293),
.A2(n_278),
.B(n_273),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_263),
.Y(n_295)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_296),
.Y(n_306)
);

AOI31xp67_ASAP7_75t_L g297 ( 
.A1(n_285),
.A2(n_283),
.A3(n_275),
.B(n_274),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_299),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_298),
.A2(n_304),
.B(n_286),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_291),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_258),
.B(n_256),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_302),
.A2(n_287),
.B(n_288),
.Y(n_305)
);

AOI21x1_ASAP7_75t_SL g312 ( 
.A1(n_305),
.A2(n_309),
.B(n_7),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_308),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_294),
.C(n_290),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_300),
.A2(n_5),
.B1(n_7),
.B2(n_303),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_5),
.Y(n_310)
);

NAND2xp33_ASAP7_75t_R g313 ( 
.A(n_310),
.B(n_7),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_312),
.A2(n_306),
.B(n_311),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_313),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_315),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_314),
.B1(n_308),
.B2(n_316),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_309),
.Y(n_319)
);


endmodule