module real_jpeg_28793_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_343, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_342, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_343;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_342;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_0),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_0),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_0),
.A2(n_27),
.B1(n_56),
.B2(n_57),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_0),
.A2(n_27),
.B1(n_62),
.B2(n_63),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_1),
.Y(n_116)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_1),
.Y(n_119)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_1),
.Y(n_208)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_3),
.A2(n_37),
.B1(n_62),
.B2(n_63),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_3),
.A2(n_37),
.B1(n_56),
.B2(n_57),
.Y(n_158)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_5),
.Y(n_108)
);

AOI21xp33_ASAP7_75t_SL g113 ( 
.A1(n_5),
.A2(n_29),
.B(n_33),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_5),
.B(n_31),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_5),
.A2(n_62),
.B(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_5),
.B(n_62),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_5),
.B(n_74),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_5),
.A2(n_136),
.B1(n_204),
.B2(n_208),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_5),
.A2(n_32),
.B(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_6),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_110),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_6),
.A2(n_62),
.B1(n_63),
.B2(n_110),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_6),
.A2(n_56),
.B1(n_57),
.B2(n_110),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_8),
.A2(n_49),
.B1(n_56),
.B2(n_57),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_8),
.A2(n_49),
.B1(n_62),
.B2(n_63),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_49),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_9),
.A2(n_62),
.B1(n_63),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_9),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_101),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_9),
.A2(n_56),
.B1(n_57),
.B2(n_101),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_101),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_10),
.A2(n_62),
.B1(n_63),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_10),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_10),
.A2(n_56),
.B1(n_57),
.B2(n_104),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_104),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_104),
.Y(n_290)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_12),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_96),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_12),
.A2(n_56),
.B1(n_57),
.B2(n_96),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_12),
.A2(n_62),
.B1(n_63),
.B2(n_96),
.Y(n_224)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_14),
.A2(n_62),
.B1(n_63),
.B2(n_70),
.Y(n_72)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_14),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_15),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_94),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_15),
.A2(n_62),
.B1(n_63),
.B2(n_94),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_15),
.A2(n_56),
.B1(n_57),
.B2(n_94),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_16),
.A2(n_25),
.B1(n_26),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_16),
.A2(n_51),
.B1(n_56),
.B2(n_57),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_16),
.A2(n_51),
.B1(n_62),
.B2(n_63),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_51),
.Y(n_282)
);

INVx11_ASAP7_75t_SL g59 ( 
.A(n_17),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_38),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_22),
.B(n_43),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_24),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_25),
.B(n_29),
.Y(n_30)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_26),
.A2(n_35),
.B(n_108),
.C(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_31),
.B(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_28),
.A2(n_31),
.B1(n_47),
.B2(n_50),
.Y(n_46)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_28),
.A2(n_31),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_28),
.A2(n_31),
.B1(n_146),
.B2(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_28),
.A2(n_31),
.B1(n_165),
.B2(n_262),
.Y(n_261)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_31),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_32),
.A2(n_69),
.B(n_71),
.C(n_72),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_32),
.B(n_69),
.Y(n_71)
);

OAI32xp33_ASAP7_75t_L g228 ( 
.A1(n_32),
.A2(n_63),
.A3(n_221),
.B1(n_229),
.B2(n_231),
.Y(n_228)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_33),
.B(n_108),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_82),
.B(n_338),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_75),
.C(n_77),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_44),
.A2(n_45),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_52),
.C(n_65),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_46),
.B(n_322),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_48),
.A2(n_79),
.B1(n_81),
.B2(n_290),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_52),
.A2(n_313),
.B1(n_315),
.B2(n_316),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_52),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_52),
.A2(n_65),
.B1(n_316),
.B2(n_323),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_60),
.B(n_64),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_53),
.B(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_53),
.A2(n_60),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_53),
.A2(n_60),
.B1(n_134),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_53),
.A2(n_60),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_53),
.A2(n_60),
.B1(n_179),
.B2(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_53),
.B(n_108),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_53),
.A2(n_60),
.B1(n_100),
.B2(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_53),
.A2(n_60),
.B1(n_64),
.B2(n_271),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_54),
.A2(n_55),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_54),
.A2(n_57),
.A3(n_62),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_55),
.B(n_56),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_56),
.B(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_56),
.B(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_62),
.B(n_232),
.Y(n_231)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_65),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_73),
.B2(n_74),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_66),
.A2(n_67),
.B1(n_74),
.B2(n_314),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_67),
.A2(n_74),
.B1(n_93),
.B2(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_67),
.A2(n_74),
.B1(n_149),
.B2(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_67),
.A2(n_74),
.B1(n_167),
.B2(n_264),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_72),
.B(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_72),
.B1(n_92),
.B2(n_95),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_68),
.A2(n_72),
.B1(n_95),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_68),
.A2(n_72),
.B1(n_125),
.B2(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_68),
.A2(n_72),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_73),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_75),
.A2(n_77),
.B1(n_78),
.B2(n_336),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_75),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_79),
.A2(n_81),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_79),
.A2(n_81),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_331),
.B(n_337),
.Y(n_82)
);

OAI321xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_307),
.A3(n_326),
.B1(n_329),
.B2(n_330),
.C(n_342),
.Y(n_83)
);

AOI321xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_258),
.A3(n_296),
.B1(n_301),
.B2(n_306),
.C(n_343),
.Y(n_84)
);

NOR3xp33_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_151),
.C(n_169),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_129),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_87),
.B(n_129),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_111),
.C(n_121),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_88),
.B(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_106),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_97),
.B2(n_98),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_98),
.C(n_106),
.Y(n_140)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_102),
.A2(n_105),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_102),
.A2(n_105),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_108),
.B(n_119),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_109),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_111),
.A2(n_121),
.B1(n_122),
.B2(n_256),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_111),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_114),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_115),
.A2(n_117),
.B1(n_118),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_115),
.A2(n_118),
.B1(n_197),
.B2(n_199),
.Y(n_196)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

INVx5_ASAP7_75t_SL g274 ( 
.A(n_118),
.Y(n_274)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.C(n_128),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_123),
.B(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_126),
.B(n_128),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_127),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_141),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_140),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_140),
.C(n_141),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_135),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_138),
.B1(n_139),
.B2(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_136),
.A2(n_138),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_136),
.A2(n_138),
.B1(n_198),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_136),
.A2(n_138),
.B1(n_193),
.B2(n_234),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_136),
.A2(n_158),
.B(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_150),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_147),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_147),
.C(n_150),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_L g302 ( 
.A1(n_152),
.A2(n_303),
.B(n_304),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_153),
.B(n_154),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_168),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_161),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_156),
.B(n_161),
.C(n_168),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_157),
.B(n_159),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_160),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_162),
.B(n_164),
.C(n_166),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_252),
.B(n_257),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_238),
.B(n_251),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_214),
.B(n_237),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_194),
.B(n_213),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_184),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_174),
.B(n_184),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_180),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_175),
.A2(n_176),
.B1(n_180),
.B2(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_178),
.Y(n_182)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_191),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_189),
.C(n_191),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_190),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_192),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_201),
.B(n_212),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_200),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_196),
.B(n_200),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_206),
.B(n_211),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_203),
.B(n_205),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_215),
.B(n_216),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_227),
.B1(n_235),
.B2(n_236),
.Y(n_216)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_217),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_222),
.B1(n_225),
.B2(n_226),
.Y(n_217)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_218),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_222),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_226),
.C(n_236),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_224),
.Y(n_248)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_227),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_233),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_233),
.Y(n_246)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_229),
.Y(n_232)
);

INVx8_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_239),
.B(n_240),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_244),
.B2(n_245),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_247),
.C(n_249),
.Y(n_253)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_249),
.B2(n_250),
.Y(n_245)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_246),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_247),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_253),
.B(n_254),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_276),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_259),
.B(n_276),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_266),
.C(n_275),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_260),
.B(n_266),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g340 ( 
.A(n_260),
.Y(n_340)
);

FAx1_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_263),
.CI(n_265),
.CON(n_260),
.SN(n_260)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_261),
.B(n_263),
.C(n_265),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_262),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_264),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_272),
.B2(n_273),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_267),
.B(n_273),
.Y(n_292)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_272),
.A2(n_273),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_272),
.A2(n_288),
.B(n_291),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_300),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_294),
.B2(n_295),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_285),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_279),
.B(n_285),
.C(n_295),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_283),
.B(n_284),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_283),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_282),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_309),
.C(n_318),
.Y(n_308)
);

FAx1_ASAP7_75t_SL g328 ( 
.A(n_284),
.B(n_309),
.CI(n_318),
.CON(n_328),
.SN(n_328)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_285)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_286),
.Y(n_293)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_294),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_297),
.A2(n_302),
.B(n_305),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_298),
.B(n_299),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_319),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_319),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_312),
.B2(n_317),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_310),
.A2(n_311),
.B1(n_321),
.B2(n_324),
.Y(n_320)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_313),
.C(n_316),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_311),
.B(n_324),
.C(n_325),
.Y(n_332)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_312),
.Y(n_317)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_313),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_325),
.Y(n_319)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_321),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_327),
.B(n_328),
.Y(n_329)
);

BUFx24_ASAP7_75t_SL g341 ( 
.A(n_328),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_333),
.Y(n_337)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);


endmodule