module real_jpeg_116_n_16 (n_5, n_4, n_8, n_0, n_12, n_327, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_327;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_1),
.A2(n_30),
.B1(n_37),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_1),
.A2(n_40),
.B1(n_46),
.B2(n_47),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_1),
.A2(n_40),
.B1(n_64),
.B2(n_66),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_1),
.A2(n_40),
.B1(n_59),
.B2(n_60),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_2),
.A2(n_30),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_2),
.A2(n_36),
.B1(n_46),
.B2(n_47),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_2),
.A2(n_36),
.B1(n_64),
.B2(n_66),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_2),
.A2(n_36),
.B1(n_59),
.B2(n_60),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_3),
.A2(n_59),
.B1(n_60),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_68),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_3),
.A2(n_30),
.B1(n_37),
.B2(n_68),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_3),
.A2(n_64),
.B1(n_66),
.B2(n_68),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_5),
.A2(n_59),
.B1(n_60),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_5),
.A2(n_64),
.B1(n_66),
.B2(n_70),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_5),
.A2(n_30),
.B1(n_37),
.B2(n_70),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_5),
.A2(n_46),
.B1(n_47),
.B2(n_70),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_6),
.A2(n_59),
.B1(n_60),
.B2(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_6),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_6),
.A2(n_46),
.B1(n_47),
.B2(n_110),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_6),
.A2(n_30),
.B1(n_37),
.B2(n_110),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_6),
.A2(n_64),
.B1(n_66),
.B2(n_110),
.Y(n_192)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_11),
.A2(n_64),
.B1(n_66),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_11),
.A2(n_30),
.B1(n_37),
.B2(n_73),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_11),
.A2(n_59),
.B1(n_60),
.B2(n_73),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_73),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_12),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_12),
.B(n_30),
.C(n_44),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_12),
.A2(n_46),
.B1(n_47),
.B2(n_99),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_12),
.B(n_33),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_12),
.B(n_120),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_12),
.B(n_66),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_12),
.A2(n_66),
.B(n_183),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_12),
.B(n_127),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_12),
.A2(n_59),
.B(n_221),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_45)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_14),
.A2(n_30),
.B1(n_37),
.B2(n_49),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_14),
.A2(n_49),
.B1(n_64),
.B2(n_66),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_14),
.A2(n_49),
.B1(n_59),
.B2(n_60),
.Y(n_278)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_319),
.C(n_324),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_317),
.B(n_321),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_307),
.B(n_316),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_273),
.B(n_304),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_250),
.B(n_272),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_136),
.B(n_249),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_111),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_23),
.B(n_111),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_83),
.C(n_94),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_24),
.B(n_83),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_54),
.B2(n_55),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_25),
.B(n_56),
.C(n_71),
.Y(n_112)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_41),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_27),
.B(n_41),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_34),
.B(n_38),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_28),
.A2(n_32),
.B(n_87),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_28),
.A2(n_32),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_28),
.A2(n_38),
.B(n_87),
.Y(n_185)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_29),
.B(n_39),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_29),
.A2(n_33),
.B1(n_35),
.B2(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_29),
.A2(n_86),
.B(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_29),
.A2(n_33),
.B1(n_99),
.B2(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_29),
.A2(n_33),
.B1(n_163),
.B2(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_37),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_30),
.B(n_161),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_32),
.B(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_32),
.A2(n_89),
.B(n_103),
.Y(n_211)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_33),
.B(n_39),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_45),
.B(n_50),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_42),
.A2(n_45),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_42),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_42),
.A2(n_92),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_42),
.B(n_200),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_53)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OA22x2_ASAP7_75t_SL g79 ( 
.A1(n_46),
.A2(n_47),
.B1(n_76),
.B2(n_78),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_46),
.B(n_78),
.Y(n_184)
);

CKINVDCx6p67_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_47),
.B(n_153),
.Y(n_152)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_47),
.A2(n_66),
.A3(n_76),
.B1(n_182),
.B2(n_184),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_50),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_51),
.B(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_52),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_52),
.A2(n_120),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_52),
.A2(n_120),
.B1(n_148),
.B2(n_156),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_52),
.A2(n_198),
.B(n_199),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_52),
.A2(n_120),
.B(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_71),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_63),
.B1(n_67),
.B2(n_69),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_57),
.A2(n_63),
.B1(n_67),
.B2(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_57),
.A2(n_69),
.B(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_57),
.A2(n_63),
.B1(n_109),
.B2(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_57),
.A2(n_260),
.B(n_261),
.Y(n_259)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_57),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_57),
.A2(n_63),
.B1(n_278),
.B2(n_288),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_57),
.A2(n_261),
.B(n_288),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_63),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_99),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_62),
.C(n_66),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_61),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_66),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_64),
.B(n_98),
.C(n_100),
.Y(n_97)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_63),
.A2(n_278),
.B(n_279),
.Y(n_277)
);

CKINVDCx6p67_ASAP7_75t_R g66 ( 
.A(n_64),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_66),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_74),
.B(n_80),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_72),
.A2(n_74),
.B(n_79),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_105),
.B(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_74),
.A2(n_79),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_74),
.A2(n_79),
.B1(n_105),
.B2(n_206),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_79),
.A2(n_130),
.B(n_131),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_79),
.B(n_99),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_80),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_81),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_82),
.B(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_82),
.A2(n_132),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_82),
.A2(n_132),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_90),
.B2(n_91),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_84),
.B(n_91),
.Y(n_133)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

INVxp33_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_92),
.A2(n_93),
.B(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_92),
.A2(n_119),
.B(n_200),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_94),
.B(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_104),
.C(n_108),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_95),
.B(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_101),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_96),
.A2(n_97),
.B1(n_101),
.B2(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_98),
.Y(n_221)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_101),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_104),
.B(n_108),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_106),
.B(n_131),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_135),
.Y(n_111)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_122),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_115),
.B(n_122),
.C(n_135),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_121),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_116),
.A2(n_117),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_117),
.B(n_118),
.Y(n_263)
);

AOI21xp33_ASAP7_75t_L g300 ( 
.A1(n_117),
.A2(n_258),
.B(n_263),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_118),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_133),
.B2(n_134),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_129),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_125),
.B(n_129),
.C(n_134),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_126),
.B(n_279),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_127),
.B(n_262),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_127),
.A2(n_128),
.B(n_280),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_128),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_130),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_132),
.A2(n_269),
.B(n_282),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_133),
.Y(n_134)
);

AOI321xp33_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_231),
.A3(n_241),
.B1(n_247),
.B2(n_248),
.C(n_327),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_214),
.B(n_230),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_194),
.B(n_213),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_176),
.B(n_193),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_157),
.B(n_175),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_150),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_150),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_147),
.C(n_178),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_144),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_149),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_151),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_169),
.B(n_174),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_164),
.B(n_168),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_167),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_173),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_179),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_186),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_187),
.C(n_190),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_185),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_185),
.Y(n_201)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_192),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_212),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_212),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_202),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_201),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_201),
.C(n_202),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_199),
.B(n_266),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_200),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_207),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_209),
.C(n_210),
.Y(n_227)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_216),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_225),
.B2(n_226),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_227),
.C(n_228),
.Y(n_242)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_222),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_223),
.C(n_224),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_234),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_238),
.C(n_240),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_235),
.A2(n_236),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_240),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_243),
.Y(n_247)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_271),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_271),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_252),
.B(n_256),
.C(n_264),
.Y(n_302)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_264),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_263),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_262),
.B(n_280),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_267),
.B(n_270),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_267),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_296),
.C(n_300),
.Y(n_295)
);

FAx1_ASAP7_75t_SL g303 ( 
.A(n_270),
.B(n_296),
.CI(n_300),
.CON(n_303),
.SN(n_303)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_301),
.Y(n_273)
);

AOI21xp33_ASAP7_75t_L g304 ( 
.A1(n_274),
.A2(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_295),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_275),
.B(n_295),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_285),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_276),
.B(n_277),
.C(n_294),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_281),
.C(n_283),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_277),
.A2(n_286),
.B1(n_293),
.B2(n_294),
.Y(n_285)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_277),
.A2(n_293),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_281),
.A2(n_283),
.B1(n_292),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_281),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_283),
.A2(n_290),
.B1(n_291),
.B2(n_292),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_283),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_283),
.B(n_287),
.C(n_291),
.Y(n_315)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_286),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_303),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g325 ( 
.A(n_303),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_309),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_315),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B1(n_313),
.B2(n_314),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_313),
.C(n_315),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_314),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_320),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_320),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);


endmodule