module fake_jpeg_22208_n_287 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_287);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_287;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx8_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_13),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_42),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_23),
.C(n_27),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_45),
.B(n_18),
.Y(n_77)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_29),
.B1(n_26),
.B2(n_15),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_58),
.B1(n_18),
.B2(n_15),
.Y(n_78)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_55),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_32),
.A2(n_20),
.B1(n_27),
.B2(n_18),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_29),
.B1(n_26),
.B2(n_22),
.Y(n_70)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_37),
.B(n_21),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_56),
.B(n_57),
.Y(n_68)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_59),
.B(n_21),
.Y(n_73)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_64),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_39),
.B1(n_34),
.B2(n_33),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_57),
.B1(n_53),
.B2(n_28),
.Y(n_84)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_29),
.B1(n_26),
.B2(n_20),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_66),
.A2(n_69),
.B1(n_54),
.B2(n_28),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

AO22x1_ASAP7_75t_SL g69 ( 
.A1(n_54),
.A2(n_38),
.B1(n_20),
.B2(n_27),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_76),
.B1(n_28),
.B2(n_18),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_44),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_59),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_56),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_22),
.B1(n_31),
.B2(n_15),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_55),
.C(n_43),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_42),
.B1(n_19),
.B2(n_17),
.Y(n_94)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_84),
.A2(n_86),
.B1(n_76),
.B2(n_63),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_88),
.B(n_91),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_95),
.Y(n_112)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_53),
.B1(n_54),
.B2(n_22),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_92),
.A2(n_66),
.B1(n_69),
.B2(n_65),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_102),
.B1(n_67),
.B2(n_80),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_SL g127 ( 
.A(n_94),
.B(n_96),
.C(n_97),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_43),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_25),
.B(n_16),
.C(n_46),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_69),
.A2(n_72),
.B1(n_67),
.B2(n_42),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_41),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_68),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_69),
.A2(n_48),
.B1(n_46),
.B2(n_24),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_68),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_104),
.B(n_106),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_82),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_105),
.Y(n_131)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_107),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_109),
.B(n_110),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_SL g113 ( 
.A1(n_102),
.A2(n_77),
.B(n_60),
.C(n_64),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_51),
.B(n_80),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_79),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_82),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_115),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_116),
.A2(n_124),
.B1(n_125),
.B2(n_83),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_99),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_117),
.Y(n_146)
);

MAJx2_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_90),
.C(n_89),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_96),
.C(n_71),
.Y(n_135)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_87),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_103),
.B(n_89),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_121),
.A2(n_119),
.B(n_108),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_98),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_122),
.Y(n_143)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_67),
.B1(n_81),
.B2(n_79),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_92),
.A2(n_71),
.B1(n_19),
.B2(n_21),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_126),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_145),
.B1(n_105),
.B2(n_115),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_127),
.A2(n_88),
.B1(n_87),
.B2(n_86),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_130),
.A2(n_134),
.B(n_142),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_121),
.C(n_120),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_107),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_136),
.B(n_126),
.Y(n_161)
);

OAI32xp33_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_110),
.A3(n_125),
.B1(n_122),
.B2(n_61),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_84),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_151),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_83),
.Y(n_140)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_127),
.A2(n_80),
.B(n_99),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_116),
.A2(n_24),
.B1(n_19),
.B2(n_51),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_124),
.B1(n_113),
.B2(n_106),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_51),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_113),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_0),
.Y(n_151)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_153),
.A2(n_173),
.B1(n_136),
.B2(n_133),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_156),
.C(n_166),
.Y(n_179)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_158),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_118),
.C(n_113),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_157),
.B(n_171),
.Y(n_188)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_167),
.B(n_175),
.Y(n_187)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_169),
.Y(n_186)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_161),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_109),
.Y(n_163)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_164),
.A2(n_165),
.B1(n_137),
.B2(n_25),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_129),
.C(n_145),
.Y(n_166)
);

AND2x2_ASAP7_75t_SL g167 ( 
.A(n_131),
.B(n_123),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_122),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_139),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_61),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_131),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_170),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_13),
.C(n_2),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_141),
.B(n_130),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_172),
.Y(n_199)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_174),
.A2(n_141),
.B1(n_146),
.B2(n_150),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_1),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_185),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_149),
.C(n_148),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_189),
.C(n_194),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_182),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_156),
.B(n_148),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_166),
.C(n_154),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_148),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_196),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_191),
.Y(n_200)
);

OAI22x1_ASAP7_75t_L g209 ( 
.A1(n_192),
.A2(n_167),
.B1(n_153),
.B2(n_169),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_162),
.A2(n_149),
.B(n_147),
.C(n_138),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_193),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_146),
.C(n_133),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_144),
.B1(n_143),
.B2(n_137),
.Y(n_195)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_143),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_197),
.A2(n_173),
.B1(n_152),
.B2(n_155),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_16),
.B1(n_2),
.B2(n_3),
.Y(n_198)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_185),
.B(n_159),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_205),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_163),
.Y(n_204)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_159),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_200),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_191),
.A2(n_152),
.B1(n_160),
.B2(n_165),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_1),
.Y(n_212)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_1),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_214),
.Y(n_233)
);

NOR2x1_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_2),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_215),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_3),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_217),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_194),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_202),
.A2(n_177),
.B1(n_190),
.B2(n_192),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_222),
.A2(n_230),
.B1(n_207),
.B2(n_218),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_189),
.C(n_179),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_231),
.C(n_232),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_196),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_228),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_215),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_227),
.A2(n_219),
.B(n_221),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_181),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_179),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_211),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_206),
.A2(n_188),
.B1(n_193),
.B2(n_195),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_187),
.C(n_198),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_187),
.C(n_4),
.Y(n_232)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_234),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_3),
.Y(n_235)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_222),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_238),
.B(n_229),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_231),
.A2(n_209),
.B(n_213),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_243),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_220),
.A2(n_208),
.B1(n_232),
.B2(n_204),
.Y(n_241)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_211),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_224),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_233),
.A2(n_214),
.B1(n_203),
.B2(n_7),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_6),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_4),
.C(n_6),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_248),
.C(n_226),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_4),
.C(n_6),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_240),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_251),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_255),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_247),
.B(n_225),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_258),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_4),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_240),
.C(n_239),
.Y(n_266)
);

AOI21xp33_ASAP7_75t_L g260 ( 
.A1(n_246),
.A2(n_12),
.B(n_7),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_260),
.A2(n_249),
.B(n_8),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_6),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_248),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_259),
.A2(n_237),
.B(n_241),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_262),
.A2(n_266),
.B(n_268),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_261),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_265),
.B(n_9),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_7),
.B(n_9),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_251),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_270),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_262),
.Y(n_272)
);

AO21x1_ASAP7_75t_L g277 ( 
.A1(n_272),
.A2(n_273),
.B(n_275),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_264),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_266),
.C(n_257),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_276),
.Y(n_278)
);

AO21x1_ASAP7_75t_L g282 ( 
.A1(n_278),
.A2(n_279),
.B(n_280),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_267),
.Y(n_280)
);

AOI21xp33_ASAP7_75t_L g281 ( 
.A1(n_277),
.A2(n_269),
.B(n_267),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_281),
.A2(n_282),
.B(n_252),
.Y(n_283)
);

NAND3xp33_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_252),
.C(n_253),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_9),
.C(n_10),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_11),
.Y(n_286)
);

AOI321xp33_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_11),
.A3(n_12),
.B1(n_235),
.B2(n_275),
.C(n_215),
.Y(n_287)
);


endmodule