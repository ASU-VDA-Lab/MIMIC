module fake_ariane_356_n_903 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_903);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_903;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_819;
wire n_717;
wire n_706;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_320;
wire n_331;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_840;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_795;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_218;
wire n_839;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_365;
wire n_238;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_889;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_705;
wire n_630;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_772;
wire n_747;
wire n_847;
wire n_371;
wire n_845;
wire n_888;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_856;
wire n_782;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

INVx2_ASAP7_75t_L g200 ( 
.A(n_97),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_110),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_192),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_92),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_107),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_35),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_42),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_82),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_143),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_90),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_158),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_71),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_33),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_12),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_193),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_172),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_51),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_16),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_185),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_83),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_127),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_147),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_195),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_154),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_186),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_68),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_45),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_168),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_160),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_6),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_58),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_113),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_102),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_165),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_84),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_132),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_194),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_91),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_78),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_136),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_81),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_76),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_162),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_109),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_101),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_99),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_183),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_123),
.Y(n_248)
);

INVxp67_ASAP7_75t_SL g249 ( 
.A(n_2),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_88),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_177),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_116),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_86),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_16),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_133),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_5),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_163),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_50),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_139),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_12),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_191),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_189),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_198),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_2),
.Y(n_264)
);

BUFx8_ASAP7_75t_SL g265 ( 
.A(n_155),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_128),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_72),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_1),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_187),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_57),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_156),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_138),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_13),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_21),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_53),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_175),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_197),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_61),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_135),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_52),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_31),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_54),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_32),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_26),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_190),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_5),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_204),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_206),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_213),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_208),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_216),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_213),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_264),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_218),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_260),
.Y(n_296)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_274),
.Y(n_297)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_274),
.Y(n_298)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_274),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_254),
.Y(n_300)
);

AND2x4_ASAP7_75t_L g301 ( 
.A(n_273),
.B(n_0),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_231),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_217),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_230),
.Y(n_304)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_279),
.Y(n_305)
);

XNOR2x2_ASAP7_75t_L g306 ( 
.A(n_207),
.B(n_0),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_200),
.B(n_1),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_249),
.Y(n_308)
);

OA21x2_ASAP7_75t_L g309 ( 
.A1(n_219),
.A2(n_3),
.B(n_4),
.Y(n_309)
);

AOI22x1_ASAP7_75t_SL g310 ( 
.A1(n_227),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_256),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_220),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_279),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_235),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_236),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_286),
.Y(n_317)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_279),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_279),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_240),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_255),
.B(n_7),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_241),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_245),
.B(n_7),
.Y(n_323)
);

AND2x4_ASAP7_75t_L g324 ( 
.A(n_200),
.B(n_8),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_233),
.B(n_8),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_248),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_250),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_253),
.B(n_9),
.Y(n_328)
);

BUFx12f_ASAP7_75t_L g329 ( 
.A(n_201),
.Y(n_329)
);

BUFx8_ASAP7_75t_L g330 ( 
.A(n_233),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_258),
.B(n_9),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_261),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_262),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_255),
.Y(n_334)
);

BUFx8_ASAP7_75t_L g335 ( 
.A(n_266),
.Y(n_335)
);

AND2x4_ASAP7_75t_L g336 ( 
.A(n_272),
.B(n_10),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_280),
.B(n_10),
.Y(n_337)
);

INVx5_ASAP7_75t_L g338 ( 
.A(n_265),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_283),
.B(n_11),
.Y(n_339)
);

OA21x2_ASAP7_75t_L g340 ( 
.A1(n_281),
.A2(n_11),
.B(n_13),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_202),
.Y(n_341)
);

BUFx12f_ASAP7_75t_L g342 ( 
.A(n_203),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_302),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_334),
.B(n_221),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_329),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_315),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_342),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_302),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_338),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_338),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_R g351 ( 
.A(n_334),
.B(n_244),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_295),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_338),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_315),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_338),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_341),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_295),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_341),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_341),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_335),
.Y(n_360)
);

NAND2xp33_ASAP7_75t_R g361 ( 
.A(n_293),
.B(n_205),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_335),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_300),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_330),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_311),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_330),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_311),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_291),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_296),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_317),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_303),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_303),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_295),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_289),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_291),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_304),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_304),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_333),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_313),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_312),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_312),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_321),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_292),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_292),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_333),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_333),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_R g387 ( 
.A(n_320),
.B(n_263),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_287),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_297),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_313),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_313),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_297),
.Y(n_392)
);

BUFx10_ASAP7_75t_L g393 ( 
.A(n_324),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_298),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_R g395 ( 
.A(n_322),
.B(n_285),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_298),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_301),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_326),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_380),
.B(n_339),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_371),
.B(n_332),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_381),
.B(n_336),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_398),
.B(n_336),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_356),
.B(n_324),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_378),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_369),
.B(n_308),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_372),
.B(n_314),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_376),
.B(n_287),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_383),
.B(n_325),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_351),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_374),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_384),
.B(n_325),
.Y(n_411)
);

NOR3xp33_ASAP7_75t_L g412 ( 
.A(n_346),
.B(n_331),
.C(n_323),
.Y(n_412)
);

INVxp33_ASAP7_75t_L g413 ( 
.A(n_387),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_389),
.B(n_288),
.Y(n_414)
);

NAND2xp33_ASAP7_75t_L g415 ( 
.A(n_377),
.B(n_323),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_363),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_373),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_392),
.B(n_288),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_388),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_368),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_393),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_379),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_365),
.B(n_290),
.Y(n_423)
);

NAND3xp33_ASAP7_75t_L g424 ( 
.A(n_367),
.B(n_328),
.C(n_331),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_393),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_385),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_386),
.Y(n_427)
);

NOR2xp67_ASAP7_75t_L g428 ( 
.A(n_390),
.B(n_299),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_391),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_394),
.B(n_290),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_396),
.B(n_397),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_357),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_357),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_352),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_375),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_352),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_358),
.B(n_294),
.Y(n_437)
);

OR2x6_ASAP7_75t_L g438 ( 
.A(n_344),
.B(n_307),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_361),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_352),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_352),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_359),
.B(n_294),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_348),
.B(n_316),
.Y(n_443)
);

OAI22xp33_ASAP7_75t_L g444 ( 
.A1(n_361),
.A2(n_337),
.B1(n_307),
.B2(n_301),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_395),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_349),
.Y(n_446)
);

BUFx6f_ASAP7_75t_SL g447 ( 
.A(n_343),
.Y(n_447)
);

INVxp33_ASAP7_75t_SL g448 ( 
.A(n_345),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_350),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_370),
.B(n_316),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_353),
.B(n_327),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_355),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_364),
.B(n_327),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_366),
.B(n_328),
.Y(n_454)
);

NOR2xp67_ASAP7_75t_L g455 ( 
.A(n_347),
.B(n_299),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_354),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_382),
.B(n_337),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_360),
.B(n_222),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_362),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_380),
.B(n_299),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_378),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_345),
.B(n_225),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_371),
.B(n_232),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_380),
.B(n_299),
.Y(n_464)
);

NAND2xp33_ASAP7_75t_L g465 ( 
.A(n_371),
.B(n_209),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_361),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_374),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_378),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_380),
.B(n_305),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_371),
.B(n_305),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_410),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_444),
.A2(n_340),
.B1(n_309),
.B2(n_310),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_407),
.B(n_309),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_L g474 ( 
.A1(n_438),
.A2(n_306),
.B1(n_340),
.B2(n_319),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_434),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_456),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_412),
.A2(n_247),
.B1(n_211),
.B2(n_212),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_467),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_435),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_443),
.B(n_14),
.Y(n_480)
);

INVx2_ASAP7_75t_SL g481 ( 
.A(n_420),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_416),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_438),
.A2(n_319),
.B1(n_251),
.B2(n_246),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_463),
.B(n_210),
.Y(n_484)
);

NOR3xp33_ASAP7_75t_SL g485 ( 
.A(n_424),
.B(n_215),
.C(n_214),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_400),
.B(n_223),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_419),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_448),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_450),
.B(n_406),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_414),
.B(n_224),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_405),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_423),
.B(n_226),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_404),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_461),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_439),
.B(n_228),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_434),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_466),
.B(n_229),
.Y(n_497)
);

NOR3xp33_ASAP7_75t_SL g498 ( 
.A(n_424),
.B(n_237),
.C(n_234),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_447),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_434),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_449),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_418),
.B(n_238),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_413),
.B(n_14),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_409),
.B(n_15),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_438),
.A2(n_319),
.B1(n_271),
.B2(n_270),
.Y(n_505)
);

BUFx8_ASAP7_75t_L g506 ( 
.A(n_447),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_468),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_433),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_431),
.B(n_239),
.Y(n_509)
);

BUFx8_ASAP7_75t_L g510 ( 
.A(n_459),
.Y(n_510)
);

NOR3xp33_ASAP7_75t_SL g511 ( 
.A(n_454),
.B(n_243),
.C(n_242),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_440),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_430),
.B(n_252),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_432),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_457),
.B(n_15),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_445),
.B(n_257),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_408),
.B(n_259),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_417),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_440),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_440),
.Y(n_520)
);

AND2x2_ASAP7_75t_SL g521 ( 
.A(n_462),
.B(n_267),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_411),
.B(n_269),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_437),
.B(n_275),
.Y(n_523)
);

O2A1O1Ixp5_ASAP7_75t_L g524 ( 
.A1(n_401),
.A2(n_284),
.B(n_282),
.C(n_278),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_422),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_429),
.Y(n_526)
);

NOR2x1_ASAP7_75t_L g527 ( 
.A(n_455),
.B(n_276),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_449),
.B(n_402),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_403),
.A2(n_442),
.B1(n_399),
.B2(n_427),
.Y(n_529)
);

INVx5_ASAP7_75t_L g530 ( 
.A(n_449),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_436),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_441),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_428),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_426),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_421),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_451),
.B(n_277),
.Y(n_536)
);

AND2x4_ASAP7_75t_SL g537 ( 
.A(n_425),
.B(n_17),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_452),
.B(n_305),
.Y(n_538)
);

INVxp67_ASAP7_75t_SL g539 ( 
.A(n_453),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_428),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_446),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_470),
.B(n_305),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_455),
.B(n_318),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_460),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_458),
.B(n_318),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_493),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_522),
.A2(n_517),
.B(n_415),
.Y(n_547)
);

NAND3xp33_ASAP7_75t_SL g548 ( 
.A(n_477),
.B(n_469),
.C(n_464),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_530),
.B(n_465),
.Y(n_549)
);

OAI22x1_ASAP7_75t_L g550 ( 
.A1(n_472),
.A2(n_318),
.B1(n_19),
.B2(n_20),
.Y(n_550)
);

NOR2xp67_ASAP7_75t_SL g551 ( 
.A(n_488),
.B(n_530),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_476),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_530),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_522),
.A2(n_318),
.B(n_22),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_489),
.B(n_18),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_514),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_539),
.B(n_199),
.Y(n_557)
);

INVx5_ASAP7_75t_L g558 ( 
.A(n_541),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_536),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_501),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_509),
.B(n_27),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_506),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_490),
.A2(n_28),
.B(n_29),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_521),
.A2(n_30),
.B1(n_34),
.B2(n_36),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_541),
.B(n_37),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_477),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_566)
);

OR2x6_ASAP7_75t_L g567 ( 
.A(n_481),
.B(n_41),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_491),
.B(n_43),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_502),
.A2(n_44),
.B(n_46),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_513),
.A2(n_47),
.B(n_48),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_526),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_471),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_491),
.B(n_196),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_480),
.B(n_49),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_478),
.Y(n_575)
);

NOR3xp33_ASAP7_75t_SL g576 ( 
.A(n_516),
.B(n_55),
.C(n_56),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_541),
.B(n_59),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_535),
.B(n_60),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_536),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_473),
.A2(n_65),
.B(n_66),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_497),
.B(n_484),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_497),
.B(n_67),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_482),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_515),
.B(n_69),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_492),
.B(n_70),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_494),
.Y(n_586)
);

OAI21xp33_ASAP7_75t_SL g587 ( 
.A1(n_487),
.A2(n_73),
.B(n_74),
.Y(n_587)
);

A2O1A1Ixp33_ASAP7_75t_L g588 ( 
.A1(n_472),
.A2(n_75),
.B(n_77),
.C(n_79),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_499),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_508),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_479),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_534),
.A2(n_80),
.B1(n_85),
.B2(n_87),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_529),
.B(n_523),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_507),
.Y(n_594)
);

AND2x6_ASAP7_75t_L g595 ( 
.A(n_503),
.B(n_89),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_492),
.B(n_93),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_518),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_504),
.B(n_94),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_544),
.B(n_95),
.Y(n_599)
);

NAND2xp33_ASAP7_75t_SL g600 ( 
.A(n_485),
.B(n_96),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_473),
.A2(n_528),
.B(n_486),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_525),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_495),
.B(n_98),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_537),
.Y(n_604)
);

NOR2xp67_ASAP7_75t_L g605 ( 
.A(n_533),
.B(n_100),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_532),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_581),
.B(n_483),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_558),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_558),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_552),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_L g611 ( 
.A1(n_601),
.A2(n_524),
.B(n_531),
.Y(n_611)
);

AO21x2_ASAP7_75t_L g612 ( 
.A1(n_547),
.A2(n_545),
.B(n_498),
.Y(n_612)
);

CKINVDCx11_ASAP7_75t_R g613 ( 
.A(n_589),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_553),
.Y(n_614)
);

NAND2x1p5_ASAP7_75t_L g615 ( 
.A(n_558),
.B(n_553),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_556),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_586),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_594),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_595),
.Y(n_619)
);

OAI21x1_ASAP7_75t_L g620 ( 
.A1(n_580),
.A2(n_531),
.B(n_519),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g621 ( 
.A(n_591),
.Y(n_621)
);

AOI22x1_ASAP7_75t_L g622 ( 
.A1(n_554),
.A2(n_500),
.B1(n_496),
.B2(n_512),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_560),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_560),
.B(n_496),
.Y(n_624)
);

INVx6_ASAP7_75t_SL g625 ( 
.A(n_567),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_595),
.Y(n_626)
);

AOI22x1_ASAP7_75t_L g627 ( 
.A1(n_550),
.A2(n_512),
.B1(n_519),
.B2(n_500),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_595),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_562),
.Y(n_629)
);

OAI21x1_ASAP7_75t_L g630 ( 
.A1(n_563),
.A2(n_527),
.B(n_540),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_604),
.Y(n_631)
);

OAI21x1_ASAP7_75t_L g632 ( 
.A1(n_569),
.A2(n_542),
.B(n_543),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_590),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_572),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_575),
.Y(n_635)
);

OR2x6_ASAP7_75t_L g636 ( 
.A(n_549),
.B(n_475),
.Y(n_636)
);

AO21x2_ASAP7_75t_L g637 ( 
.A1(n_585),
.A2(n_538),
.B(n_511),
.Y(n_637)
);

AO21x2_ASAP7_75t_L g638 ( 
.A1(n_596),
.A2(n_474),
.B(n_475),
.Y(n_638)
);

OAI21x1_ASAP7_75t_L g639 ( 
.A1(n_570),
.A2(n_505),
.B(n_520),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_583),
.Y(n_640)
);

AO21x2_ASAP7_75t_L g641 ( 
.A1(n_574),
.A2(n_520),
.B(n_475),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_606),
.Y(n_642)
);

AO21x2_ASAP7_75t_L g643 ( 
.A1(n_593),
.A2(n_520),
.B(n_104),
.Y(n_643)
);

AO21x2_ASAP7_75t_L g644 ( 
.A1(n_548),
.A2(n_561),
.B(n_584),
.Y(n_644)
);

OAI21x1_ASAP7_75t_L g645 ( 
.A1(n_599),
.A2(n_103),
.B(n_105),
.Y(n_645)
);

INVxp67_ASAP7_75t_SL g646 ( 
.A(n_551),
.Y(n_646)
);

OAI21x1_ASAP7_75t_L g647 ( 
.A1(n_559),
.A2(n_579),
.B(n_555),
.Y(n_647)
);

OAI21x1_ASAP7_75t_L g648 ( 
.A1(n_565),
.A2(n_106),
.B(n_108),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_557),
.A2(n_111),
.B(n_112),
.Y(n_649)
);

BUFx12f_ASAP7_75t_L g650 ( 
.A(n_567),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_L g651 ( 
.A1(n_582),
.A2(n_114),
.B(n_115),
.Y(n_651)
);

OR2x6_ASAP7_75t_L g652 ( 
.A(n_598),
.B(n_506),
.Y(n_652)
);

AOI22x1_ASAP7_75t_L g653 ( 
.A1(n_597),
.A2(n_510),
.B1(n_118),
.B2(n_119),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_617),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_640),
.Y(n_655)
);

OAI22xp33_ASAP7_75t_L g656 ( 
.A1(n_607),
.A2(n_564),
.B1(n_566),
.B2(n_592),
.Y(n_656)
);

BUFx4_ASAP7_75t_SL g657 ( 
.A(n_652),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_617),
.Y(n_658)
);

CKINVDCx8_ASAP7_75t_R g659 ( 
.A(n_652),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_629),
.Y(n_660)
);

BUFx2_ASAP7_75t_R g661 ( 
.A(n_629),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_635),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_618),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_610),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_618),
.Y(n_665)
);

OAI22xp33_ASAP7_75t_L g666 ( 
.A1(n_652),
.A2(n_573),
.B1(n_568),
.B2(n_602),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_624),
.B(n_614),
.Y(n_667)
);

AO21x1_ASAP7_75t_L g668 ( 
.A1(n_649),
.A2(n_600),
.B(n_603),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_SL g669 ( 
.A1(n_650),
.A2(n_510),
.B1(n_578),
.B2(n_587),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_616),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_616),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_634),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_634),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_614),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_642),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_642),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_633),
.Y(n_677)
);

BUFx12f_ASAP7_75t_L g678 ( 
.A(n_613),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_633),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_613),
.Y(n_680)
);

AOI21x1_ASAP7_75t_L g681 ( 
.A1(n_647),
.A2(n_605),
.B(n_577),
.Y(n_681)
);

BUFx12f_ASAP7_75t_L g682 ( 
.A(n_650),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_628),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_SL g684 ( 
.A1(n_628),
.A2(n_588),
.B1(n_546),
.B2(n_571),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_633),
.Y(n_685)
);

AOI21xp33_ASAP7_75t_L g686 ( 
.A1(n_638),
.A2(n_576),
.B(n_120),
.Y(n_686)
);

INVx1_ASAP7_75t_SL g687 ( 
.A(n_621),
.Y(n_687)
);

AO21x1_ASAP7_75t_L g688 ( 
.A1(n_651),
.A2(n_117),
.B(n_121),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_SL g689 ( 
.A1(n_628),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_615),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_623),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_652),
.A2(n_126),
.B1(n_129),
.B2(n_130),
.Y(n_692)
);

OAI21x1_ASAP7_75t_L g693 ( 
.A1(n_620),
.A2(n_622),
.B(n_632),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_666),
.B(n_619),
.Y(n_694)
);

OR2x2_ASAP7_75t_SL g695 ( 
.A(n_657),
.B(n_625),
.Y(n_695)
);

AND2x4_ASAP7_75t_SL g696 ( 
.A(n_667),
.B(n_690),
.Y(n_696)
);

BUFx2_ASAP7_75t_L g697 ( 
.A(n_664),
.Y(n_697)
);

A2O1A1Ixp33_ASAP7_75t_L g698 ( 
.A1(n_669),
.A2(n_647),
.B(n_626),
.C(n_619),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_R g699 ( 
.A(n_667),
.B(n_619),
.Y(n_699)
);

CKINVDCx20_ASAP7_75t_R g700 ( 
.A(n_691),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_656),
.A2(n_626),
.B1(n_646),
.B2(n_636),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_654),
.Y(n_702)
);

NOR3xp33_ASAP7_75t_SL g703 ( 
.A(n_656),
.B(n_611),
.C(n_625),
.Y(n_703)
);

CKINVDCx16_ASAP7_75t_R g704 ( 
.A(n_678),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_687),
.B(n_624),
.Y(n_705)
);

AO31x2_ASAP7_75t_L g706 ( 
.A1(n_688),
.A2(n_643),
.A3(n_644),
.B(n_638),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_672),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_662),
.Y(n_708)
);

OR2x6_ASAP7_75t_L g709 ( 
.A(n_672),
.B(n_626),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_665),
.Y(n_710)
);

NAND2xp33_ASAP7_75t_R g711 ( 
.A(n_683),
.B(n_624),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_658),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_655),
.B(n_615),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_663),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_R g715 ( 
.A(n_683),
.B(n_673),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_671),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_670),
.Y(n_717)
);

NOR2xp67_ASAP7_75t_R g718 ( 
.A(n_657),
.B(n_608),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_676),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_676),
.Y(n_720)
);

NOR3xp33_ASAP7_75t_SL g721 ( 
.A(n_680),
.B(n_625),
.C(n_637),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_687),
.B(n_661),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_661),
.B(n_631),
.Y(n_723)
);

CKINVDCx16_ASAP7_75t_R g724 ( 
.A(n_682),
.Y(n_724)
);

OAI21xp5_ASAP7_75t_L g725 ( 
.A1(n_684),
.A2(n_639),
.B(n_627),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_675),
.B(n_631),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_690),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_685),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_685),
.B(n_644),
.Y(n_729)
);

NAND2xp33_ASAP7_75t_R g730 ( 
.A(n_659),
.B(n_608),
.Y(n_730)
);

BUFx4f_ASAP7_75t_SL g731 ( 
.A(n_660),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_677),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_674),
.B(n_609),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_679),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_690),
.B(n_608),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_669),
.B(n_641),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_692),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_681),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_668),
.B(n_609),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_686),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_693),
.B(n_636),
.Y(n_741)
);

OR2x6_ASAP7_75t_L g742 ( 
.A(n_736),
.B(n_636),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_708),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_729),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_697),
.B(n_684),
.Y(n_745)
);

BUFx2_ASAP7_75t_L g746 ( 
.A(n_707),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_729),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_710),
.Y(n_748)
);

NOR2x1p5_ASAP7_75t_L g749 ( 
.A(n_737),
.B(n_653),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_705),
.B(n_612),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_722),
.B(n_612),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_719),
.B(n_641),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_716),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_720),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_728),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_734),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_723),
.B(n_612),
.Y(n_757)
);

OR2x2_ASAP7_75t_L g758 ( 
.A(n_726),
.B(n_636),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_694),
.A2(n_686),
.B1(n_689),
.B2(n_637),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_732),
.Y(n_760)
);

NOR2x1_ASAP7_75t_L g761 ( 
.A(n_739),
.B(n_643),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_713),
.B(n_689),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_736),
.B(n_643),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_733),
.B(n_639),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_702),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_715),
.Y(n_766)
);

INVxp67_ASAP7_75t_SL g767 ( 
.A(n_738),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_731),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_712),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_714),
.Y(n_770)
);

INVxp33_ASAP7_75t_L g771 ( 
.A(n_718),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_709),
.B(n_645),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_701),
.B(n_630),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_709),
.B(n_630),
.Y(n_774)
);

OAI221xp5_ASAP7_75t_SL g775 ( 
.A1(n_701),
.A2(n_645),
.B1(n_648),
.B2(n_137),
.C(n_140),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_727),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_703),
.B(n_620),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_717),
.Y(n_778)
);

OR2x2_ASAP7_75t_L g779 ( 
.A(n_709),
.B(n_648),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_721),
.B(n_131),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_756),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_769),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_746),
.B(n_740),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_756),
.B(n_698),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_769),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_748),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_748),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_754),
.B(n_755),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_764),
.B(n_741),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_757),
.B(n_741),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_774),
.B(n_725),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_744),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_743),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_744),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_765),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_753),
.B(n_718),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_776),
.Y(n_797)
);

OR2x2_ASAP7_75t_L g798 ( 
.A(n_750),
.B(n_704),
.Y(n_798)
);

AND2x4_ASAP7_75t_L g799 ( 
.A(n_772),
.B(n_725),
.Y(n_799)
);

NOR3xp33_ASAP7_75t_L g800 ( 
.A(n_775),
.B(n_724),
.C(n_727),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_747),
.B(n_695),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_762),
.A2(n_700),
.B1(n_735),
.B2(n_696),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_760),
.Y(n_803)
);

BUFx2_ASAP7_75t_L g804 ( 
.A(n_766),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_751),
.B(n_735),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_752),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_747),
.B(n_745),
.Y(n_807)
);

AND2x2_ASAP7_75t_SL g808 ( 
.A(n_773),
.B(n_699),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_770),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_789),
.B(n_766),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_790),
.B(n_742),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_797),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_808),
.B(n_784),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_792),
.B(n_773),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_798),
.B(n_768),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_789),
.B(n_804),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_801),
.B(n_742),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_781),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_792),
.B(n_761),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_786),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_794),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_794),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_799),
.B(n_742),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_807),
.B(n_763),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_797),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_808),
.A2(n_800),
.B1(n_749),
.B2(n_759),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_799),
.B(n_771),
.Y(n_827)
);

OAI32xp33_ASAP7_75t_L g828 ( 
.A1(n_814),
.A2(n_783),
.A3(n_796),
.B1(n_771),
.B2(n_788),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_816),
.B(n_799),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_814),
.B(n_818),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_821),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_812),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_822),
.Y(n_833)
);

AOI22xp5_ASAP7_75t_L g834 ( 
.A1(n_826),
.A2(n_759),
.B1(n_802),
.B2(n_791),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_820),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_827),
.B(n_791),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_826),
.A2(n_791),
.B1(n_802),
.B2(n_780),
.Y(n_837)
);

OAI32xp33_ASAP7_75t_L g838 ( 
.A1(n_813),
.A2(n_793),
.A3(n_777),
.B1(n_779),
.B2(n_806),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_810),
.B(n_805),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_835),
.Y(n_840)
);

AOI221xp5_ASAP7_75t_L g841 ( 
.A1(n_838),
.A2(n_819),
.B1(n_775),
.B2(n_803),
.C(n_824),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_830),
.B(n_819),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_831),
.Y(n_843)
);

INVx1_ASAP7_75t_SL g844 ( 
.A(n_832),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_844),
.B(n_829),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_L g846 ( 
.A1(n_841),
.A2(n_834),
.B(n_837),
.Y(n_846)
);

INVxp67_ASAP7_75t_L g847 ( 
.A(n_840),
.Y(n_847)
);

NOR2x1_ASAP7_75t_L g848 ( 
.A(n_843),
.B(n_815),
.Y(n_848)
);

INVxp67_ASAP7_75t_SL g849 ( 
.A(n_842),
.Y(n_849)
);

NAND3xp33_ASAP7_75t_L g850 ( 
.A(n_846),
.B(n_834),
.C(n_833),
.Y(n_850)
);

O2A1O1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_847),
.A2(n_828),
.B(n_825),
.C(n_836),
.Y(n_851)
);

INVx1_ASAP7_75t_SL g852 ( 
.A(n_845),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_848),
.B(n_839),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_850),
.A2(n_849),
.B(n_823),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_SL g855 ( 
.A1(n_852),
.A2(n_817),
.B(n_811),
.Y(n_855)
);

AND4x1_ASAP7_75t_L g856 ( 
.A(n_851),
.B(n_730),
.C(n_711),
.D(n_817),
.Y(n_856)
);

NAND4xp25_ASAP7_75t_L g857 ( 
.A(n_853),
.B(n_758),
.C(n_811),
.D(n_795),
.Y(n_857)
);

NOR2x1p5_ASAP7_75t_L g858 ( 
.A(n_857),
.B(n_809),
.Y(n_858)
);

NOR2x1_ASAP7_75t_L g859 ( 
.A(n_855),
.B(n_809),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_854),
.A2(n_795),
.B1(n_787),
.B2(n_778),
.Y(n_860)
);

NAND2xp33_ASAP7_75t_L g861 ( 
.A(n_856),
.B(n_787),
.Y(n_861)
);

NOR2x1_ASAP7_75t_L g862 ( 
.A(n_861),
.B(n_785),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_860),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_859),
.A2(n_785),
.B1(n_782),
.B2(n_767),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_858),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_860),
.B(n_134),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_860),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_865),
.A2(n_767),
.B1(n_782),
.B2(n_706),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_867),
.Y(n_869)
);

OAI211xp5_ASAP7_75t_L g870 ( 
.A1(n_863),
.A2(n_632),
.B(n_142),
.C(n_144),
.Y(n_870)
);

NOR2x1_ASAP7_75t_L g871 ( 
.A(n_866),
.B(n_141),
.Y(n_871)
);

XOR2x1_ASAP7_75t_L g872 ( 
.A(n_862),
.B(n_145),
.Y(n_872)
);

NOR2x1_ASAP7_75t_L g873 ( 
.A(n_864),
.B(n_146),
.Y(n_873)
);

INVx3_ASAP7_75t_SL g874 ( 
.A(n_869),
.Y(n_874)
);

NAND2x1p5_ASAP7_75t_L g875 ( 
.A(n_871),
.B(n_148),
.Y(n_875)
);

BUFx4f_ASAP7_75t_SL g876 ( 
.A(n_872),
.Y(n_876)
);

INVx1_ASAP7_75t_SL g877 ( 
.A(n_873),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_870),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_868),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_869),
.A2(n_706),
.B1(n_150),
.B2(n_151),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_869),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_881),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_874),
.A2(n_706),
.B1(n_152),
.B2(n_153),
.Y(n_883)
);

AO22x2_ASAP7_75t_L g884 ( 
.A1(n_877),
.A2(n_879),
.B1(n_876),
.B2(n_880),
.Y(n_884)
);

XOR2xp5_ASAP7_75t_L g885 ( 
.A(n_875),
.B(n_149),
.Y(n_885)
);

INVxp67_ASAP7_75t_L g886 ( 
.A(n_878),
.Y(n_886)
);

AO22x2_ASAP7_75t_L g887 ( 
.A1(n_878),
.A2(n_157),
.B1(n_159),
.B2(n_161),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_874),
.B(n_164),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_881),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_876),
.A2(n_166),
.B1(n_167),
.B2(n_169),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_886),
.B(n_170),
.Y(n_891)
);

OAI22xp33_ASAP7_75t_L g892 ( 
.A1(n_888),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_887),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_885),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_894)
);

BUFx2_ASAP7_75t_SL g895 ( 
.A(n_882),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_893),
.Y(n_896)
);

OAI22x1_ASAP7_75t_L g897 ( 
.A1(n_891),
.A2(n_889),
.B1(n_890),
.B2(n_894),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_895),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_898),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_899),
.A2(n_897),
.B(n_896),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_900),
.A2(n_884),
.B1(n_883),
.B2(n_892),
.Y(n_901)
);

OR2x6_ASAP7_75t_L g902 ( 
.A(n_901),
.B(n_180),
.Y(n_902)
);

AOI211xp5_ASAP7_75t_L g903 ( 
.A1(n_902),
.A2(n_181),
.B(n_182),
.C(n_184),
.Y(n_903)
);


endmodule