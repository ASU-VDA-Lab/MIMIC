module fake_ariane_2891_n_2477 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_240, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_236, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_226, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_229, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_227, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_232, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_54, n_25, n_2477);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_240;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_236;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_226;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_229;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_54;
input n_25;

output n_2477;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2334;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_2407;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2374;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_2288;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_259;
wire n_2442;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_2233;
wire n_2370;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_2433;
wire n_352;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_2427;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_2456;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_461;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_249;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_2426;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_2415;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_967;
wire n_274;
wire n_1083;
wire n_437;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_2439;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_2400;
wire n_632;
wire n_477;
wire n_650;
wire n_2388;
wire n_425;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_489;
wire n_2294;
wire n_2274;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_397;
wire n_2467;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_307;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_2328;
wire n_347;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_299;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_2262;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_552;
wire n_348;
wire n_2312;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2059;
wire n_2437;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_677;
wire n_604;
wire n_439;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_321;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_2379;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_2266;
wire n_2449;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_2366;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_2474;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_2460;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1769;
wire n_1632;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_516;
wire n_2364;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_374;
wire n_1352;
wire n_2405;
wire n_1824;
wire n_643;
wire n_1492;
wire n_2383;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2320;
wire n_979;
wire n_2329;
wire n_1642;
wire n_2417;
wire n_1815;
wire n_897;
wire n_949;
wire n_2454;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_354;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2331;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_2444;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_243;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_2402;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_2395;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2440;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_2268;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_2445;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2463;
wire n_309;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_2397;
wire n_369;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_248;
wire n_1152;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_2422;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_2097;
wire n_1982;
wire n_662;
wire n_641;
wire n_2430;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_2381;
wire n_1967;
wire n_2384;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2318;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_2336;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_19),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_135),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_203),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_109),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_103),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_142),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_227),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_87),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_26),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_240),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_117),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_160),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_234),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_58),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_44),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_220),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_122),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_53),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_217),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_93),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_239),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_189),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_128),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_51),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_210),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_178),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_233),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_48),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_149),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_192),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_68),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_14),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_19),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_212),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_50),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_139),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_18),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_90),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_213),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_78),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_190),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_96),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_172),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_73),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_60),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_214),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_24),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_80),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_21),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_82),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_61),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_224),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_154),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_173),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_219),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_144),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_32),
.Y(n_297)
);

BUFx8_ASAP7_75t_SL g298 ( 
.A(n_40),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_147),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_8),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_99),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_65),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_131),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_140),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_93),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_82),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_113),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_36),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_0),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_67),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_6),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_202),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_2),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_27),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_31),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_17),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_41),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_132),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_111),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_18),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_24),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_26),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_127),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_0),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_183),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_22),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_158),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_62),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_185),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_123),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_138),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_35),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_99),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_237),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_141),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_94),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_230),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_226),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_80),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_114),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_155),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_164),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_216),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_58),
.Y(n_344)
);

BUFx5_ASAP7_75t_L g345 ( 
.A(n_59),
.Y(n_345)
);

INVx4_ASAP7_75t_R g346 ( 
.A(n_235),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_165),
.Y(n_347)
);

BUFx10_ASAP7_75t_L g348 ( 
.A(n_56),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_72),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_171),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_215),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_167),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_85),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_181),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_199),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_67),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_102),
.Y(n_357)
);

BUFx10_ASAP7_75t_L g358 ( 
.A(n_100),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_221),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_41),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_81),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_198),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_204),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_8),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_56),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_152),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_177),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_228),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_4),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_13),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_169),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_85),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_231),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_225),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_229),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_176),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_106),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_17),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_3),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_63),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_47),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_2),
.Y(n_382)
);

CKINVDCx14_ASAP7_75t_R g383 ( 
.A(n_146),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_197),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_143),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_95),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_223),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_73),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_42),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_168),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_110),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_1),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_211),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_207),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_64),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_107),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_27),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_236),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_61),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_35),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_89),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_13),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_104),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_74),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_83),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_5),
.Y(n_406)
);

BUFx2_ASAP7_75t_SL g407 ( 
.A(n_25),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_79),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_49),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_66),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_118),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_16),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_39),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_39),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_9),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_180),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_208),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_95),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_52),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_36),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_194),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_175),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_193),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_200),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_104),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_195),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_76),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_179),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_62),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_65),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_187),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_46),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_16),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_89),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_64),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_20),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_112),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_33),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_43),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_60),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_48),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_4),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_49),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_50),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_46),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_184),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_63),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_43),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_157),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_40),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_126),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_136),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_145),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_102),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_188),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_87),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_101),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_88),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_28),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_201),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_57),
.Y(n_461)
);

CKINVDCx14_ASAP7_75t_R g462 ( 
.A(n_68),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_25),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_33),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_137),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_125),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_55),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_11),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_103),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_88),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_6),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_166),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_269),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_345),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_436),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_345),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_345),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_298),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_345),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_345),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_345),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_345),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_268),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_269),
.B(n_1),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_302),
.B(n_3),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_345),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_345),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_268),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_243),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_251),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_462),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_246),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_253),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_251),
.B(n_5),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_279),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_286),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_252),
.Y(n_497)
);

BUFx6f_ASAP7_75t_SL g498 ( 
.A(n_263),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_252),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_257),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_330),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_257),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_340),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_436),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_367),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_373),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_261),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_421),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_261),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_270),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_432),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_296),
.B(n_7),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_432),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_463),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_280),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_270),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_276),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_276),
.B(n_7),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_241),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_324),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_294),
.Y(n_521)
);

INVxp33_ASAP7_75t_SL g522 ( 
.A(n_463),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_311),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_248),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_294),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_303),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_249),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_254),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_311),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_303),
.Y(n_530)
);

INVxp67_ASAP7_75t_SL g531 ( 
.A(n_438),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_318),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_318),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_272),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_323),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_323),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_273),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_275),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_284),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_337),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_438),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_326),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_400),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_337),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_351),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_351),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_354),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_285),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_287),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_354),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_288),
.Y(n_551)
);

INVxp67_ASAP7_75t_SL g552 ( 
.A(n_441),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_404),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_355),
.Y(n_554)
);

CKINVDCx16_ASAP7_75t_R g555 ( 
.A(n_341),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_355),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_362),
.Y(n_557)
);

NOR2xp67_ASAP7_75t_L g558 ( 
.A(n_322),
.B(n_9),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_268),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_362),
.Y(n_560)
);

INVxp67_ASAP7_75t_SL g561 ( 
.A(n_441),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_289),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_363),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_290),
.Y(n_564)
);

BUFx2_ASAP7_75t_SL g565 ( 
.A(n_263),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_420),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_322),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_297),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_300),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_407),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_363),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_371),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_371),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_341),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_375),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_305),
.Y(n_576)
);

BUFx6f_ASAP7_75t_SL g577 ( 
.A(n_263),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_308),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_375),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_313),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_428),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_384),
.B(n_10),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_428),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_384),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_385),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_385),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_390),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_314),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_316),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_390),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_465),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_391),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_320),
.Y(n_593)
);

INVxp33_ASAP7_75t_L g594 ( 
.A(n_245),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_391),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_332),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_349),
.Y(n_597)
);

INVxp67_ASAP7_75t_SL g598 ( 
.A(n_268),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_393),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_393),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_268),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_465),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_353),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_483),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_474),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_483),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_489),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_485),
.B(n_264),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_483),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_488),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_492),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_515),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_495),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_496),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_488),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_475),
.B(n_245),
.Y(n_616)
);

OA21x2_ASAP7_75t_L g617 ( 
.A1(n_490),
.A2(n_411),
.B(n_398),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_505),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_488),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_511),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_513),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_493),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_501),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_503),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_559),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_474),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_476),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_559),
.Y(n_628)
);

NOR2x1_ASAP7_75t_L g629 ( 
.A(n_565),
.B(n_293),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_476),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_506),
.Y(n_631)
);

INVxp67_ASAP7_75t_L g632 ( 
.A(n_565),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_601),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_601),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_477),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_485),
.B(n_317),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_477),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_574),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_479),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_479),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_490),
.B(n_383),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_480),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_480),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_R g644 ( 
.A(n_519),
.B(n_242),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_481),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_481),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_482),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_508),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_520),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_482),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_486),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_486),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_487),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_487),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_598),
.Y(n_655)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_581),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_570),
.B(n_455),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_478),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_524),
.Y(n_659)
);

XNOR2xp5_ASAP7_75t_L g660 ( 
.A(n_542),
.B(n_258),
.Y(n_660)
);

AND2x4_ASAP7_75t_L g661 ( 
.A(n_497),
.B(n_499),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_497),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_499),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_543),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_500),
.B(n_502),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_527),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_500),
.B(n_502),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_528),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_507),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_553),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_507),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_509),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_512),
.B(n_317),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_534),
.Y(n_674)
);

OAI21x1_ASAP7_75t_L g675 ( 
.A1(n_509),
.A2(n_411),
.B(n_398),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_537),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_538),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_510),
.B(n_264),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_539),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_566),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_510),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_516),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_516),
.B(n_278),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_491),
.Y(n_684)
);

OAI21x1_ASAP7_75t_L g685 ( 
.A1(n_517),
.A2(n_417),
.B(n_416),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_517),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_521),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_521),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_525),
.Y(n_689)
);

AND2x6_ASAP7_75t_L g690 ( 
.A(n_525),
.B(n_460),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_526),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_526),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_530),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_530),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_531),
.B(n_416),
.Y(n_695)
);

OA21x2_ASAP7_75t_L g696 ( 
.A1(n_532),
.A2(n_446),
.B(n_417),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_532),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_533),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_533),
.Y(n_699)
);

CKINVDCx20_ASAP7_75t_R g700 ( 
.A(n_583),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_535),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_548),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_642),
.Y(n_703)
);

INVx4_ASAP7_75t_L g704 ( 
.A(n_661),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_665),
.B(n_667),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_658),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_662),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_642),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_662),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_641),
.B(n_473),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_629),
.B(n_541),
.Y(n_711)
);

BUFx4f_ASAP7_75t_L g712 ( 
.A(n_617),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_669),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_663),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_641),
.B(n_473),
.Y(n_715)
);

INVx5_ASAP7_75t_L g716 ( 
.A(n_690),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_616),
.B(n_555),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_608),
.A2(n_522),
.B1(n_484),
.B2(n_518),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_605),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_642),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_663),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_682),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_605),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_682),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_616),
.B(n_475),
.Y(n_725)
);

INVx4_ASAP7_75t_SL g726 ( 
.A(n_690),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_669),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_642),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_632),
.B(n_549),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_669),
.Y(n_730)
);

AND2x6_ASAP7_75t_L g731 ( 
.A(n_641),
.B(n_446),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_694),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_629),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_616),
.B(n_514),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_655),
.B(n_498),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_694),
.Y(n_736)
);

XOR2xp5_ASAP7_75t_SL g737 ( 
.A(n_678),
.B(n_535),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_644),
.B(n_551),
.Y(n_738)
);

NAND2xp33_ASAP7_75t_R g739 ( 
.A(n_620),
.B(n_562),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_661),
.B(n_536),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_665),
.B(n_552),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_661),
.B(n_665),
.Y(n_742)
);

INVx4_ASAP7_75t_L g743 ( 
.A(n_661),
.Y(n_743)
);

AND2x6_ASAP7_75t_L g744 ( 
.A(n_661),
.B(n_449),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_697),
.Y(n_745)
);

INVx5_ASAP7_75t_L g746 ( 
.A(n_690),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_669),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_607),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_669),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_611),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_647),
.Y(n_751)
);

BUFx2_ASAP7_75t_L g752 ( 
.A(n_620),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_667),
.Y(n_753)
);

AND2x2_ASAP7_75t_SL g754 ( 
.A(n_617),
.B(n_494),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_613),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_626),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_626),
.Y(n_757)
);

AND2x6_ASAP7_75t_L g758 ( 
.A(n_667),
.B(n_449),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_627),
.Y(n_759)
);

AO21x2_ASAP7_75t_L g760 ( 
.A1(n_673),
.A2(n_453),
.B(n_451),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_686),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_647),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_686),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_657),
.B(n_498),
.Y(n_764)
);

INVx5_ASAP7_75t_L g765 ( 
.A(n_690),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_614),
.Y(n_766)
);

INVxp67_ASAP7_75t_L g767 ( 
.A(n_620),
.Y(n_767)
);

AND2x6_ASAP7_75t_L g768 ( 
.A(n_608),
.B(n_451),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_647),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_644),
.B(n_564),
.Y(n_770)
);

BUFx2_ASAP7_75t_L g771 ( 
.A(n_621),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_686),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_657),
.A2(n_568),
.B1(n_578),
.B2(n_569),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_605),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_618),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_636),
.B(n_498),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_636),
.B(n_577),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_627),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_608),
.B(n_536),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_617),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_647),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_659),
.B(n_580),
.Y(n_782)
);

AO21x2_ASAP7_75t_L g783 ( 
.A1(n_673),
.A2(n_685),
.B(n_675),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_669),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_669),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_608),
.B(n_540),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_687),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_608),
.B(n_577),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_605),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_666),
.B(n_588),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_687),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_687),
.Y(n_792)
);

INVx4_ASAP7_75t_L g793 ( 
.A(n_697),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_635),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_668),
.B(n_577),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_692),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_674),
.B(n_589),
.Y(n_797)
);

OR2x2_ASAP7_75t_L g798 ( 
.A(n_621),
.B(n_514),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_635),
.Y(n_799)
);

INVx4_ASAP7_75t_L g800 ( 
.A(n_697),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_669),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_692),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_635),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_637),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_672),
.Y(n_805)
);

INVx4_ASAP7_75t_L g806 ( 
.A(n_697),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_676),
.B(n_593),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_695),
.A2(n_582),
.B1(n_504),
.B2(n_567),
.Y(n_808)
);

BUFx2_ASAP7_75t_L g809 ( 
.A(n_621),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_678),
.B(n_561),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_637),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_692),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_605),
.Y(n_813)
);

OR2x6_ASAP7_75t_L g814 ( 
.A(n_678),
.B(n_558),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_677),
.B(n_596),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_672),
.Y(n_816)
);

BUFx4f_ASAP7_75t_L g817 ( 
.A(n_617),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_693),
.Y(n_818)
);

BUFx10_ASAP7_75t_L g819 ( 
.A(n_679),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_617),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_683),
.B(n_594),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_637),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_651),
.Y(n_823)
);

INVx4_ASAP7_75t_SL g824 ( 
.A(n_690),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_693),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_612),
.Y(n_826)
);

INVx1_ASAP7_75t_SL g827 ( 
.A(n_656),
.Y(n_827)
);

AND2x6_ASAP7_75t_L g828 ( 
.A(n_671),
.B(n_453),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_656),
.B(n_576),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_651),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_651),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_693),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_702),
.B(n_597),
.Y(n_833)
);

OR2x6_ASAP7_75t_L g834 ( 
.A(n_683),
.B(n_407),
.Y(n_834)
);

INVx4_ASAP7_75t_SL g835 ( 
.A(n_690),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_697),
.B(n_540),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_630),
.B(n_544),
.Y(n_837)
);

AND2x6_ASAP7_75t_L g838 ( 
.A(n_671),
.B(n_472),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_630),
.B(n_544),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_701),
.Y(n_840)
);

AND2x6_ASAP7_75t_L g841 ( 
.A(n_671),
.B(n_472),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_695),
.B(n_603),
.Y(n_842)
);

BUFx10_ASAP7_75t_L g843 ( 
.A(n_622),
.Y(n_843)
);

AO21x2_ASAP7_75t_L g844 ( 
.A1(n_675),
.A2(n_546),
.B(n_545),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_640),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_639),
.B(n_545),
.Y(n_846)
);

BUFx8_ASAP7_75t_SL g847 ( 
.A(n_612),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_683),
.B(n_567),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_672),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_701),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_701),
.B(n_546),
.Y(n_851)
);

INVx4_ASAP7_75t_L g852 ( 
.A(n_672),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_639),
.B(n_547),
.Y(n_853)
);

OR2x6_ASAP7_75t_L g854 ( 
.A(n_638),
.B(n_529),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_671),
.B(n_547),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_689),
.Y(n_856)
);

AND2x6_ASAP7_75t_L g857 ( 
.A(n_689),
.B(n_274),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_617),
.A2(n_554),
.B1(n_556),
.B2(n_550),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_696),
.Y(n_859)
);

NAND2x1p5_ASAP7_75t_L g860 ( 
.A(n_696),
.B(n_550),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_689),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_645),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_672),
.Y(n_863)
);

CKINVDCx20_ASAP7_75t_R g864 ( 
.A(n_649),
.Y(n_864)
);

OR2x2_ASAP7_75t_L g865 ( 
.A(n_638),
.B(n_523),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_842),
.B(n_591),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_704),
.B(n_602),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_758),
.A2(n_696),
.B1(n_691),
.B2(n_689),
.Y(n_868)
);

NAND2x1p5_ASAP7_75t_L g869 ( 
.A(n_704),
.B(n_696),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_764),
.B(n_640),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_731),
.B(n_735),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_731),
.B(n_640),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_731),
.B(n_640),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_856),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_731),
.B(n_654),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_731),
.B(n_654),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_794),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_731),
.B(n_654),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_745),
.A2(n_646),
.B(n_645),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_704),
.A2(n_698),
.B1(n_699),
.B2(n_691),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_743),
.A2(n_698),
.B1(n_699),
.B2(n_691),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_705),
.B(n_654),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_745),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_745),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_754),
.A2(n_696),
.B1(n_556),
.B2(n_557),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_712),
.A2(n_685),
.B(n_675),
.Y(n_886)
);

AO22x1_ASAP7_75t_L g887 ( 
.A1(n_758),
.A2(n_698),
.B1(n_699),
.B2(n_691),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_861),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_743),
.B(n_672),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_793),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_797),
.B(n_638),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_743),
.B(n_698),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_705),
.B(n_654),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_821),
.B(n_699),
.Y(n_894)
);

INVxp67_ASAP7_75t_L g895 ( 
.A(n_752),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_807),
.B(n_623),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_761),
.Y(n_897)
);

NAND2x1p5_ASAP7_75t_L g898 ( 
.A(n_712),
.B(n_696),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_711),
.B(n_646),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_758),
.A2(n_754),
.B1(n_744),
.B2(n_768),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_815),
.B(n_624),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_763),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_711),
.B(n_652),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_711),
.B(n_652),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_767),
.B(n_631),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_758),
.A2(n_653),
.B1(n_681),
.B2(n_672),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_793),
.A2(n_653),
.B(n_643),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_712),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_817),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_834),
.B(n_554),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_773),
.B(n_672),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_795),
.B(n_681),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_733),
.B(n_681),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_758),
.A2(n_688),
.B1(n_681),
.B2(n_327),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_772),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_718),
.A2(n_361),
.B1(n_369),
.B2(n_357),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_729),
.B(n_648),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_752),
.B(n_681),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_L g919 ( 
.A1(n_758),
.A2(n_560),
.B1(n_563),
.B2(n_557),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_821),
.B(n_560),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_733),
.B(n_681),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_771),
.B(n_681),
.Y(n_922)
);

BUFx8_ASAP7_75t_L g923 ( 
.A(n_771),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_817),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_717),
.B(n_700),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_741),
.B(n_563),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_817),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_794),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_788),
.B(n_681),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_741),
.B(n_688),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_742),
.A2(n_685),
.B(n_572),
.C(n_573),
.Y(n_931)
);

INVx3_ASAP7_75t_L g932 ( 
.A(n_793),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_799),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_829),
.Y(n_934)
);

NOR3xp33_ASAP7_75t_L g935 ( 
.A(n_809),
.B(n_301),
.C(n_271),
.Y(n_935)
);

OR2x6_ASAP7_75t_L g936 ( 
.A(n_834),
.B(n_278),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_787),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_799),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_768),
.A2(n_744),
.B1(n_810),
.B2(n_834),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_810),
.B(n_688),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_800),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_810),
.B(n_688),
.Y(n_942)
);

OR2x6_ASAP7_75t_L g943 ( 
.A(n_834),
.B(n_310),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_803),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_740),
.B(n_851),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_791),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_809),
.B(n_688),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_800),
.Y(n_948)
);

INVxp67_ASAP7_75t_L g949 ( 
.A(n_829),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_800),
.Y(n_950)
);

AOI22xp33_ASAP7_75t_L g951 ( 
.A1(n_768),
.A2(n_572),
.B1(n_573),
.B2(n_571),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_776),
.B(n_688),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_803),
.Y(n_953)
);

CKINVDCx16_ASAP7_75t_R g954 ( 
.A(n_739),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_848),
.B(n_571),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_806),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_777),
.B(n_688),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_753),
.B(n_575),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_819),
.Y(n_959)
);

AO22x1_ASAP7_75t_L g960 ( 
.A1(n_744),
.A2(n_579),
.B1(n_584),
.B2(n_575),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_779),
.B(n_579),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_806),
.A2(n_643),
.B(n_605),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_804),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_804),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_819),
.B(n_348),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_819),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_806),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_768),
.A2(n_327),
.B1(n_244),
.B2(n_584),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_811),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_786),
.B(n_585),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_855),
.B(n_768),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_738),
.B(n_348),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_780),
.A2(n_609),
.B(n_606),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_855),
.B(n_585),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_792),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_855),
.B(n_586),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_768),
.B(n_586),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_770),
.B(n_348),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_707),
.B(n_587),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_717),
.B(n_700),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_848),
.B(n_587),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_709),
.B(n_590),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_714),
.B(n_721),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_811),
.Y(n_984)
);

INVxp67_ASAP7_75t_L g985 ( 
.A(n_827),
.Y(n_985)
);

HB1xp67_ASAP7_75t_L g986 ( 
.A(n_865),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_798),
.B(n_649),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_722),
.B(n_590),
.Y(n_988)
);

NOR2xp67_ASAP7_75t_SL g989 ( 
.A(n_780),
.B(n_820),
.Y(n_989)
);

AND2x6_ASAP7_75t_SL g990 ( 
.A(n_847),
.B(n_255),
.Y(n_990)
);

NAND2x1_ASAP7_75t_L g991 ( 
.A(n_852),
.B(n_690),
.Y(n_991)
);

NAND2x1_ASAP7_75t_L g992 ( 
.A(n_852),
.B(n_690),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_724),
.B(n_592),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_860),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_719),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_750),
.B(n_348),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_750),
.B(n_358),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_732),
.B(n_592),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_755),
.B(n_358),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_755),
.B(n_766),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_736),
.B(n_595),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_756),
.B(n_595),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_854),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_756),
.B(n_599),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_757),
.B(n_599),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_744),
.A2(n_600),
.B1(n_263),
.B2(n_281),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_757),
.B(n_600),
.Y(n_1007)
);

OAI22x1_ASAP7_75t_SL g1008 ( 
.A1(n_826),
.A2(n_670),
.B1(n_680),
.B2(n_664),
.Y(n_1008)
);

AOI22xp33_ASAP7_75t_L g1009 ( 
.A1(n_744),
.A2(n_281),
.B1(n_447),
.B2(n_358),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_766),
.B(n_358),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_759),
.A2(n_378),
.B1(n_379),
.B2(n_370),
.Y(n_1011)
);

A2O1A1Ixp33_ASAP7_75t_SL g1012 ( 
.A1(n_713),
.A2(n_604),
.B(n_609),
.C(n_606),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_775),
.B(n_380),
.Y(n_1013)
);

AOI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_744),
.A2(n_838),
.B1(n_841),
.B2(n_828),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_822),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_796),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_759),
.B(n_604),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_706),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_778),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_719),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_798),
.B(n_664),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_775),
.B(n_381),
.Y(n_1022)
);

AOI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_814),
.A2(n_244),
.B1(n_374),
.B2(n_283),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_706),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_843),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_814),
.A2(n_250),
.B1(n_256),
.B2(n_247),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_782),
.B(n_670),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_778),
.B(n_604),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_862),
.Y(n_1029)
);

AND2x6_ASAP7_75t_SL g1030 ( 
.A(n_847),
.B(n_255),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_790),
.B(n_386),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_862),
.B(n_604),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_808),
.A2(n_395),
.B1(n_402),
.B2(n_389),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_822),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_710),
.B(n_604),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_715),
.B(n_610),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_833),
.B(n_680),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_802),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_940),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_949),
.B(n_865),
.Y(n_1040)
);

INVxp67_ASAP7_75t_L g1041 ( 
.A(n_934),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_942),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_R g1043 ( 
.A(n_1018),
.B(n_826),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_892),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_926),
.B(n_814),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_926),
.B(n_920),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_959),
.Y(n_1047)
);

NOR3xp33_ASAP7_75t_SL g1048 ( 
.A(n_1018),
.B(n_405),
.C(n_403),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_920),
.B(n_814),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_908),
.Y(n_1050)
);

AOI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_866),
.A2(n_748),
.B1(n_854),
.B2(n_820),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_894),
.B(n_837),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_908),
.Y(n_1053)
);

INVxp67_ASAP7_75t_L g1054 ( 
.A(n_987),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_877),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_900),
.A2(n_828),
.B1(n_841),
.B2(n_838),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_908),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_892),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_892),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_894),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_923),
.Y(n_1061)
);

BUFx3_ASAP7_75t_L g1062 ( 
.A(n_1024),
.Y(n_1062)
);

INVx4_ASAP7_75t_L g1063 ( 
.A(n_959),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_900),
.B(n_719),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_897),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_955),
.B(n_981),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_955),
.B(n_839),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_908),
.B(n_719),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_891),
.B(n_854),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_981),
.B(n_846),
.Y(n_1070)
);

INVx4_ASAP7_75t_L g1071 ( 
.A(n_966),
.Y(n_1071)
);

INVx5_ASAP7_75t_L g1072 ( 
.A(n_908),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_910),
.B(n_853),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_910),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_910),
.B(n_836),
.Y(n_1075)
);

INVx5_ASAP7_75t_L g1076 ( 
.A(n_927),
.Y(n_1076)
);

BUFx3_ASAP7_75t_L g1077 ( 
.A(n_1024),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_986),
.B(n_725),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_1019),
.Y(n_1079)
);

AOI222xp33_ASAP7_75t_L g1080 ( 
.A1(n_1008),
.A2(n_660),
.B1(n_864),
.B2(n_684),
.C1(n_364),
.C2(n_333),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_895),
.B(n_854),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_927),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_1025),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_927),
.B(n_719),
.Y(n_1084)
);

NOR2x1_ASAP7_75t_L g1085 ( 
.A(n_1025),
.B(n_725),
.Y(n_1085)
);

OR2x2_ASAP7_75t_L g1086 ( 
.A(n_1021),
.B(n_734),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_945),
.B(n_858),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_1019),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_927),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_897),
.Y(n_1090)
);

NOR3xp33_ASAP7_75t_SL g1091 ( 
.A(n_1000),
.B(n_410),
.C(n_408),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_954),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_927),
.B(n_723),
.Y(n_1093)
);

INVxp67_ASAP7_75t_L g1094 ( 
.A(n_985),
.Y(n_1094)
);

NOR3xp33_ASAP7_75t_L g1095 ( 
.A(n_896),
.B(n_734),
.C(n_277),
.Y(n_1095)
);

AOI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_939),
.A2(n_859),
.B1(n_843),
.B2(n_860),
.Y(n_1096)
);

AND2x6_ASAP7_75t_L g1097 ( 
.A(n_1014),
.B(n_737),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_902),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_899),
.B(n_860),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_903),
.B(n_859),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_954),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_904),
.B(n_845),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_918),
.B(n_845),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_877),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_909),
.B(n_723),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_1019),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_885),
.A2(n_828),
.B1(n_841),
.B2(n_838),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_901),
.B(n_843),
.Y(n_1108)
);

INVx5_ASAP7_75t_L g1109 ( 
.A(n_995),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_966),
.B(n_726),
.Y(n_1110)
);

OR2x6_ASAP7_75t_L g1111 ( 
.A(n_936),
.B(n_737),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_SL g1112 ( 
.A1(n_925),
.A2(n_864),
.B1(n_684),
.B2(n_660),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_928),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_905),
.B(n_660),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_1029),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_923),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_928),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_902),
.Y(n_1118)
);

INVx5_ASAP7_75t_L g1119 ( 
.A(n_995),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_915),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_882),
.B(n_812),
.Y(n_1121)
);

XNOR2xp5_ASAP7_75t_L g1122 ( 
.A(n_1008),
.B(n_1003),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_933),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_893),
.B(n_818),
.Y(n_1124)
);

NOR3xp33_ASAP7_75t_SL g1125 ( 
.A(n_1013),
.B(n_414),
.C(n_412),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_995),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_915),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_933),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1002),
.B(n_825),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_1029),
.Y(n_1130)
);

BUFx10_ASAP7_75t_L g1131 ( 
.A(n_980),
.Y(n_1131)
);

NOR3xp33_ASAP7_75t_SL g1132 ( 
.A(n_1022),
.B(n_425),
.C(n_418),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_995),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_916),
.A2(n_840),
.B(n_850),
.C(n_832),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_1003),
.B(n_703),
.Y(n_1135)
);

NOR3xp33_ASAP7_75t_SL g1136 ( 
.A(n_922),
.B(n_433),
.C(n_427),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_936),
.B(n_726),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_923),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_937),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_936),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_938),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_937),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_946),
.Y(n_1143)
);

INVx5_ASAP7_75t_L g1144 ( 
.A(n_995),
.Y(n_1144)
);

OR2x2_ASAP7_75t_L g1145 ( 
.A(n_1027),
.B(n_760),
.Y(n_1145)
);

INVxp33_ASAP7_75t_SL g1146 ( 
.A(n_1037),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_936),
.B(n_726),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_971),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_946),
.Y(n_1149)
);

AND2x6_ASAP7_75t_L g1150 ( 
.A(n_1014),
.B(n_703),
.Y(n_1150)
);

CKINVDCx6p67_ASAP7_75t_R g1151 ( 
.A(n_943),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_943),
.B(n_947),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_938),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_909),
.B(n_723),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_1020),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1009),
.A2(n_917),
.B1(n_943),
.B2(n_871),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1004),
.B(n_823),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1005),
.B(n_823),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_1020),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_867),
.B(n_852),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_975),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_R g1162 ( 
.A(n_924),
.B(n_713),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_1020),
.Y(n_1163)
);

NOR3xp33_ASAP7_75t_SL g1164 ( 
.A(n_889),
.B(n_435),
.C(n_434),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_975),
.Y(n_1165)
);

AND2x6_ASAP7_75t_L g1166 ( 
.A(n_868),
.B(n_708),
.Y(n_1166)
);

CKINVDCx20_ASAP7_75t_R g1167 ( 
.A(n_1031),
.Y(n_1167)
);

BUFx8_ASAP7_75t_SL g1168 ( 
.A(n_943),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_960),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1007),
.B(n_830),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_944),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_935),
.B(n_708),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_930),
.B(n_830),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1016),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1016),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_974),
.B(n_831),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_976),
.B(n_720),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_1029),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_960),
.Y(n_1179)
);

NAND3xp33_ASAP7_75t_L g1180 ( 
.A(n_1033),
.B(n_784),
.C(n_747),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_944),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_924),
.B(n_723),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_958),
.B(n_720),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1038),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_977),
.Y(n_1185)
);

INVx2_ASAP7_75t_SL g1186 ( 
.A(n_965),
.Y(n_1186)
);

INVx4_ASAP7_75t_L g1187 ( 
.A(n_1020),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_953),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_883),
.B(n_723),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_961),
.B(n_728),
.Y(n_1190)
);

INVx5_ASAP7_75t_L g1191 ( 
.A(n_1020),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_869),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1038),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_870),
.A2(n_727),
.B1(n_730),
.B2(n_713),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1023),
.B(n_727),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_874),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_874),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_953),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_963),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_994),
.B(n_726),
.Y(n_1200)
);

AOI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1006),
.A2(n_730),
.B1(n_749),
.B2(n_727),
.Y(n_1201)
);

NOR3xp33_ASAP7_75t_SL g1202 ( 
.A(n_996),
.B(n_442),
.C(n_440),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_970),
.B(n_728),
.Y(n_1203)
);

AND2x6_ASAP7_75t_L g1204 ( 
.A(n_868),
.B(n_751),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_888),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_888),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1011),
.B(n_751),
.Y(n_1207)
);

OR2x2_ASAP7_75t_SL g1208 ( 
.A(n_990),
.B(n_310),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_983),
.B(n_1036),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1035),
.B(n_730),
.Y(n_1210)
);

CKINVDCx20_ASAP7_75t_R g1211 ( 
.A(n_997),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_963),
.Y(n_1212)
);

AND3x1_ASAP7_75t_SL g1213 ( 
.A(n_1030),
.B(n_277),
.C(n_260),
.Y(n_1213)
);

AOI21x1_ASAP7_75t_L g1214 ( 
.A1(n_989),
.A2(n_784),
.B(n_747),
.Y(n_1214)
);

NOR3xp33_ASAP7_75t_SL g1215 ( 
.A(n_999),
.B(n_444),
.C(n_443),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_994),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1026),
.B(n_762),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_964),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_911),
.A2(n_785),
.B1(n_816),
.B2(n_749),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_964),
.Y(n_1220)
);

OR2x2_ASAP7_75t_SL g1221 ( 
.A(n_979),
.B(n_336),
.Y(n_1221)
);

AND2x4_ASAP7_75t_SL g1222 ( 
.A(n_919),
.B(n_951),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_883),
.B(n_774),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_898),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_982),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_988),
.B(n_762),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_1010),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_993),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_969),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_998),
.B(n_1001),
.Y(n_1230)
);

NAND3xp33_ASAP7_75t_SL g1231 ( 
.A(n_968),
.B(n_450),
.C(n_445),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1214),
.A2(n_886),
.B(n_898),
.Y(n_1232)
);

NAND2xp33_ASAP7_75t_L g1233 ( 
.A(n_1126),
.B(n_883),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1074),
.B(n_884),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1062),
.Y(n_1235)
);

A2O1A1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1069),
.A2(n_931),
.B(n_879),
.C(n_973),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1069),
.B(n_887),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1103),
.A2(n_873),
.B(n_872),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1209),
.A2(n_929),
.B(n_890),
.Y(n_1239)
);

AOI221x1_ASAP7_75t_L g1240 ( 
.A1(n_1095),
.A2(n_952),
.B1(n_957),
.B2(n_881),
.C(n_880),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1146),
.B(n_972),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1103),
.A2(n_876),
.B(n_875),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1210),
.A2(n_878),
.B(n_869),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_1043),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1068),
.A2(n_898),
.B(n_962),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1046),
.B(n_887),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1068),
.A2(n_907),
.B(n_869),
.Y(n_1247)
);

NAND2x1_ASAP7_75t_L g1248 ( 
.A(n_1187),
.B(n_884),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1210),
.A2(n_906),
.B(n_1017),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1180),
.A2(n_1032),
.B(n_1028),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1066),
.B(n_969),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1067),
.B(n_984),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1070),
.B(n_984),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1084),
.A2(n_921),
.B(n_913),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1230),
.A2(n_890),
.B1(n_932),
.B2(n_884),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_1126),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1084),
.A2(n_1034),
.B(n_1015),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1055),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1126),
.Y(n_1259)
);

CKINVDCx16_ASAP7_75t_R g1260 ( 
.A(n_1043),
.Y(n_1260)
);

NOR2xp67_ASAP7_75t_L g1261 ( 
.A(n_1094),
.B(n_978),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1074),
.B(n_890),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1065),
.Y(n_1263)
);

INVx4_ASAP7_75t_L g1264 ( 
.A(n_1109),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1093),
.A2(n_1034),
.B(n_1015),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1099),
.A2(n_914),
.B(n_932),
.Y(n_1266)
);

AO21x2_ASAP7_75t_L g1267 ( 
.A1(n_1093),
.A2(n_912),
.B(n_1012),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1064),
.A2(n_781),
.B(n_769),
.Y(n_1268)
);

INVx3_ASAP7_75t_L g1269 ( 
.A(n_1126),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1137),
.B(n_932),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1064),
.A2(n_781),
.B(n_801),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1225),
.B(n_941),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1055),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1086),
.B(n_760),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1113),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1114),
.B(n_456),
.Y(n_1276)
);

BUFx8_ASAP7_75t_SL g1277 ( 
.A(n_1061),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1194),
.A2(n_805),
.B(n_801),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1090),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1078),
.B(n_457),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1095),
.B(n_458),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1062),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1105),
.A2(n_863),
.B(n_805),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1228),
.B(n_941),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1060),
.B(n_948),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1098),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1072),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1105),
.A2(n_863),
.B(n_991),
.Y(n_1288)
);

NAND2x1p5_ASAP7_75t_L g1289 ( 
.A(n_1072),
.B(n_1076),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1154),
.A2(n_992),
.B(n_991),
.Y(n_1290)
);

BUFx12f_ASAP7_75t_L g1291 ( 
.A(n_1116),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1137),
.B(n_948),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1108),
.B(n_950),
.Y(n_1293)
);

AOI21xp33_ASAP7_75t_L g1294 ( 
.A1(n_1054),
.A2(n_760),
.B(n_992),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1102),
.A2(n_956),
.B(n_950),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1072),
.B(n_950),
.Y(n_1296)
);

OR2x2_ASAP7_75t_L g1297 ( 
.A(n_1040),
.B(n_1041),
.Y(n_1297)
);

AO31x2_ASAP7_75t_L g1298 ( 
.A1(n_1113),
.A2(n_628),
.A3(n_633),
.B(n_625),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1052),
.A2(n_967),
.B(n_956),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1045),
.B(n_967),
.Y(n_1300)
);

AO31x2_ASAP7_75t_L g1301 ( 
.A1(n_1117),
.A2(n_628),
.A3(n_633),
.B(n_625),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1051),
.B(n_749),
.Y(n_1302)
);

INVxp67_ASAP7_75t_L g1303 ( 
.A(n_1081),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1072),
.B(n_774),
.Y(n_1304)
);

NAND3x1_ASAP7_75t_L g1305 ( 
.A(n_1156),
.B(n_282),
.C(n_260),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1154),
.A2(n_816),
.B(n_785),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1049),
.B(n_785),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1073),
.B(n_816),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1183),
.A2(n_989),
.B(n_789),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1118),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1182),
.A2(n_849),
.B(n_628),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1077),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1182),
.A2(n_849),
.B(n_633),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1117),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1121),
.A2(n_789),
.B(n_774),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_1076),
.B(n_774),
.Y(n_1316)
);

AO32x2_ASAP7_75t_L g1317 ( 
.A1(n_1140),
.A2(n_844),
.A3(n_841),
.B1(n_838),
.B2(n_828),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1123),
.Y(n_1318)
);

INVx4_ASAP7_75t_L g1319 ( 
.A(n_1109),
.Y(n_1319)
);

INVx4_ASAP7_75t_L g1320 ( 
.A(n_1109),
.Y(n_1320)
);

NAND2x1p5_ASAP7_75t_L g1321 ( 
.A(n_1076),
.B(n_849),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1076),
.B(n_774),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1134),
.A2(n_634),
.B(n_625),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1173),
.A2(n_634),
.B(n_295),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_SL g1325 ( 
.A(n_1050),
.B(n_789),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1039),
.B(n_789),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_SL g1327 ( 
.A1(n_1187),
.A2(n_377),
.B(n_336),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1124),
.A2(n_1203),
.B(n_1190),
.Y(n_1328)
);

AOI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1189),
.A2(n_634),
.B(n_615),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1042),
.B(n_789),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1081),
.B(n_813),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1189),
.A2(n_295),
.B(n_274),
.Y(n_1332)
);

AOI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1223),
.A2(n_615),
.B(n_610),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1148),
.B(n_813),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1148),
.B(n_813),
.Y(n_1335)
);

AOI211x1_ASAP7_75t_L g1336 ( 
.A1(n_1120),
.A2(n_306),
.B(n_309),
.C(n_315),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1223),
.A2(n_813),
.B(n_844),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1131),
.B(n_813),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1226),
.A2(n_844),
.B(n_783),
.Y(n_1339)
);

INVx3_ASAP7_75t_L g1340 ( 
.A(n_1133),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1157),
.A2(n_1170),
.B(n_1158),
.Y(n_1341)
);

OAI21xp33_ASAP7_75t_L g1342 ( 
.A1(n_1075),
.A2(n_461),
.B(n_459),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1044),
.B(n_828),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1219),
.A2(n_838),
.B(n_828),
.Y(n_1344)
);

AND2x6_ASAP7_75t_SL g1345 ( 
.A(n_1195),
.B(n_282),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1058),
.B(n_838),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1131),
.B(n_467),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1138),
.B(n_1092),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1129),
.A2(n_350),
.B(n_619),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1100),
.A2(n_783),
.B(n_643),
.Y(n_1350)
);

AOI21xp33_ASAP7_75t_L g1351 ( 
.A1(n_1145),
.A2(n_783),
.B(n_469),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1123),
.A2(n_350),
.B(n_619),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1128),
.A2(n_306),
.B(n_291),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1177),
.A2(n_643),
.B(n_605),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1059),
.B(n_841),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1087),
.A2(n_643),
.B(n_605),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1147),
.B(n_824),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1172),
.B(n_841),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1127),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1139),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1142),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1201),
.A2(n_857),
.B(n_690),
.Y(n_1362)
);

AOI21x1_ASAP7_75t_SL g1363 ( 
.A1(n_1207),
.A2(n_857),
.B(n_10),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1143),
.B(n_468),
.Y(n_1364)
);

BUFx3_ASAP7_75t_L g1365 ( 
.A(n_1077),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1176),
.A2(n_650),
.B(n_643),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1138),
.B(n_291),
.Y(n_1367)
);

OAI21xp33_ASAP7_75t_L g1368 ( 
.A1(n_1149),
.A2(n_315),
.B(n_309),
.Y(n_1368)
);

OA21x2_ASAP7_75t_L g1369 ( 
.A1(n_1128),
.A2(n_1181),
.B(n_1153),
.Y(n_1369)
);

NOR2x1_ASAP7_75t_L g1370 ( 
.A(n_1083),
.B(n_293),
.Y(n_1370)
);

AOI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1161),
.A2(n_333),
.B(n_321),
.Y(n_1371)
);

AO21x2_ASAP7_75t_L g1372 ( 
.A1(n_1196),
.A2(n_339),
.B(n_321),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1165),
.B(n_339),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1153),
.A2(n_1188),
.B(n_1181),
.Y(n_1374)
);

A2O1A1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1195),
.A2(n_382),
.B(n_399),
.C(n_401),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1174),
.B(n_356),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1147),
.B(n_824),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1188),
.A2(n_360),
.B(n_356),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1197),
.A2(n_650),
.B(n_643),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1175),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1184),
.B(n_360),
.Y(n_1381)
);

AO31x2_ASAP7_75t_L g1382 ( 
.A1(n_1198),
.A2(n_415),
.A3(n_364),
.B(n_365),
.Y(n_1382)
);

AO31x2_ASAP7_75t_L g1383 ( 
.A1(n_1198),
.A2(n_419),
.A3(n_365),
.B(n_372),
.Y(n_1383)
);

BUFx2_ASAP7_75t_SL g1384 ( 
.A(n_1083),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1193),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1199),
.A2(n_382),
.B(n_372),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1110),
.B(n_824),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1205),
.Y(n_1388)
);

AOI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1206),
.A2(n_392),
.B(n_388),
.Y(n_1389)
);

A2O1A1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1160),
.A2(n_392),
.B(n_415),
.C(n_419),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_SL g1391 ( 
.A1(n_1056),
.A2(n_397),
.B(n_377),
.Y(n_1391)
);

OAI21xp33_ASAP7_75t_L g1392 ( 
.A1(n_1125),
.A2(n_399),
.B(n_388),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1133),
.A2(n_650),
.B(n_643),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1133),
.A2(n_650),
.B(n_262),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1110),
.B(n_824),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1104),
.Y(n_1396)
);

AOI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1112),
.A2(n_857),
.B1(n_397),
.B2(n_413),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1133),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1141),
.Y(n_1399)
);

AO31x2_ASAP7_75t_L g1400 ( 
.A1(n_1240),
.A2(n_1199),
.A3(n_1218),
.B(n_1212),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1369),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1270),
.B(n_1111),
.Y(n_1402)
);

AO21x1_ASAP7_75t_L g1403 ( 
.A1(n_1351),
.A2(n_1302),
.B(n_1328),
.Y(n_1403)
);

NAND2x1p5_ASAP7_75t_L g1404 ( 
.A(n_1264),
.B(n_1192),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1233),
.A2(n_1119),
.B(n_1109),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1263),
.Y(n_1406)
);

AO21x2_ASAP7_75t_L g1407 ( 
.A1(n_1356),
.A2(n_1096),
.B(n_1162),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1279),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1369),
.Y(n_1409)
);

BUFx10_ASAP7_75t_L g1410 ( 
.A(n_1338),
.Y(n_1410)
);

OAI211xp5_ASAP7_75t_L g1411 ( 
.A1(n_1281),
.A2(n_1080),
.B(n_1091),
.C(n_1125),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1286),
.B(n_1111),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1234),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1324),
.A2(n_1218),
.B(n_1212),
.Y(n_1414)
);

INVx3_ASAP7_75t_L g1415 ( 
.A(n_1264),
.Y(n_1415)
);

OAI21xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1293),
.A2(n_1056),
.B(n_1107),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1324),
.A2(n_1229),
.B(n_1220),
.Y(n_1417)
);

OA21x2_ASAP7_75t_L g1418 ( 
.A1(n_1349),
.A2(n_1229),
.B(n_1220),
.Y(n_1418)
);

AO21x2_ASAP7_75t_L g1419 ( 
.A1(n_1339),
.A2(n_1162),
.B(n_1179),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1349),
.A2(n_1171),
.B(n_1088),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1310),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1332),
.A2(n_1088),
.B(n_1079),
.Y(n_1422)
);

AO21x2_ASAP7_75t_L g1423 ( 
.A1(n_1350),
.A2(n_1179),
.B(n_1160),
.Y(n_1423)
);

OAI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1266),
.A2(n_1217),
.B(n_1231),
.Y(n_1424)
);

BUFx12f_ASAP7_75t_L g1425 ( 
.A(n_1291),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1270),
.B(n_1111),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1369),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1332),
.A2(n_1106),
.B(n_1079),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1297),
.B(n_1101),
.Y(n_1429)
);

O2A1O1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1375),
.A2(n_1186),
.B(n_1132),
.C(n_1091),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1270),
.B(n_1292),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1280),
.B(n_1085),
.Y(n_1432)
);

AO31x2_ASAP7_75t_L g1433 ( 
.A1(n_1236),
.A2(n_1169),
.A3(n_1204),
.B(n_1166),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1352),
.A2(n_1115),
.B(n_1106),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1374),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1352),
.A2(n_1130),
.B(n_1115),
.Y(n_1436)
);

A2O1A1Ixp33_ASAP7_75t_L g1437 ( 
.A1(n_1375),
.A2(n_1222),
.B(n_1132),
.C(n_1107),
.Y(n_1437)
);

NAND2x1_ASAP7_75t_L g1438 ( 
.A(n_1264),
.B(n_1155),
.Y(n_1438)
);

OA21x2_ASAP7_75t_L g1439 ( 
.A1(n_1278),
.A2(n_1341),
.B(n_1232),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1278),
.A2(n_1178),
.B(n_1130),
.Y(n_1440)
);

OAI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1260),
.A2(n_1227),
.B1(n_1211),
.B2(n_1167),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1233),
.A2(n_1144),
.B(n_1119),
.Y(n_1442)
);

INVxp67_ASAP7_75t_SL g1443 ( 
.A(n_1234),
.Y(n_1443)
);

OA21x2_ASAP7_75t_L g1444 ( 
.A1(n_1341),
.A2(n_1164),
.B(n_1136),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1235),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1234),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1303),
.B(n_1135),
.Y(n_1447)
);

OAI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1249),
.A2(n_1204),
.B(n_1166),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1359),
.Y(n_1449)
);

AO21x2_ASAP7_75t_L g1450 ( 
.A1(n_1337),
.A2(n_1164),
.B(n_1136),
.Y(n_1450)
);

NAND3xp33_ASAP7_75t_L g1451 ( 
.A(n_1390),
.B(n_1215),
.C(n_1202),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1360),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1276),
.A2(n_1097),
.B1(n_1222),
.B2(n_1122),
.Y(n_1453)
);

O2A1O1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1392),
.A2(n_1390),
.B(n_1347),
.C(n_1241),
.Y(n_1454)
);

AOI22x1_ASAP7_75t_L g1455 ( 
.A1(n_1239),
.A2(n_1178),
.B1(n_1159),
.B2(n_1163),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1361),
.B(n_1152),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1235),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1380),
.Y(n_1458)
);

INVxp67_ASAP7_75t_L g1459 ( 
.A(n_1367),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1241),
.B(n_1047),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1262),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1385),
.B(n_1151),
.Y(n_1462)
);

INVxp33_ASAP7_75t_L g1463 ( 
.A(n_1347),
.Y(n_1463)
);

AO21x2_ASAP7_75t_L g1464 ( 
.A1(n_1243),
.A2(n_1152),
.B(n_1202),
.Y(n_1464)
);

INVxp67_ASAP7_75t_L g1465 ( 
.A(n_1244),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1299),
.A2(n_1204),
.B(n_1166),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1397),
.A2(n_1097),
.B1(n_1185),
.B2(n_1166),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1388),
.B(n_1047),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1345),
.B(n_1063),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1374),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1282),
.B(n_1312),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1245),
.A2(n_1204),
.B(n_1166),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1245),
.A2(n_1204),
.B(n_1224),
.Y(n_1473)
);

AO31x2_ASAP7_75t_L g1474 ( 
.A1(n_1236),
.A2(n_1354),
.A3(n_1366),
.B(n_1315),
.Y(n_1474)
);

AND2x2_ASAP7_75t_SL g1475 ( 
.A(n_1237),
.B(n_1097),
.Y(n_1475)
);

AO31x2_ASAP7_75t_L g1476 ( 
.A1(n_1258),
.A2(n_413),
.A3(n_430),
.B(n_401),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1291),
.A2(n_1208),
.B1(n_1221),
.B2(n_1213),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1232),
.A2(n_1313),
.B(n_1311),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1282),
.B(n_1063),
.Y(n_1479)
);

INVx2_ASAP7_75t_SL g1480 ( 
.A(n_1287),
.Y(n_1480)
);

INVx2_ASAP7_75t_SL g1481 ( 
.A(n_1287),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1274),
.B(n_1216),
.Y(n_1482)
);

NAND2xp33_ASAP7_75t_L g1483 ( 
.A(n_1255),
.B(n_1097),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_1312),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1258),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1311),
.A2(n_1224),
.B(n_1192),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1365),
.B(n_1071),
.Y(n_1487)
);

INVx8_ASAP7_75t_L g1488 ( 
.A(n_1357),
.Y(n_1488)
);

BUFx12f_ASAP7_75t_L g1489 ( 
.A(n_1348),
.Y(n_1489)
);

BUFx12f_ASAP7_75t_L g1490 ( 
.A(n_1365),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1273),
.Y(n_1491)
);

OAI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1238),
.A2(n_1150),
.B(n_1215),
.Y(n_1492)
);

CKINVDCx11_ASAP7_75t_R g1493 ( 
.A(n_1277),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1313),
.A2(n_1224),
.B(n_409),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1252),
.B(n_1071),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1242),
.A2(n_1150),
.B(n_1097),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1277),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1273),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_1384),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1305),
.A2(n_1150),
.B1(n_1213),
.B2(n_1048),
.Y(n_1500)
);

BUFx6f_ASAP7_75t_L g1501 ( 
.A(n_1287),
.Y(n_1501)
);

INVx3_ASAP7_75t_L g1502 ( 
.A(n_1319),
.Y(n_1502)
);

AOI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1309),
.A2(n_1144),
.B(n_1119),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1275),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1396),
.Y(n_1505)
);

OA21x2_ASAP7_75t_L g1506 ( 
.A1(n_1306),
.A2(n_409),
.B(n_406),
.Y(n_1506)
);

AOI221xp5_ASAP7_75t_L g1507 ( 
.A1(n_1368),
.A2(n_1048),
.B1(n_471),
.B2(n_454),
.C(n_448),
.Y(n_1507)
);

OA21x2_ASAP7_75t_L g1508 ( 
.A1(n_1306),
.A2(n_429),
.B(n_406),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1246),
.A2(n_1262),
.B1(n_1331),
.B2(n_1284),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1275),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1314),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1342),
.B(n_1168),
.Y(n_1512)
);

CKINVDCx14_ASAP7_75t_R g1513 ( 
.A(n_1338),
.Y(n_1513)
);

AND2x6_ASAP7_75t_L g1514 ( 
.A(n_1287),
.B(n_1224),
.Y(n_1514)
);

A2O1A1Ixp33_ASAP7_75t_L g1515 ( 
.A1(n_1307),
.A2(n_1053),
.B(n_1050),
.C(n_1057),
.Y(n_1515)
);

OAI21x1_ASAP7_75t_L g1516 ( 
.A1(n_1247),
.A2(n_430),
.B(n_429),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1314),
.Y(n_1517)
);

CKINVDCx20_ASAP7_75t_R g1518 ( 
.A(n_1364),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1387),
.Y(n_1519)
);

BUFx2_ASAP7_75t_L g1520 ( 
.A(n_1262),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1247),
.A2(n_454),
.B(n_448),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1271),
.A2(n_471),
.B(n_1150),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1292),
.B(n_1144),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_SL g1524 ( 
.A(n_1292),
.B(n_1191),
.Y(n_1524)
);

NAND2x1p5_ASAP7_75t_L g1525 ( 
.A(n_1319),
.B(n_1191),
.Y(n_1525)
);

OAI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1261),
.A2(n_1082),
.B1(n_1050),
.B2(n_1053),
.Y(n_1526)
);

BUFx2_ASAP7_75t_L g1527 ( 
.A(n_1256),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1399),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1272),
.A2(n_1191),
.B1(n_1155),
.B2(n_1163),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1319),
.Y(n_1530)
);

AO31x2_ASAP7_75t_L g1531 ( 
.A1(n_1318),
.A2(n_1150),
.A3(n_857),
.B(n_1216),
.Y(n_1531)
);

AOI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1295),
.A2(n_1159),
.B(n_1155),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1318),
.Y(n_1533)
);

INVx4_ASAP7_75t_SL g1534 ( 
.A(n_1382),
.Y(n_1534)
);

OAI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1307),
.A2(n_857),
.B(n_1200),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1271),
.A2(n_1159),
.B(n_1155),
.Y(n_1536)
);

OA21x2_ASAP7_75t_L g1537 ( 
.A1(n_1353),
.A2(n_1386),
.B(n_1378),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_1256),
.Y(n_1538)
);

INVx4_ASAP7_75t_L g1539 ( 
.A(n_1387),
.Y(n_1539)
);

OAI21x1_ASAP7_75t_L g1540 ( 
.A1(n_1268),
.A2(n_1163),
.B(n_1053),
.Y(n_1540)
);

INVx2_ASAP7_75t_SL g1541 ( 
.A(n_1387),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1373),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1376),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1358),
.A2(n_281),
.B1(n_857),
.B2(n_1216),
.Y(n_1544)
);

OAI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1250),
.A2(n_1200),
.B(n_690),
.Y(n_1545)
);

BUFx6f_ASAP7_75t_L g1546 ( 
.A(n_1395),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1381),
.Y(n_1547)
);

INVxp67_ASAP7_75t_SL g1548 ( 
.A(n_1289),
.Y(n_1548)
);

OAI221xp5_ASAP7_75t_L g1549 ( 
.A1(n_1344),
.A2(n_1050),
.B1(n_1053),
.B2(n_1089),
.C(n_1082),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1382),
.Y(n_1550)
);

NAND2x1p5_ASAP7_75t_L g1551 ( 
.A(n_1320),
.B(n_1057),
.Y(n_1551)
);

BUFx3_ASAP7_75t_L g1552 ( 
.A(n_1395),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1257),
.Y(n_1553)
);

NAND2x1p5_ASAP7_75t_L g1554 ( 
.A(n_1320),
.B(n_1057),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1372),
.A2(n_281),
.B1(n_1216),
.B2(n_1089),
.Y(n_1555)
);

OAI21x1_ASAP7_75t_L g1556 ( 
.A1(n_1268),
.A2(n_1163),
.B(n_1082),
.Y(n_1556)
);

OAI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1305),
.A2(n_265),
.B(n_259),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1357),
.B(n_1057),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1257),
.A2(n_1089),
.B(n_1082),
.Y(n_1559)
);

NOR2x1_ASAP7_75t_SL g1560 ( 
.A(n_1320),
.B(n_1089),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1256),
.Y(n_1561)
);

OA21x2_ASAP7_75t_L g1562 ( 
.A1(n_1353),
.A2(n_267),
.B(n_266),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1259),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1265),
.A2(n_835),
.B(n_650),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1382),
.Y(n_1565)
);

AO21x2_ASAP7_75t_L g1566 ( 
.A1(n_1378),
.A2(n_346),
.B(n_835),
.Y(n_1566)
);

OAI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1251),
.A2(n_299),
.B(n_292),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1265),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1298),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1372),
.A2(n_317),
.B1(n_328),
.B2(n_344),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1298),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1382),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1300),
.A2(n_328),
.B1(n_470),
.B2(n_464),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1370),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1357),
.B(n_835),
.Y(n_1575)
);

AOI21xp33_ASAP7_75t_SL g1576 ( 
.A1(n_1296),
.A2(n_11),
.B(n_12),
.Y(n_1576)
);

AO21x2_ASAP7_75t_L g1577 ( 
.A1(n_1386),
.A2(n_346),
.B(n_835),
.Y(n_1577)
);

CKINVDCx20_ASAP7_75t_R g1578 ( 
.A(n_1259),
.Y(n_1578)
);

INVx6_ASAP7_75t_SL g1579 ( 
.A(n_1377),
.Y(n_1579)
);

OAI21x1_ASAP7_75t_L g1580 ( 
.A1(n_1254),
.A2(n_650),
.B(n_746),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1298),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1298),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1377),
.B(n_108),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1253),
.B(n_650),
.Y(n_1584)
);

AOI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1483),
.A2(n_1325),
.B(n_1296),
.Y(n_1585)
);

OR2x6_ASAP7_75t_L g1586 ( 
.A(n_1496),
.B(n_1413),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1420),
.A2(n_1254),
.B(n_1283),
.Y(n_1587)
);

OAI22x1_ASAP7_75t_L g1588 ( 
.A1(n_1500),
.A2(n_1371),
.B1(n_1389),
.B2(n_1317),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1488),
.Y(n_1589)
);

NAND3xp33_ASAP7_75t_SL g1590 ( 
.A(n_1454),
.B(n_307),
.C(n_304),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1453),
.A2(n_1391),
.B1(n_1343),
.B2(n_1346),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1493),
.Y(n_1592)
);

A2O1A1Ixp33_ASAP7_75t_L g1593 ( 
.A1(n_1437),
.A2(n_1362),
.B(n_1294),
.C(n_1285),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1402),
.B(n_1259),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1459),
.B(n_1383),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1406),
.Y(n_1596)
);

AOI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1483),
.A2(n_1325),
.B(n_1316),
.Y(n_1597)
);

AOI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1518),
.A2(n_1395),
.B1(n_1377),
.B2(n_1355),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1463),
.B(n_1383),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1451),
.A2(n_1308),
.B1(n_470),
.B2(n_439),
.Y(n_1600)
);

AND2x4_ASAP7_75t_L g1601 ( 
.A(n_1402),
.B(n_1269),
.Y(n_1601)
);

AOI221xp5_ASAP7_75t_L g1602 ( 
.A1(n_1411),
.A2(n_1336),
.B1(n_317),
.B2(n_328),
.C(n_344),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1408),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1542),
.B(n_1383),
.Y(n_1604)
);

OAI221xp5_ASAP7_75t_L g1605 ( 
.A1(n_1507),
.A2(n_1334),
.B1(n_1335),
.B2(n_1330),
.C(n_1326),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1543),
.B(n_1547),
.Y(n_1606)
);

INVx1_ASAP7_75t_SL g1607 ( 
.A(n_1484),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1463),
.B(n_1383),
.Y(n_1608)
);

OR2x6_ASAP7_75t_L g1609 ( 
.A(n_1413),
.B(n_1289),
.Y(n_1609)
);

INVx3_ASAP7_75t_L g1610 ( 
.A(n_1488),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1401),
.Y(n_1611)
);

AO21x2_ASAP7_75t_L g1612 ( 
.A1(n_1403),
.A2(n_1327),
.B(n_1329),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1518),
.A2(n_439),
.B1(n_317),
.B2(n_328),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1421),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1447),
.B(n_1269),
.Y(n_1615)
);

NAND3xp33_ASAP7_75t_L g1616 ( 
.A(n_1557),
.B(n_344),
.C(n_328),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1456),
.B(n_12),
.Y(n_1617)
);

AO221x2_ASAP7_75t_L g1618 ( 
.A1(n_1448),
.A2(n_14),
.B1(n_15),
.B2(n_20),
.C(n_21),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1475),
.A2(n_470),
.B1(n_464),
.B2(n_439),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1460),
.B(n_1269),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1449),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1475),
.A2(n_439),
.B1(n_344),
.B2(n_464),
.Y(n_1622)
);

AO22x1_ASAP7_75t_SL g1623 ( 
.A1(n_1402),
.A2(n_1317),
.B1(n_22),
.B2(n_23),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1452),
.Y(n_1624)
);

INVx4_ASAP7_75t_SL g1625 ( 
.A(n_1514),
.Y(n_1625)
);

OAI211xp5_ASAP7_75t_SL g1626 ( 
.A1(n_1465),
.A2(n_1379),
.B(n_1394),
.C(n_1393),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1578),
.Y(n_1627)
);

O2A1O1Ixp33_ASAP7_75t_SL g1628 ( 
.A1(n_1492),
.A2(n_1248),
.B(n_1316),
.C(n_1304),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1409),
.Y(n_1629)
);

NAND2xp33_ASAP7_75t_SL g1630 ( 
.A(n_1538),
.B(n_1340),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1458),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_SL g1632 ( 
.A1(n_1464),
.A2(n_1317),
.B1(n_464),
.B2(n_470),
.Y(n_1632)
);

AND2x4_ASAP7_75t_L g1633 ( 
.A(n_1426),
.B(n_1431),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1427),
.Y(n_1634)
);

BUFx2_ASAP7_75t_L g1635 ( 
.A(n_1578),
.Y(n_1635)
);

CKINVDCx20_ASAP7_75t_R g1636 ( 
.A(n_1493),
.Y(n_1636)
);

OAI221xp5_ASAP7_75t_L g1637 ( 
.A1(n_1430),
.A2(n_1424),
.B1(n_1477),
.B2(n_1432),
.C(n_1469),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1425),
.Y(n_1638)
);

AOI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1466),
.A2(n_1322),
.B(n_1304),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_1499),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1433),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1456),
.B(n_15),
.Y(n_1642)
);

CKINVDCx11_ASAP7_75t_R g1643 ( 
.A(n_1425),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1446),
.B(n_1461),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1471),
.B(n_1340),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1505),
.Y(n_1646)
);

INVx6_ASAP7_75t_L g1647 ( 
.A(n_1490),
.Y(n_1647)
);

OAI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1443),
.A2(n_1398),
.B1(n_1340),
.B2(n_1321),
.Y(n_1648)
);

BUFx2_ASAP7_75t_L g1649 ( 
.A(n_1490),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1467),
.A2(n_1464),
.B1(n_1512),
.B2(n_1412),
.Y(n_1650)
);

INVx6_ASAP7_75t_L g1651 ( 
.A(n_1488),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1528),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1485),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1485),
.Y(n_1654)
);

INVx3_ASAP7_75t_L g1655 ( 
.A(n_1488),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1499),
.B(n_1398),
.Y(n_1656)
);

INVx3_ASAP7_75t_L g1657 ( 
.A(n_1539),
.Y(n_1657)
);

NAND2x1p5_ASAP7_75t_L g1658 ( 
.A(n_1523),
.B(n_1398),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1498),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1429),
.A2(n_1321),
.B1(n_1322),
.B2(n_1333),
.Y(n_1660)
);

OAI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1446),
.A2(n_1520),
.B1(n_1461),
.B2(n_1576),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1427),
.Y(n_1662)
);

OAI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1520),
.A2(n_344),
.B1(n_439),
.B2(n_464),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1431),
.B(n_23),
.Y(n_1664)
);

OAI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1567),
.A2(n_470),
.B1(n_1363),
.B2(n_1317),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1513),
.A2(n_325),
.B1(n_319),
.B2(n_312),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1464),
.A2(n_1412),
.B1(n_1416),
.B2(n_1403),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1498),
.Y(n_1668)
);

AOI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1441),
.A2(n_1267),
.B1(n_329),
.B2(n_396),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1491),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1426),
.A2(n_1267),
.B1(n_460),
.B2(n_1323),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1482),
.B(n_1301),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1489),
.Y(n_1673)
);

INVx3_ASAP7_75t_L g1674 ( 
.A(n_1539),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_1489),
.Y(n_1675)
);

AO21x2_ASAP7_75t_L g1676 ( 
.A1(n_1550),
.A2(n_1323),
.B(n_1283),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1431),
.B(n_28),
.Y(n_1677)
);

AOI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1509),
.A2(n_331),
.B1(n_334),
.B2(n_335),
.C(n_338),
.Y(n_1678)
);

CKINVDCx16_ASAP7_75t_R g1679 ( 
.A(n_1497),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1445),
.B(n_29),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1457),
.B(n_29),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1426),
.B(n_1290),
.Y(n_1682)
);

NOR3xp33_ASAP7_75t_SL g1683 ( 
.A(n_1538),
.B(n_1487),
.C(n_1479),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1513),
.B(n_30),
.Y(n_1684)
);

OAI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1468),
.A2(n_342),
.B1(n_343),
.B2(n_347),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1482),
.B(n_1301),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1497),
.Y(n_1687)
);

INVx3_ASAP7_75t_L g1688 ( 
.A(n_1539),
.Y(n_1688)
);

NOR3xp33_ASAP7_75t_SL g1689 ( 
.A(n_1526),
.B(n_352),
.C(n_359),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1495),
.B(n_30),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_SL g1691 ( 
.A1(n_1450),
.A2(n_460),
.B1(n_1290),
.B2(n_1288),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_1579),
.Y(n_1692)
);

AO22x2_ASAP7_75t_L g1693 ( 
.A1(n_1534),
.A2(n_1301),
.B1(n_1288),
.B2(n_34),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1570),
.A2(n_460),
.B1(n_366),
.B2(n_426),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1450),
.A2(n_460),
.B1(n_368),
.B2(n_431),
.Y(n_1695)
);

INVx4_ASAP7_75t_L g1696 ( 
.A(n_1501),
.Y(n_1696)
);

AO31x2_ASAP7_75t_L g1697 ( 
.A1(n_1571),
.A2(n_1582),
.A3(n_1581),
.B(n_1569),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1504),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1504),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_SL g1700 ( 
.A1(n_1450),
.A2(n_437),
.B1(n_387),
.B2(n_394),
.Y(n_1700)
);

INVx3_ASAP7_75t_SL g1701 ( 
.A(n_1523),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1433),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1552),
.B(n_31),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1565),
.A2(n_466),
.B1(n_422),
.B2(n_423),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1552),
.B(n_32),
.Y(n_1705)
);

OR2x6_ASAP7_75t_L g1706 ( 
.A(n_1583),
.B(n_1301),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1519),
.Y(n_1707)
);

AOI21xp33_ASAP7_75t_L g1708 ( 
.A1(n_1444),
.A2(n_376),
.B(n_424),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_1523),
.B(n_34),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1510),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1572),
.A2(n_1574),
.B1(n_1534),
.B2(n_1562),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1519),
.B(n_37),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1462),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1519),
.B(n_37),
.Y(n_1714)
);

CKINVDCx20_ASAP7_75t_R g1715 ( 
.A(n_1563),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_1579),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1534),
.A2(n_452),
.B1(n_746),
.B2(n_716),
.Y(n_1717)
);

A2O1A1Ixp33_ASAP7_75t_L g1718 ( 
.A1(n_1583),
.A2(n_38),
.B(n_42),
.C(n_44),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_SL g1719 ( 
.A(n_1583),
.B(n_716),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1527),
.B(n_1561),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1433),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1555),
.A2(n_38),
.B1(n_45),
.B2(n_47),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1511),
.Y(n_1723)
);

AOI22xp33_ASAP7_75t_SL g1724 ( 
.A1(n_1444),
.A2(n_765),
.B1(n_746),
.B2(n_716),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1541),
.B(n_45),
.Y(n_1725)
);

INVx3_ASAP7_75t_L g1726 ( 
.A(n_1519),
.Y(n_1726)
);

OAI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1535),
.A2(n_1544),
.B1(n_1444),
.B2(n_1545),
.C(n_1573),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1546),
.B(n_51),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1546),
.B(n_52),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1546),
.B(n_1541),
.Y(n_1730)
);

OAI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1532),
.A2(n_765),
.B(n_746),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1549),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1546),
.B(n_54),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1517),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1546),
.B(n_57),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1558),
.B(n_59),
.Y(n_1736)
);

OAI22xp33_ASAP7_75t_L g1737 ( 
.A1(n_1584),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1558),
.B(n_69),
.Y(n_1738)
);

NAND3xp33_ASAP7_75t_SL g1739 ( 
.A(n_1515),
.B(n_1561),
.C(n_1527),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1558),
.B(n_70),
.Y(n_1740)
);

INVx4_ASAP7_75t_L g1741 ( 
.A(n_1501),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1480),
.B(n_1481),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1476),
.B(n_71),
.Y(n_1743)
);

BUFx2_ASAP7_75t_L g1744 ( 
.A(n_1501),
.Y(n_1744)
);

NAND2x1p5_ASAP7_75t_L g1745 ( 
.A(n_1524),
.B(n_765),
.Y(n_1745)
);

AOI211xp5_ASAP7_75t_L g1746 ( 
.A1(n_1529),
.A2(n_71),
.B(n_72),
.C(n_74),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1548),
.B(n_75),
.Y(n_1747)
);

OAI221xp5_ASAP7_75t_L g1748 ( 
.A1(n_1562),
.A2(n_765),
.B1(n_746),
.B2(n_716),
.C(n_78),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1433),
.B(n_75),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1480),
.B(n_76),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1517),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1481),
.B(n_77),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1533),
.Y(n_1753)
);

OAI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1415),
.A2(n_77),
.B1(n_79),
.B2(n_81),
.Y(n_1754)
);

OAI221xp5_ASAP7_75t_L g1755 ( 
.A1(n_1562),
.A2(n_765),
.B1(n_716),
.B2(n_86),
.C(n_90),
.Y(n_1755)
);

CKINVDCx6p67_ASAP7_75t_R g1756 ( 
.A(n_1501),
.Y(n_1756)
);

AOI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1534),
.A2(n_1419),
.B1(n_1569),
.B2(n_1579),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_SL g1758 ( 
.A1(n_1419),
.A2(n_83),
.B1(n_84),
.B2(n_86),
.Y(n_1758)
);

BUFx2_ASAP7_75t_L g1759 ( 
.A(n_1501),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1533),
.B(n_84),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1433),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1476),
.Y(n_1762)
);

NAND2xp33_ASAP7_75t_SL g1763 ( 
.A(n_1415),
.B(n_91),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1476),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1571),
.Y(n_1765)
);

OAI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1405),
.A2(n_91),
.B1(n_92),
.B2(n_94),
.Y(n_1766)
);

OAI221xp5_ASAP7_75t_L g1767 ( 
.A1(n_1455),
.A2(n_92),
.B1(n_96),
.B2(n_97),
.C(n_98),
.Y(n_1767)
);

NAND3xp33_ASAP7_75t_L g1768 ( 
.A(n_1455),
.B(n_97),
.C(n_98),
.Y(n_1768)
);

NAND2xp33_ASAP7_75t_SL g1769 ( 
.A(n_1415),
.B(n_100),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1419),
.A2(n_101),
.B1(n_105),
.B2(n_106),
.Y(n_1770)
);

INVx6_ASAP7_75t_L g1771 ( 
.A(n_1575),
.Y(n_1771)
);

AOI211x1_ASAP7_75t_L g1772 ( 
.A1(n_1442),
.A2(n_105),
.B(n_115),
.C(n_116),
.Y(n_1772)
);

BUFx12f_ASAP7_75t_L g1773 ( 
.A(n_1410),
.Y(n_1773)
);

BUFx3_ASAP7_75t_L g1774 ( 
.A(n_1514),
.Y(n_1774)
);

AOI221xp5_ASAP7_75t_L g1775 ( 
.A1(n_1423),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.C(n_124),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1476),
.B(n_129),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1410),
.B(n_238),
.Y(n_1777)
);

BUFx3_ASAP7_75t_L g1778 ( 
.A(n_1514),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1476),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1407),
.A2(n_130),
.B1(n_133),
.B2(n_134),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1581),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1400),
.Y(n_1782)
);

OAI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1551),
.A2(n_1554),
.B1(n_1502),
.B2(n_1530),
.Y(n_1783)
);

OAI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1551),
.A2(n_148),
.B1(n_150),
.B2(n_151),
.Y(n_1784)
);

INVx2_ASAP7_75t_SL g1785 ( 
.A(n_1410),
.Y(n_1785)
);

AOI221xp5_ASAP7_75t_L g1786 ( 
.A1(n_1423),
.A2(n_153),
.B1(n_156),
.B2(n_159),
.C(n_161),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_SL g1787 ( 
.A1(n_1618),
.A2(n_1577),
.B1(n_1566),
.B2(n_1407),
.Y(n_1787)
);

NAND3xp33_ASAP7_75t_SL g1788 ( 
.A(n_1746),
.B(n_1438),
.C(n_1554),
.Y(n_1788)
);

OAI221xp5_ASAP7_75t_L g1789 ( 
.A1(n_1613),
.A2(n_1506),
.B1(n_1508),
.B2(n_1404),
.C(n_1438),
.Y(n_1789)
);

OAI21xp33_ASAP7_75t_SL g1790 ( 
.A1(n_1770),
.A2(n_1472),
.B(n_1440),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1618),
.A2(n_1407),
.B1(n_1423),
.B2(n_1577),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1627),
.B(n_1531),
.Y(n_1792)
);

OAI221xp5_ASAP7_75t_L g1793 ( 
.A1(n_1613),
.A2(n_1508),
.B1(n_1506),
.B2(n_1404),
.C(n_1551),
.Y(n_1793)
);

OAI221xp5_ASAP7_75t_L g1794 ( 
.A1(n_1718),
.A2(n_1506),
.B1(n_1508),
.B2(n_1404),
.C(n_1553),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_SL g1795 ( 
.A1(n_1618),
.A2(n_1566),
.B1(n_1577),
.B2(n_1472),
.Y(n_1795)
);

CKINVDCx20_ASAP7_75t_R g1796 ( 
.A(n_1636),
.Y(n_1796)
);

AOI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1749),
.A2(n_1566),
.B1(n_1582),
.B2(n_1537),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1602),
.A2(n_1619),
.B1(n_1622),
.B2(n_1770),
.Y(n_1798)
);

AOI221xp5_ASAP7_75t_L g1799 ( 
.A1(n_1737),
.A2(n_1695),
.B1(n_1766),
.B2(n_1637),
.C(n_1590),
.Y(n_1799)
);

AOI221xp5_ASAP7_75t_L g1800 ( 
.A1(n_1737),
.A2(n_1568),
.B1(n_1553),
.B2(n_1435),
.C(n_1470),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1596),
.Y(n_1801)
);

OAI211xp5_ASAP7_75t_L g1802 ( 
.A1(n_1669),
.A2(n_1690),
.B(n_1695),
.C(n_1767),
.Y(n_1802)
);

OR2x6_ASAP7_75t_L g1803 ( 
.A(n_1706),
.B(n_1473),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1630),
.A2(n_1769),
.B(n_1763),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1635),
.B(n_1531),
.Y(n_1805)
);

AOI211xp5_ASAP7_75t_L g1806 ( 
.A1(n_1766),
.A2(n_1521),
.B(n_1516),
.C(n_1503),
.Y(n_1806)
);

A2O1A1Ixp33_ASAP7_75t_L g1807 ( 
.A1(n_1619),
.A2(n_1473),
.B(n_1522),
.C(n_1516),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1617),
.B(n_1642),
.Y(n_1808)
);

AOI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1763),
.A2(n_1439),
.B(n_1560),
.Y(n_1809)
);

AOI222xp33_ASAP7_75t_L g1810 ( 
.A1(n_1622),
.A2(n_1575),
.B1(n_1514),
.B2(n_1435),
.C1(n_1470),
.C2(n_1560),
.Y(n_1810)
);

OAI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1690),
.A2(n_1502),
.B1(n_1530),
.B2(n_1525),
.Y(n_1811)
);

OAI221xp5_ASAP7_75t_L g1812 ( 
.A1(n_1758),
.A2(n_1568),
.B1(n_1439),
.B2(n_1537),
.C(n_1525),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1664),
.B(n_1531),
.Y(n_1813)
);

BUFx3_ASAP7_75t_L g1814 ( 
.A(n_1649),
.Y(n_1814)
);

AND2x2_ASAP7_75t_SL g1815 ( 
.A(n_1641),
.B(n_1439),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1677),
.B(n_1531),
.Y(n_1816)
);

OAI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1700),
.A2(n_1600),
.B1(n_1715),
.B2(n_1661),
.Y(n_1817)
);

AOI222xp33_ASAP7_75t_L g1818 ( 
.A1(n_1650),
.A2(n_1575),
.B1(n_1514),
.B2(n_1522),
.C1(n_1521),
.C2(n_1417),
.Y(n_1818)
);

HB1xp67_ASAP7_75t_L g1819 ( 
.A(n_1782),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1615),
.B(n_1400),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1603),
.Y(n_1821)
);

OAI211xp5_ASAP7_75t_L g1822 ( 
.A1(n_1769),
.A2(n_1440),
.B(n_1494),
.C(n_1422),
.Y(n_1822)
);

OR2x6_ASAP7_75t_L g1823 ( 
.A(n_1706),
.B(n_1486),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_SL g1824 ( 
.A1(n_1623),
.A2(n_1514),
.B1(n_1537),
.B2(n_1418),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1606),
.B(n_1400),
.Y(n_1825)
);

INVx2_ASAP7_75t_SL g1826 ( 
.A(n_1647),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1652),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_L g1828 ( 
.A1(n_1632),
.A2(n_1418),
.B1(n_1414),
.B2(n_1417),
.Y(n_1828)
);

HB1xp67_ASAP7_75t_L g1829 ( 
.A(n_1676),
.Y(n_1829)
);

HB1xp67_ASAP7_75t_L g1830 ( 
.A(n_1676),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1614),
.Y(n_1831)
);

NOR4xp25_ASAP7_75t_L g1832 ( 
.A(n_1754),
.B(n_1474),
.C(n_1400),
.D(n_1494),
.Y(n_1832)
);

O2A1O1Ixp33_ASAP7_75t_L g1833 ( 
.A1(n_1732),
.A2(n_1722),
.B(n_1684),
.C(n_1661),
.Y(n_1833)
);

AOI33xp33_ASAP7_75t_L g1834 ( 
.A1(n_1680),
.A2(n_1474),
.A3(n_1400),
.B1(n_170),
.B2(n_174),
.B3(n_182),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1644),
.B(n_1474),
.Y(n_1835)
);

OAI21x1_ASAP7_75t_L g1836 ( 
.A1(n_1587),
.A2(n_1478),
.B(n_1580),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1703),
.B(n_1486),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1621),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1705),
.B(n_1536),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1624),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_SL g1841 ( 
.A1(n_1719),
.A2(n_1559),
.B1(n_1536),
.B2(n_1414),
.Y(n_1841)
);

OAI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1709),
.A2(n_1434),
.B1(n_1436),
.B2(n_1422),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1709),
.B(n_1559),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1631),
.Y(n_1844)
);

NAND3xp33_ASAP7_75t_L g1845 ( 
.A(n_1678),
.B(n_1474),
.C(n_1428),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1738),
.B(n_1556),
.Y(n_1846)
);

NOR2x1_ASAP7_75t_R g1847 ( 
.A(n_1643),
.B(n_162),
.Y(n_1847)
);

OAI221xp5_ASAP7_75t_L g1848 ( 
.A1(n_1708),
.A2(n_1474),
.B1(n_1428),
.B2(n_1436),
.C(n_1556),
.Y(n_1848)
);

AOI221x1_ASAP7_75t_SL g1849 ( 
.A1(n_1681),
.A2(n_163),
.B1(n_186),
.B2(n_191),
.C(n_196),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1620),
.B(n_1540),
.Y(n_1850)
);

INVx3_ASAP7_75t_L g1851 ( 
.A(n_1696),
.Y(n_1851)
);

AOI22xp33_ASAP7_75t_SL g1852 ( 
.A1(n_1616),
.A2(n_1540),
.B1(n_1564),
.B2(n_209),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1720),
.B(n_1564),
.Y(n_1853)
);

AOI21xp33_ASAP7_75t_L g1854 ( 
.A1(n_1588),
.A2(n_1755),
.B(n_1604),
.Y(n_1854)
);

OAI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1743),
.A2(n_205),
.B1(n_206),
.B2(n_218),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1650),
.A2(n_222),
.B1(n_232),
.B2(n_1599),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1670),
.Y(n_1857)
);

OAI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1598),
.A2(n_1586),
.B1(n_1701),
.B2(n_1665),
.Y(n_1858)
);

HB1xp67_ASAP7_75t_L g1859 ( 
.A(n_1641),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1738),
.A2(n_1740),
.B1(n_1736),
.B2(n_1713),
.Y(n_1860)
);

NOR2xp33_ASAP7_75t_L g1861 ( 
.A(n_1714),
.B(n_1736),
.Y(n_1861)
);

INVx2_ASAP7_75t_SL g1862 ( 
.A(n_1647),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1653),
.Y(n_1863)
);

HB1xp67_ASAP7_75t_L g1864 ( 
.A(n_1702),
.Y(n_1864)
);

CKINVDCx14_ASAP7_75t_R g1865 ( 
.A(n_1643),
.Y(n_1865)
);

NAND3xp33_ASAP7_75t_L g1866 ( 
.A(n_1775),
.B(n_1786),
.C(n_1772),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1608),
.A2(n_1776),
.B1(n_1595),
.B2(n_1780),
.Y(n_1867)
);

OAI21x1_ASAP7_75t_L g1868 ( 
.A1(n_1597),
.A2(n_1585),
.B(n_1671),
.Y(n_1868)
);

OAI22xp33_ASAP7_75t_L g1869 ( 
.A1(n_1586),
.A2(n_1701),
.B1(n_1768),
.B2(n_1747),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1654),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_SL g1871 ( 
.A1(n_1702),
.A2(n_1761),
.B1(n_1721),
.B2(n_1693),
.Y(n_1871)
);

AOI22xp33_ASAP7_75t_SL g1872 ( 
.A1(n_1721),
.A2(n_1761),
.B1(n_1693),
.B2(n_1748),
.Y(n_1872)
);

OAI22xp33_ASAP7_75t_L g1873 ( 
.A1(n_1586),
.A2(n_1784),
.B1(n_1727),
.B2(n_1740),
.Y(n_1873)
);

BUFx3_ASAP7_75t_L g1874 ( 
.A(n_1647),
.Y(n_1874)
);

AOI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_1780),
.A2(n_1667),
.B1(n_1693),
.B2(n_1694),
.Y(n_1875)
);

OAI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1683),
.A2(n_1704),
.B1(n_1640),
.B2(n_1714),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1712),
.B(n_1728),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_SL g1878 ( 
.A(n_1783),
.B(n_1683),
.Y(n_1878)
);

OAI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1704),
.A2(n_1675),
.B1(n_1673),
.B2(n_1591),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1659),
.Y(n_1880)
);

AOI221xp5_ASAP7_75t_L g1881 ( 
.A1(n_1667),
.A2(n_1666),
.B1(n_1711),
.B2(n_1784),
.C(n_1663),
.Y(n_1881)
);

OAI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1591),
.A2(n_1656),
.B1(n_1733),
.B2(n_1735),
.Y(n_1882)
);

A2O1A1Ixp33_ASAP7_75t_L g1883 ( 
.A1(n_1593),
.A2(n_1689),
.B(n_1671),
.C(n_1691),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1694),
.A2(n_1711),
.B1(n_1605),
.B2(n_1706),
.Y(n_1884)
);

OAI221xp5_ASAP7_75t_L g1885 ( 
.A1(n_1689),
.A2(n_1593),
.B1(n_1607),
.B2(n_1725),
.C(n_1685),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_SL g1886 ( 
.A1(n_1774),
.A2(n_1778),
.B1(n_1773),
.B2(n_1771),
.Y(n_1886)
);

BUFx3_ASAP7_75t_L g1887 ( 
.A(n_1687),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1762),
.A2(n_1779),
.B1(n_1764),
.B2(n_1686),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1672),
.B(n_1668),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1698),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1699),
.Y(n_1891)
);

OAI332xp33_ASAP7_75t_L g1892 ( 
.A1(n_1750),
.A2(n_1752),
.A3(n_1760),
.B1(n_1679),
.B2(n_1645),
.B3(n_1785),
.C1(n_1777),
.C2(n_1660),
.Y(n_1892)
);

OAI22xp33_ASAP7_75t_L g1893 ( 
.A1(n_1774),
.A2(n_1778),
.B1(n_1651),
.B2(n_1773),
.Y(n_1893)
);

AOI22xp33_ASAP7_75t_SL g1894 ( 
.A1(n_1771),
.A2(n_1729),
.B1(n_1651),
.B2(n_1682),
.Y(n_1894)
);

OAI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1657),
.A2(n_1674),
.B1(n_1688),
.B2(n_1589),
.Y(n_1895)
);

AOI22xp33_ASAP7_75t_SL g1896 ( 
.A1(n_1771),
.A2(n_1651),
.B1(n_1633),
.B2(n_1648),
.Y(n_1896)
);

AOI22xp33_ASAP7_75t_L g1897 ( 
.A1(n_1594),
.A2(n_1601),
.B1(n_1633),
.B2(n_1739),
.Y(n_1897)
);

OAI21xp5_ASAP7_75t_L g1898 ( 
.A1(n_1639),
.A2(n_1626),
.B(n_1628),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1730),
.B(n_1594),
.Y(n_1899)
);

OAI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1657),
.A2(n_1674),
.B1(n_1688),
.B2(n_1589),
.Y(n_1900)
);

OAI22xp33_ASAP7_75t_L g1901 ( 
.A1(n_1609),
.A2(n_1716),
.B1(n_1692),
.B2(n_1655),
.Y(n_1901)
);

AOI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1628),
.A2(n_1783),
.B(n_1609),
.Y(n_1902)
);

AOI22xp33_ASAP7_75t_SL g1903 ( 
.A1(n_1601),
.A2(n_1707),
.B1(n_1609),
.B2(n_1655),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1726),
.B(n_1744),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1742),
.B(n_1726),
.Y(n_1905)
);

AOI221xp5_ASAP7_75t_L g1906 ( 
.A1(n_1757),
.A2(n_1638),
.B1(n_1753),
.B2(n_1717),
.C(n_1612),
.Y(n_1906)
);

AOI22xp33_ASAP7_75t_L g1907 ( 
.A1(n_1717),
.A2(n_1757),
.B1(n_1723),
.B2(n_1751),
.Y(n_1907)
);

AOI222xp33_ASAP7_75t_L g1908 ( 
.A1(n_1625),
.A2(n_1723),
.B1(n_1710),
.B2(n_1751),
.C1(n_1734),
.C2(n_1611),
.Y(n_1908)
);

OAI221xp5_ASAP7_75t_L g1909 ( 
.A1(n_1658),
.A2(n_1610),
.B1(n_1759),
.B2(n_1724),
.C(n_1592),
.Y(n_1909)
);

OAI221xp5_ASAP7_75t_L g1910 ( 
.A1(n_1610),
.A2(n_1745),
.B1(n_1741),
.B2(n_1731),
.C(n_1734),
.Y(n_1910)
);

AOI22xp33_ASAP7_75t_L g1911 ( 
.A1(n_1710),
.A2(n_1781),
.B1(n_1765),
.B2(n_1629),
.Y(n_1911)
);

AOI211xp5_ASAP7_75t_SL g1912 ( 
.A1(n_1765),
.A2(n_1781),
.B(n_1629),
.C(n_1634),
.Y(n_1912)
);

AOI21xp5_ASAP7_75t_SL g1913 ( 
.A1(n_1662),
.A2(n_1718),
.B(n_1618),
.Y(n_1913)
);

AOI22xp33_ASAP7_75t_L g1914 ( 
.A1(n_1697),
.A2(n_1080),
.B1(n_1618),
.B2(n_1095),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1697),
.B(n_1615),
.Y(n_1915)
);

AOI221xp5_ASAP7_75t_L g1916 ( 
.A1(n_1697),
.A2(n_1095),
.B1(n_866),
.B2(n_1454),
.C(n_1281),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_1643),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1596),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1646),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1627),
.B(n_1635),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_L g1921 ( 
.A1(n_1618),
.A2(n_1080),
.B1(n_1095),
.B2(n_1112),
.Y(n_1921)
);

OAI22xp5_ASAP7_75t_L g1922 ( 
.A1(n_1718),
.A2(n_1069),
.B1(n_1500),
.B2(n_866),
.Y(n_1922)
);

AOI22xp5_ASAP7_75t_L g1923 ( 
.A1(n_1618),
.A2(n_866),
.B1(n_1069),
.B2(n_1095),
.Y(n_1923)
);

AOI22xp33_ASAP7_75t_L g1924 ( 
.A1(n_1618),
.A2(n_1080),
.B1(n_1095),
.B2(n_1112),
.Y(n_1924)
);

A2O1A1Ixp33_ASAP7_75t_L g1925 ( 
.A1(n_1718),
.A2(n_1454),
.B(n_1437),
.C(n_1069),
.Y(n_1925)
);

BUFx3_ASAP7_75t_L g1926 ( 
.A(n_1649),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1627),
.B(n_1635),
.Y(n_1927)
);

AO31x2_ASAP7_75t_L g1928 ( 
.A1(n_1588),
.A2(n_1403),
.A3(n_1665),
.B(n_1762),
.Y(n_1928)
);

OAI22xp5_ASAP7_75t_L g1929 ( 
.A1(n_1718),
.A2(n_1069),
.B1(n_1500),
.B2(n_866),
.Y(n_1929)
);

INVx5_ASAP7_75t_SL g1930 ( 
.A(n_1756),
.Y(n_1930)
);

NAND2x1_ASAP7_75t_L g1931 ( 
.A(n_1785),
.B(n_1696),
.Y(n_1931)
);

AND2x4_ASAP7_75t_L g1932 ( 
.A(n_1625),
.B(n_1682),
.Y(n_1932)
);

CKINVDCx20_ASAP7_75t_R g1933 ( 
.A(n_1636),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1627),
.B(n_1635),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1596),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1596),
.Y(n_1936)
);

OA21x2_ASAP7_75t_L g1937 ( 
.A1(n_1587),
.A2(n_1711),
.B(n_1521),
.Y(n_1937)
);

AOI22xp33_ASAP7_75t_L g1938 ( 
.A1(n_1618),
.A2(n_1080),
.B1(n_1095),
.B2(n_1112),
.Y(n_1938)
);

OAI22xp5_ASAP7_75t_L g1939 ( 
.A1(n_1718),
.A2(n_1069),
.B1(n_1500),
.B2(n_866),
.Y(n_1939)
);

AOI22xp33_ASAP7_75t_L g1940 ( 
.A1(n_1618),
.A2(n_1080),
.B1(n_1095),
.B2(n_1112),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_SL g1941 ( 
.A(n_1661),
.B(n_1509),
.Y(n_1941)
);

AOI22xp33_ASAP7_75t_SL g1942 ( 
.A1(n_1618),
.A2(n_866),
.B1(n_1112),
.B2(n_1411),
.Y(n_1942)
);

AND2x4_ASAP7_75t_L g1943 ( 
.A(n_1625),
.B(n_1682),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1596),
.Y(n_1944)
);

OA21x2_ASAP7_75t_L g1945 ( 
.A1(n_1587),
.A2(n_1711),
.B(n_1521),
.Y(n_1945)
);

AO21x2_ASAP7_75t_L g1946 ( 
.A1(n_1762),
.A2(n_1779),
.B(n_1764),
.Y(n_1946)
);

OAI211xp5_ASAP7_75t_SL g1947 ( 
.A1(n_1640),
.A2(n_1054),
.B(n_1048),
.C(n_1000),
.Y(n_1947)
);

AND2x2_ASAP7_75t_SL g1948 ( 
.A(n_1749),
.B(n_1641),
.Y(n_1948)
);

AOI222xp33_ASAP7_75t_L g1949 ( 
.A1(n_1613),
.A2(n_1008),
.B1(n_1112),
.B2(n_1281),
.C1(n_1411),
.C2(n_484),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1596),
.Y(n_1950)
);

OAI22xp5_ASAP7_75t_L g1951 ( 
.A1(n_1718),
.A2(n_1069),
.B1(n_1500),
.B2(n_866),
.Y(n_1951)
);

AO221x2_ASAP7_75t_L g1952 ( 
.A1(n_1737),
.A2(n_1661),
.B1(n_1766),
.B2(n_1618),
.C(n_1448),
.Y(n_1952)
);

AOI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1618),
.A2(n_866),
.B1(n_1069),
.B2(n_1095),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1615),
.B(n_1606),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1718),
.A2(n_1069),
.B1(n_1500),
.B2(n_866),
.Y(n_1955)
);

AOI22xp33_ASAP7_75t_L g1956 ( 
.A1(n_1618),
.A2(n_1080),
.B1(n_1095),
.B2(n_1112),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1627),
.B(n_1635),
.Y(n_1957)
);

AOI22x1_ASAP7_75t_L g1958 ( 
.A1(n_1640),
.A2(n_750),
.B1(n_766),
.B2(n_755),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1615),
.B(n_1606),
.Y(n_1959)
);

INVxp67_ASAP7_75t_L g1960 ( 
.A(n_1819),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1863),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1954),
.B(n_1959),
.Y(n_1962)
);

NOR2xp67_ASAP7_75t_L g1963 ( 
.A(n_1829),
.B(n_1830),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1815),
.B(n_1835),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1815),
.B(n_1850),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1825),
.B(n_1820),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1829),
.B(n_1830),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1870),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1880),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1948),
.B(n_1792),
.Y(n_1970)
);

AOI22xp33_ASAP7_75t_L g1971 ( 
.A1(n_1952),
.A2(n_1924),
.B1(n_1940),
.B2(n_1938),
.Y(n_1971)
);

BUFx3_ASAP7_75t_L g1972 ( 
.A(n_1932),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1857),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1890),
.Y(n_1974)
);

HB1xp67_ASAP7_75t_L g1975 ( 
.A(n_1819),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1891),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1948),
.B(n_1805),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1915),
.B(n_1801),
.Y(n_1978)
);

AOI22xp33_ASAP7_75t_L g1979 ( 
.A1(n_1952),
.A2(n_1924),
.B1(n_1956),
.B2(n_1921),
.Y(n_1979)
);

NAND4xp25_ASAP7_75t_L g1980 ( 
.A(n_1923),
.B(n_1953),
.C(n_1921),
.D(n_1956),
.Y(n_1980)
);

HB1xp67_ASAP7_75t_L g1981 ( 
.A(n_1859),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1839),
.B(n_1803),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1803),
.B(n_1937),
.Y(n_1983)
);

AND2x4_ASAP7_75t_L g1984 ( 
.A(n_1932),
.B(n_1943),
.Y(n_1984)
);

AND2x4_ASAP7_75t_L g1985 ( 
.A(n_1943),
.B(n_1803),
.Y(n_1985)
);

INVxp67_ASAP7_75t_L g1986 ( 
.A(n_1859),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1937),
.B(n_1945),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1937),
.B(n_1945),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1945),
.B(n_1843),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1864),
.B(n_1821),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1864),
.B(n_1831),
.Y(n_1991)
);

BUFx3_ASAP7_75t_L g1992 ( 
.A(n_1931),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1838),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1901),
.B(n_1893),
.Y(n_1994)
);

OAI221xp5_ASAP7_75t_L g1995 ( 
.A1(n_1942),
.A2(n_1938),
.B1(n_1940),
.B2(n_1799),
.C(n_1914),
.Y(n_1995)
);

HB1xp67_ASAP7_75t_L g1996 ( 
.A(n_1840),
.Y(n_1996)
);

BUFx3_ASAP7_75t_L g1997 ( 
.A(n_1874),
.Y(n_1997)
);

INVxp67_ASAP7_75t_L g1998 ( 
.A(n_1904),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1844),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1918),
.B(n_1935),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1936),
.B(n_1944),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1950),
.B(n_1832),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1928),
.B(n_1846),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1928),
.B(n_1823),
.Y(n_2004)
);

OR2x2_ASAP7_75t_L g2005 ( 
.A(n_1889),
.B(n_1827),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1928),
.B(n_1823),
.Y(n_2006)
);

AOI221xp5_ASAP7_75t_L g2007 ( 
.A1(n_1914),
.A2(n_1916),
.B1(n_1802),
.B2(n_1817),
.C(n_1922),
.Y(n_2007)
);

BUFx2_ASAP7_75t_L g2008 ( 
.A(n_1790),
.Y(n_2008)
);

INVxp67_ASAP7_75t_L g2009 ( 
.A(n_1919),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1928),
.B(n_1791),
.Y(n_2010)
);

HB1xp67_ASAP7_75t_L g2011 ( 
.A(n_1946),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1791),
.B(n_1813),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1941),
.B(n_1834),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1853),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1836),
.Y(n_2015)
);

HB1xp67_ASAP7_75t_L g2016 ( 
.A(n_1848),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1816),
.B(n_1837),
.Y(n_2017)
);

OAI211xp5_ASAP7_75t_L g2018 ( 
.A1(n_1949),
.A2(n_1941),
.B(n_1833),
.C(n_1913),
.Y(n_2018)
);

INVxp67_ASAP7_75t_SL g2019 ( 
.A(n_1868),
.Y(n_2019)
);

OR2x2_ASAP7_75t_SL g2020 ( 
.A(n_1905),
.B(n_1788),
.Y(n_2020)
);

AOI221xp5_ASAP7_75t_L g2021 ( 
.A1(n_1929),
.A2(n_1955),
.B1(n_1951),
.B2(n_1939),
.C(n_1849),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1871),
.B(n_1795),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1800),
.B(n_1797),
.Y(n_2023)
);

BUFx2_ASAP7_75t_L g2024 ( 
.A(n_1851),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1842),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1797),
.B(n_1787),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1888),
.B(n_1841),
.Y(n_2027)
);

HB1xp67_ASAP7_75t_L g2028 ( 
.A(n_1812),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1888),
.B(n_1898),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1911),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1867),
.B(n_1824),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1867),
.B(n_1808),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1911),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1834),
.B(n_1872),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1809),
.B(n_1899),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1854),
.B(n_1807),
.Y(n_2036)
);

AOI22xp33_ASAP7_75t_L g2037 ( 
.A1(n_1875),
.A2(n_1798),
.B1(n_1881),
.B2(n_1856),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1902),
.B(n_1878),
.Y(n_2038)
);

INVxp67_ASAP7_75t_SL g2039 ( 
.A(n_1878),
.Y(n_2039)
);

OR2x2_ASAP7_75t_L g2040 ( 
.A(n_1877),
.B(n_1920),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1794),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1892),
.B(n_1873),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1845),
.B(n_1927),
.Y(n_2043)
);

OR2x2_ASAP7_75t_L g2044 ( 
.A(n_1934),
.B(n_1957),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1908),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1907),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1907),
.Y(n_2047)
);

INVxp67_ASAP7_75t_SL g2048 ( 
.A(n_1882),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1818),
.B(n_1875),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1895),
.Y(n_2050)
);

BUFx3_ASAP7_75t_L g2051 ( 
.A(n_1874),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1912),
.B(n_1861),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1900),
.Y(n_2053)
);

AOI222xp33_ASAP7_75t_SL g2054 ( 
.A1(n_1947),
.A2(n_1876),
.B1(n_1879),
.B2(n_1958),
.C1(n_1811),
.C2(n_1865),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1793),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_1861),
.B(n_1804),
.Y(n_2056)
);

INVx3_ASAP7_75t_L g2057 ( 
.A(n_1930),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1789),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1910),
.Y(n_2059)
);

HB1xp67_ASAP7_75t_L g2060 ( 
.A(n_1822),
.Y(n_2060)
);

INVx3_ASAP7_75t_L g2061 ( 
.A(n_1930),
.Y(n_2061)
);

OAI221xp5_ASAP7_75t_L g2062 ( 
.A1(n_1925),
.A2(n_1883),
.B1(n_1798),
.B2(n_1866),
.C(n_1884),
.Y(n_2062)
);

BUFx2_ASAP7_75t_L g2063 ( 
.A(n_1981),
.Y(n_2063)
);

AOI22xp33_ASAP7_75t_L g2064 ( 
.A1(n_2049),
.A2(n_1873),
.B1(n_1906),
.B2(n_1856),
.Y(n_2064)
);

NAND3xp33_ASAP7_75t_L g2065 ( 
.A(n_2007),
.B(n_1885),
.C(n_1869),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2048),
.B(n_2056),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1996),
.Y(n_2067)
);

NAND4xp25_ASAP7_75t_L g2068 ( 
.A(n_2021),
.B(n_1884),
.C(n_1887),
.D(n_1814),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1973),
.Y(n_2069)
);

OAI211xp5_ASAP7_75t_L g2070 ( 
.A1(n_2018),
.A2(n_1865),
.B(n_1860),
.C(n_1897),
.Y(n_2070)
);

HB1xp67_ASAP7_75t_L g2071 ( 
.A(n_1981),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1996),
.Y(n_2072)
);

OAI33xp33_ASAP7_75t_L g2073 ( 
.A1(n_2042),
.A2(n_1869),
.A3(n_1855),
.B1(n_1858),
.B2(n_1901),
.B3(n_1893),
.Y(n_2073)
);

INVxp67_ASAP7_75t_SL g2074 ( 
.A(n_1963),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_2052),
.B(n_1862),
.Y(n_2075)
);

NOR2xp33_ASAP7_75t_SL g2076 ( 
.A(n_2062),
.B(n_1909),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2008),
.B(n_1926),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_2008),
.B(n_1897),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1990),
.Y(n_2079)
);

NAND2xp33_ASAP7_75t_SL g2080 ( 
.A(n_2013),
.B(n_1796),
.Y(n_2080)
);

AOI22xp33_ASAP7_75t_L g2081 ( 
.A1(n_2049),
.A2(n_1855),
.B1(n_1858),
.B2(n_1896),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_2035),
.B(n_1826),
.Y(n_2082)
);

INVxp67_ASAP7_75t_L g2083 ( 
.A(n_2056),
.Y(n_2083)
);

AOI221xp5_ASAP7_75t_L g2084 ( 
.A1(n_2007),
.A2(n_1995),
.B1(n_1980),
.B2(n_1979),
.C(n_1971),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_2035),
.B(n_1894),
.Y(n_2085)
);

OAI221xp5_ASAP7_75t_L g2086 ( 
.A1(n_1980),
.A2(n_1886),
.B1(n_1903),
.B2(n_1806),
.C(n_1852),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2035),
.B(n_1810),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_1965),
.B(n_1930),
.Y(n_2088)
);

NOR2xp33_ASAP7_75t_R g2089 ( 
.A(n_2057),
.B(n_1933),
.Y(n_2089)
);

INVxp67_ASAP7_75t_L g2090 ( 
.A(n_2056),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1990),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_1965),
.B(n_1828),
.Y(n_2092)
);

NAND2xp33_ASAP7_75t_R g2093 ( 
.A(n_2052),
.B(n_1917),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1990),
.Y(n_2094)
);

OR2x2_ASAP7_75t_L g2095 ( 
.A(n_1966),
.B(n_1828),
.Y(n_2095)
);

AOI322xp5_ASAP7_75t_L g2096 ( 
.A1(n_2042),
.A2(n_1847),
.A3(n_2034),
.B1(n_2037),
.B2(n_2031),
.C1(n_2049),
.C2(n_2013),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_1965),
.B(n_1989),
.Y(n_2097)
);

AOI221xp5_ASAP7_75t_L g2098 ( 
.A1(n_1995),
.A2(n_2062),
.B1(n_2036),
.B2(n_2028),
.C(n_2034),
.Y(n_2098)
);

BUFx2_ASAP7_75t_L g2099 ( 
.A(n_1986),
.Y(n_2099)
);

AOI22xp33_ASAP7_75t_SL g2100 ( 
.A1(n_2034),
.A2(n_2031),
.B1(n_2022),
.B2(n_2026),
.Y(n_2100)
);

AOI21x1_ASAP7_75t_L g2101 ( 
.A1(n_2016),
.A2(n_1963),
.B(n_2060),
.Y(n_2101)
);

OAI321xp33_ASAP7_75t_L g2102 ( 
.A1(n_2018),
.A2(n_2021),
.A3(n_2031),
.B1(n_2036),
.B2(n_2048),
.C(n_2022),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_1989),
.B(n_2017),
.Y(n_2103)
);

OR2x2_ASAP7_75t_L g2104 ( 
.A(n_1966),
.B(n_2014),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_1989),
.B(n_2017),
.Y(n_2105)
);

AOI22xp33_ASAP7_75t_L g2106 ( 
.A1(n_2022),
.A2(n_2026),
.B1(n_2047),
.B2(n_2046),
.Y(n_2106)
);

AOI222xp33_ASAP7_75t_L g2107 ( 
.A1(n_2052),
.A2(n_2026),
.B1(n_2023),
.B2(n_2029),
.C1(n_2032),
.C2(n_2047),
.Y(n_2107)
);

AOI222xp33_ASAP7_75t_L g2108 ( 
.A1(n_2023),
.A2(n_2046),
.B1(n_2010),
.B2(n_2036),
.C1(n_2028),
.C2(n_2027),
.Y(n_2108)
);

OAI33xp33_ASAP7_75t_L g2109 ( 
.A1(n_1962),
.A2(n_1978),
.A3(n_2038),
.B1(n_2014),
.B2(n_2001),
.B3(n_2000),
.Y(n_2109)
);

BUFx2_ASAP7_75t_L g2110 ( 
.A(n_1986),
.Y(n_2110)
);

OAI31xp33_ASAP7_75t_L g2111 ( 
.A1(n_2029),
.A2(n_2038),
.A3(n_2023),
.B(n_2041),
.Y(n_2111)
);

AOI22xp33_ASAP7_75t_L g2112 ( 
.A1(n_2045),
.A2(n_2027),
.B1(n_2041),
.B2(n_2055),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2017),
.B(n_1964),
.Y(n_2113)
);

OR2x2_ASAP7_75t_L g2114 ( 
.A(n_1978),
.B(n_1975),
.Y(n_2114)
);

INVx4_ASAP7_75t_L g2115 ( 
.A(n_2057),
.Y(n_2115)
);

OAI31xp33_ASAP7_75t_SL g2116 ( 
.A1(n_2039),
.A2(n_2029),
.A3(n_1994),
.B(n_2002),
.Y(n_2116)
);

BUFx6f_ASAP7_75t_L g2117 ( 
.A(n_1992),
.Y(n_2117)
);

AND2x4_ASAP7_75t_L g2118 ( 
.A(n_1985),
.B(n_1972),
.Y(n_2118)
);

OR2x2_ASAP7_75t_L g2119 ( 
.A(n_1975),
.B(n_2003),
.Y(n_2119)
);

AOI211xp5_ASAP7_75t_SL g2120 ( 
.A1(n_2060),
.A2(n_2016),
.B(n_2010),
.C(n_2039),
.Y(n_2120)
);

INVx3_ASAP7_75t_L g2121 ( 
.A(n_2015),
.Y(n_2121)
);

AOI22xp33_ASAP7_75t_L g2122 ( 
.A1(n_2045),
.A2(n_2027),
.B1(n_2041),
.B2(n_2055),
.Y(n_2122)
);

NOR2xp33_ASAP7_75t_R g2123 ( 
.A(n_2057),
.B(n_2061),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1991),
.Y(n_2124)
);

INVx1_ASAP7_75t_SL g2125 ( 
.A(n_2024),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_1964),
.B(n_2003),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1991),
.Y(n_2127)
);

AOI22xp33_ASAP7_75t_L g2128 ( 
.A1(n_2055),
.A2(n_2058),
.B1(n_2010),
.B2(n_2012),
.Y(n_2128)
);

INVx2_ASAP7_75t_SL g2129 ( 
.A(n_1997),
.Y(n_2129)
);

OAI31xp33_ASAP7_75t_L g2130 ( 
.A1(n_2058),
.A2(n_2054),
.A3(n_2032),
.B(n_2002),
.Y(n_2130)
);

NOR2xp33_ASAP7_75t_R g2131 ( 
.A(n_2057),
.B(n_2061),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_1964),
.B(n_2003),
.Y(n_2132)
);

OAI31xp33_ASAP7_75t_SL g2133 ( 
.A1(n_2002),
.A2(n_2043),
.A3(n_2032),
.B(n_2054),
.Y(n_2133)
);

OAI221xp5_ASAP7_75t_L g2134 ( 
.A1(n_2058),
.A2(n_2059),
.B1(n_2025),
.B2(n_2004),
.C(n_2006),
.Y(n_2134)
);

INVx2_ASAP7_75t_SL g2135 ( 
.A(n_1997),
.Y(n_2135)
);

OR2x2_ASAP7_75t_L g2136 ( 
.A(n_1998),
.B(n_2005),
.Y(n_2136)
);

OR2x2_ASAP7_75t_L g2137 ( 
.A(n_1998),
.B(n_2005),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1991),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2103),
.B(n_2043),
.Y(n_2139)
);

NOR2xp67_ASAP7_75t_L g2140 ( 
.A(n_2083),
.B(n_2059),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_2121),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_2066),
.B(n_2133),
.Y(n_2142)
);

OR2x2_ASAP7_75t_L g2143 ( 
.A(n_2119),
.B(n_2040),
.Y(n_2143)
);

INVx1_ASAP7_75t_SL g2144 ( 
.A(n_2089),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2103),
.B(n_2043),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2067),
.Y(n_2146)
);

OR2x2_ASAP7_75t_L g2147 ( 
.A(n_2119),
.B(n_2040),
.Y(n_2147)
);

OR2x2_ASAP7_75t_L g2148 ( 
.A(n_2114),
.B(n_1960),
.Y(n_2148)
);

OR2x2_ASAP7_75t_L g2149 ( 
.A(n_2114),
.B(n_1960),
.Y(n_2149)
);

INVx1_ASAP7_75t_SL g2150 ( 
.A(n_2077),
.Y(n_2150)
);

BUFx2_ASAP7_75t_L g2151 ( 
.A(n_2063),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2105),
.B(n_2044),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2133),
.B(n_1962),
.Y(n_2153)
);

INVx6_ASAP7_75t_L g2154 ( 
.A(n_2115),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2067),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_2121),
.Y(n_2156)
);

OR2x6_ASAP7_75t_L g2157 ( 
.A(n_2077),
.B(n_2004),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2090),
.B(n_2050),
.Y(n_2158)
);

NOR2x1_ASAP7_75t_L g2159 ( 
.A(n_2099),
.B(n_1992),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_2116),
.B(n_2050),
.Y(n_2160)
);

OR2x2_ASAP7_75t_L g2161 ( 
.A(n_2104),
.B(n_2044),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_2105),
.B(n_2025),
.Y(n_2162)
);

AOI22xp33_ASAP7_75t_SL g2163 ( 
.A1(n_2076),
.A2(n_2065),
.B1(n_2078),
.B2(n_2087),
.Y(n_2163)
);

AND2x4_ASAP7_75t_L g2164 ( 
.A(n_2118),
.B(n_1984),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2072),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_2097),
.B(n_2025),
.Y(n_2166)
);

INVx4_ASAP7_75t_L g2167 ( 
.A(n_2115),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2072),
.Y(n_2168)
);

NOR2xp67_ASAP7_75t_L g2169 ( 
.A(n_2101),
.B(n_2059),
.Y(n_2169)
);

INVx4_ASAP7_75t_L g2170 ( 
.A(n_2115),
.Y(n_2170)
);

HB1xp67_ASAP7_75t_L g2171 ( 
.A(n_2071),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2116),
.B(n_2053),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2097),
.B(n_1982),
.Y(n_2173)
);

INVx1_ASAP7_75t_SL g2174 ( 
.A(n_2136),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_2113),
.B(n_1982),
.Y(n_2175)
);

OAI21xp5_ASAP7_75t_L g2176 ( 
.A1(n_2102),
.A2(n_2006),
.B(n_2004),
.Y(n_2176)
);

NOR2xp33_ASAP7_75t_L g2177 ( 
.A(n_2102),
.B(n_1997),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_2113),
.B(n_1982),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2104),
.B(n_2053),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_2121),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_2107),
.B(n_1967),
.Y(n_2181)
);

HB1xp67_ASAP7_75t_L g2182 ( 
.A(n_2063),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2079),
.Y(n_2183)
);

HB1xp67_ASAP7_75t_L g2184 ( 
.A(n_2099),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2107),
.B(n_1967),
.Y(n_2185)
);

NOR2xp33_ASAP7_75t_L g2186 ( 
.A(n_2068),
.B(n_2051),
.Y(n_2186)
);

OR2x2_ASAP7_75t_L g2187 ( 
.A(n_2136),
.B(n_1967),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2137),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2137),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2079),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2126),
.B(n_1977),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_2126),
.B(n_1977),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2091),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_2121),
.Y(n_2194)
);

INVx4_ASAP7_75t_L g2195 ( 
.A(n_2115),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2111),
.B(n_1993),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2091),
.Y(n_2197)
);

OR2x2_ASAP7_75t_L g2198 ( 
.A(n_2132),
.B(n_2000),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2094),
.Y(n_2199)
);

INVxp67_ASAP7_75t_SL g2200 ( 
.A(n_2101),
.Y(n_2200)
);

INVx2_ASAP7_75t_SL g2201 ( 
.A(n_2118),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_2111),
.B(n_2078),
.Y(n_2202)
);

AND2x4_ASAP7_75t_SL g2203 ( 
.A(n_2088),
.B(n_1984),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2094),
.Y(n_2204)
);

OR2x6_ASAP7_75t_L g2205 ( 
.A(n_2117),
.B(n_2006),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2124),
.Y(n_2206)
);

NAND2x1_ASAP7_75t_L g2207 ( 
.A(n_2118),
.B(n_1984),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_2069),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2146),
.Y(n_2209)
);

HB1xp67_ASAP7_75t_L g2210 ( 
.A(n_2171),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2161),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2153),
.B(n_2110),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2161),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2188),
.Y(n_2214)
);

AND2x4_ASAP7_75t_L g2215 ( 
.A(n_2157),
.B(n_2118),
.Y(n_2215)
);

INVxp67_ASAP7_75t_SL g2216 ( 
.A(n_2169),
.Y(n_2216)
);

INVxp67_ASAP7_75t_L g2217 ( 
.A(n_2177),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2142),
.B(n_2110),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2160),
.B(n_2130),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_2172),
.B(n_2130),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2155),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2165),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2168),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2183),
.Y(n_2224)
);

HB1xp67_ASAP7_75t_L g2225 ( 
.A(n_2182),
.Y(n_2225)
);

NAND2x1_ASAP7_75t_L g2226 ( 
.A(n_2159),
.B(n_2132),
.Y(n_2226)
);

BUFx2_ASAP7_75t_L g2227 ( 
.A(n_2157),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2183),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2193),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2191),
.B(n_2082),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_2208),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_2191),
.B(n_2082),
.Y(n_2232)
);

BUFx3_ASAP7_75t_L g2233 ( 
.A(n_2144),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2179),
.B(n_2100),
.Y(n_2234)
);

HB1xp67_ASAP7_75t_L g2235 ( 
.A(n_2184),
.Y(n_2235)
);

OR2x2_ASAP7_75t_L g2236 ( 
.A(n_2148),
.B(n_2149),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2189),
.Y(n_2237)
);

OR2x2_ASAP7_75t_L g2238 ( 
.A(n_2148),
.B(n_2149),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2143),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2196),
.B(n_2098),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2143),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2147),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2174),
.B(n_2158),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2166),
.B(n_2108),
.Y(n_2244)
);

OR2x2_ASAP7_75t_L g2245 ( 
.A(n_2187),
.B(n_2124),
.Y(n_2245)
);

NAND2x1p5_ASAP7_75t_L g2246 ( 
.A(n_2207),
.B(n_1992),
.Y(n_2246)
);

OR2x2_ASAP7_75t_L g2247 ( 
.A(n_2187),
.B(n_2127),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2147),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_2192),
.B(n_2127),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2198),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2198),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2166),
.B(n_2092),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_2192),
.B(n_2138),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_SL g2254 ( 
.A(n_2186),
.B(n_2065),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2193),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2197),
.Y(n_2256)
);

INVx2_ASAP7_75t_SL g2257 ( 
.A(n_2203),
.Y(n_2257)
);

OAI21xp33_ASAP7_75t_SL g2258 ( 
.A1(n_2150),
.A2(n_2075),
.B(n_2125),
.Y(n_2258)
);

NOR2xp33_ASAP7_75t_SL g2259 ( 
.A(n_2176),
.B(n_2076),
.Y(n_2259)
);

AND2x2_ASAP7_75t_L g2260 ( 
.A(n_2139),
.B(n_2138),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2190),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_2215),
.B(n_2164),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2215),
.B(n_2164),
.Y(n_2263)
);

INVx1_ASAP7_75t_SL g2264 ( 
.A(n_2233),
.Y(n_2264)
);

OR2x2_ASAP7_75t_L g2265 ( 
.A(n_2236),
.B(n_2181),
.Y(n_2265)
);

NOR2x1_ASAP7_75t_R g2266 ( 
.A(n_2233),
.B(n_2093),
.Y(n_2266)
);

NAND2xp33_ASAP7_75t_SL g2267 ( 
.A(n_2226),
.B(n_2212),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2209),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2219),
.B(n_2202),
.Y(n_2269)
);

OR2x2_ASAP7_75t_L g2270 ( 
.A(n_2236),
.B(n_2185),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2220),
.B(n_2162),
.Y(n_2271)
);

AND2x4_ASAP7_75t_SL g2272 ( 
.A(n_2215),
.B(n_2164),
.Y(n_2272)
);

HB1xp67_ASAP7_75t_L g2273 ( 
.A(n_2210),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2218),
.B(n_2162),
.Y(n_2274)
);

INVx1_ASAP7_75t_SL g2275 ( 
.A(n_2254),
.Y(n_2275)
);

AOI32xp33_ASAP7_75t_L g2276 ( 
.A1(n_2259),
.A2(n_2163),
.A3(n_2120),
.B1(n_2106),
.B2(n_2080),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2209),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_2231),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2221),
.Y(n_2279)
);

OR2x2_ASAP7_75t_L g2280 ( 
.A(n_2238),
.B(n_2151),
.Y(n_2280)
);

AND2x2_ASAP7_75t_L g2281 ( 
.A(n_2227),
.B(n_2139),
.Y(n_2281)
);

HB1xp67_ASAP7_75t_L g2282 ( 
.A(n_2235),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2234),
.B(n_2151),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2221),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_2227),
.B(n_2145),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_SL g2286 ( 
.A(n_2258),
.B(n_2167),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2222),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_2231),
.Y(n_2288)
);

INVx1_ASAP7_75t_SL g2289 ( 
.A(n_2238),
.Y(n_2289)
);

INVx1_ASAP7_75t_SL g2290 ( 
.A(n_2240),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2222),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2243),
.B(n_2145),
.Y(n_2292)
);

OR2x6_ASAP7_75t_L g2293 ( 
.A(n_2217),
.B(n_2205),
.Y(n_2293)
);

BUFx3_ASAP7_75t_L g2294 ( 
.A(n_2225),
.Y(n_2294)
);

INVx1_ASAP7_75t_SL g2295 ( 
.A(n_2244),
.Y(n_2295)
);

NOR2xp33_ASAP7_75t_L g2296 ( 
.A(n_2252),
.B(n_2109),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2211),
.B(n_2152),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2223),
.Y(n_2298)
);

HB1xp67_ASAP7_75t_L g2299 ( 
.A(n_2223),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2213),
.B(n_2152),
.Y(n_2300)
);

AND2x4_ASAP7_75t_L g2301 ( 
.A(n_2257),
.B(n_2157),
.Y(n_2301)
);

OR2x2_ASAP7_75t_L g2302 ( 
.A(n_2239),
.B(n_2197),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2214),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2237),
.B(n_2096),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2261),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2224),
.Y(n_2306)
);

OR2x2_ASAP7_75t_L g2307 ( 
.A(n_2241),
.B(n_2095),
.Y(n_2307)
);

INVx2_ASAP7_75t_SL g2308 ( 
.A(n_2257),
.Y(n_2308)
);

OAI31xp33_ASAP7_75t_L g2309 ( 
.A1(n_2216),
.A2(n_2070),
.A3(n_2134),
.B(n_2087),
.Y(n_2309)
);

AND2x4_ASAP7_75t_L g2310 ( 
.A(n_2242),
.B(n_2157),
.Y(n_2310)
);

NAND2xp33_ASAP7_75t_SL g2311 ( 
.A(n_2226),
.B(n_2207),
.Y(n_2311)
);

OR2x2_ASAP7_75t_L g2312 ( 
.A(n_2248),
.B(n_2206),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_2296),
.B(n_2250),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2299),
.Y(n_2314)
);

NOR2xp67_ASAP7_75t_L g2315 ( 
.A(n_2286),
.B(n_2201),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2306),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2296),
.B(n_2251),
.Y(n_2317)
);

NOR2x1_ASAP7_75t_L g2318 ( 
.A(n_2264),
.B(n_2068),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2268),
.Y(n_2319)
);

AOI32xp33_ASAP7_75t_L g2320 ( 
.A1(n_2275),
.A2(n_2200),
.A3(n_2084),
.B1(n_2122),
.B2(n_2112),
.Y(n_2320)
);

AOI311xp33_ASAP7_75t_L g2321 ( 
.A1(n_2305),
.A2(n_2283),
.A3(n_2279),
.B(n_2277),
.C(n_2284),
.Y(n_2321)
);

AOI21xp5_ASAP7_75t_L g2322 ( 
.A1(n_2276),
.A2(n_2073),
.B(n_2081),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2287),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2271),
.B(n_2096),
.Y(n_2324)
);

INVx2_ASAP7_75t_SL g2325 ( 
.A(n_2301),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2291),
.Y(n_2326)
);

NOR2xp33_ASAP7_75t_SL g2327 ( 
.A(n_2266),
.B(n_2167),
.Y(n_2327)
);

OR2x2_ASAP7_75t_L g2328 ( 
.A(n_2270),
.B(n_2245),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2298),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2303),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_2281),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2273),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2282),
.Y(n_2333)
);

AOI21xp33_ASAP7_75t_SL g2334 ( 
.A1(n_2286),
.A2(n_2246),
.B(n_2201),
.Y(n_2334)
);

AOI21xp33_ASAP7_75t_L g2335 ( 
.A1(n_2290),
.A2(n_2095),
.B(n_2064),
.Y(n_2335)
);

OAI21xp5_ASAP7_75t_SL g2336 ( 
.A1(n_2289),
.A2(n_2246),
.B(n_2086),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_2281),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2269),
.B(n_2230),
.Y(n_2338)
);

O2A1O1Ixp33_ASAP7_75t_L g2339 ( 
.A1(n_2304),
.A2(n_2092),
.B(n_2074),
.C(n_2128),
.Y(n_2339)
);

AOI21xp33_ASAP7_75t_SL g2340 ( 
.A1(n_2308),
.A2(n_2246),
.B(n_2247),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2294),
.B(n_2230),
.Y(n_2341)
);

A2O1A1Ixp33_ASAP7_75t_L g2342 ( 
.A1(n_2309),
.A2(n_2140),
.B(n_2085),
.C(n_1987),
.Y(n_2342)
);

OAI21xp5_ASAP7_75t_SL g2343 ( 
.A1(n_2301),
.A2(n_2203),
.B(n_2088),
.Y(n_2343)
);

AOI21xp33_ASAP7_75t_L g2344 ( 
.A1(n_2295),
.A2(n_2019),
.B(n_2224),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2302),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2302),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2294),
.B(n_2232),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2274),
.B(n_2232),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2312),
.Y(n_2349)
);

INVxp67_ASAP7_75t_L g2350 ( 
.A(n_2308),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2272),
.B(n_2260),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2312),
.Y(n_2352)
);

OAI21xp5_ASAP7_75t_L g2353 ( 
.A1(n_2267),
.A2(n_2228),
.B(n_2255),
.Y(n_2353)
);

INVxp67_ASAP7_75t_L g2354 ( 
.A(n_2318),
.Y(n_2354)
);

OAI221xp5_ASAP7_75t_L g2355 ( 
.A1(n_2342),
.A2(n_2267),
.B1(n_2270),
.B2(n_2265),
.C(n_2293),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2316),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2338),
.B(n_2285),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2316),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2319),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2322),
.B(n_2285),
.Y(n_2360)
);

NOR2x1p5_ASAP7_75t_L g2361 ( 
.A(n_2341),
.B(n_2280),
.Y(n_2361)
);

AOI221xp5_ASAP7_75t_L g2362 ( 
.A1(n_2313),
.A2(n_2307),
.B1(n_2288),
.B2(n_2278),
.C(n_2311),
.Y(n_2362)
);

OAI22xp5_ASAP7_75t_L g2363 ( 
.A1(n_2342),
.A2(n_2301),
.B1(n_2272),
.B2(n_2293),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2319),
.Y(n_2364)
);

INVxp67_ASAP7_75t_L g2365 ( 
.A(n_2325),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2346),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2331),
.B(n_2280),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2346),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2323),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2326),
.Y(n_2370)
);

NOR2xp33_ASAP7_75t_L g2371 ( 
.A(n_2325),
.B(n_2310),
.Y(n_2371)
);

OAI21xp5_ASAP7_75t_L g2372 ( 
.A1(n_2353),
.A2(n_2293),
.B(n_2310),
.Y(n_2372)
);

AOI221xp5_ASAP7_75t_L g2373 ( 
.A1(n_2317),
.A2(n_2278),
.B1(n_2288),
.B2(n_2311),
.C(n_2310),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2331),
.B(n_2292),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2329),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_2351),
.B(n_2262),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2345),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_2337),
.B(n_2297),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2337),
.B(n_2300),
.Y(n_2379)
);

AOI21xp5_ASAP7_75t_L g2380 ( 
.A1(n_2324),
.A2(n_2336),
.B(n_2339),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2349),
.Y(n_2381)
);

AOI321xp33_ASAP7_75t_L g2382 ( 
.A1(n_2321),
.A2(n_2335),
.A3(n_2344),
.B1(n_2352),
.B2(n_2334),
.C(n_2347),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2330),
.Y(n_2383)
);

OAI221xp5_ASAP7_75t_L g2384 ( 
.A1(n_2320),
.A2(n_2293),
.B1(n_2205),
.B2(n_1987),
.C(n_1988),
.Y(n_2384)
);

INVxp67_ASAP7_75t_L g2385 ( 
.A(n_2371),
.Y(n_2385)
);

AOI21xp5_ASAP7_75t_L g2386 ( 
.A1(n_2354),
.A2(n_2327),
.B(n_2315),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2356),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_SL g2388 ( 
.A(n_2382),
.B(n_2350),
.Y(n_2388)
);

NAND3xp33_ASAP7_75t_L g2389 ( 
.A(n_2380),
.B(n_2332),
.C(n_2333),
.Y(n_2389)
);

AND2x2_ASAP7_75t_L g2390 ( 
.A(n_2376),
.B(n_2351),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2360),
.B(n_2314),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2361),
.Y(n_2392)
);

INVx2_ASAP7_75t_SL g2393 ( 
.A(n_2376),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2365),
.B(n_2328),
.Y(n_2394)
);

NAND3xp33_ASAP7_75t_L g2395 ( 
.A(n_2362),
.B(n_2340),
.C(n_2328),
.Y(n_2395)
);

NOR2x1_ASAP7_75t_L g2396 ( 
.A(n_2356),
.B(n_2358),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_2358),
.Y(n_2397)
);

BUFx3_ASAP7_75t_L g2398 ( 
.A(n_2377),
.Y(n_2398)
);

INVxp67_ASAP7_75t_L g2399 ( 
.A(n_2371),
.Y(n_2399)
);

NOR2xp33_ASAP7_75t_L g2400 ( 
.A(n_2377),
.B(n_2343),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2359),
.Y(n_2401)
);

INVxp67_ASAP7_75t_SL g2402 ( 
.A(n_2367),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2357),
.B(n_2348),
.Y(n_2403)
);

NOR2xp33_ASAP7_75t_L g2404 ( 
.A(n_2383),
.B(n_2262),
.Y(n_2404)
);

CKINVDCx20_ASAP7_75t_R g2405 ( 
.A(n_2381),
.Y(n_2405)
);

NAND3xp33_ASAP7_75t_L g2406 ( 
.A(n_2373),
.B(n_2256),
.C(n_2255),
.Y(n_2406)
);

AOI22xp5_ASAP7_75t_L g2407 ( 
.A1(n_2355),
.A2(n_2085),
.B1(n_1987),
.B2(n_1988),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2364),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2366),
.Y(n_2409)
);

OAI21xp33_ASAP7_75t_SL g2410 ( 
.A1(n_2388),
.A2(n_2372),
.B(n_2368),
.Y(n_2410)
);

NOR4xp25_ASAP7_75t_L g2411 ( 
.A(n_2388),
.B(n_2369),
.C(n_2370),
.D(n_2375),
.Y(n_2411)
);

AOI31xp33_ASAP7_75t_L g2412 ( 
.A1(n_2385),
.A2(n_2379),
.A3(n_2378),
.B(n_2374),
.Y(n_2412)
);

NOR2xp67_ASAP7_75t_L g2413 ( 
.A(n_2393),
.B(n_2363),
.Y(n_2413)
);

NOR2xp33_ASAP7_75t_SL g2414 ( 
.A(n_2399),
.B(n_2384),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_2390),
.Y(n_2415)
);

OAI211xp5_ASAP7_75t_SL g2416 ( 
.A1(n_2391),
.A2(n_2247),
.B(n_2245),
.C(n_2229),
.Y(n_2416)
);

AOI22xp5_ASAP7_75t_L g2417 ( 
.A1(n_2405),
.A2(n_2205),
.B1(n_1988),
.B2(n_2263),
.Y(n_2417)
);

NOR3xp33_ASAP7_75t_L g2418 ( 
.A(n_2389),
.B(n_2263),
.C(n_2001),
.Y(n_2418)
);

NAND3xp33_ASAP7_75t_SL g2419 ( 
.A(n_2386),
.B(n_2123),
.C(n_2131),
.Y(n_2419)
);

NAND4xp25_ASAP7_75t_L g2420 ( 
.A(n_2400),
.B(n_2167),
.C(n_2195),
.D(n_2170),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2402),
.B(n_2228),
.Y(n_2421)
);

INVxp67_ASAP7_75t_L g2422 ( 
.A(n_2394),
.Y(n_2422)
);

NAND4xp25_ASAP7_75t_L g2423 ( 
.A(n_2400),
.B(n_2195),
.C(n_2170),
.D(n_2061),
.Y(n_2423)
);

NOR2xp33_ASAP7_75t_L g2424 ( 
.A(n_2405),
.B(n_2229),
.Y(n_2424)
);

OAI21xp33_ASAP7_75t_L g2425 ( 
.A1(n_2414),
.A2(n_2404),
.B(n_2407),
.Y(n_2425)
);

AOI221xp5_ASAP7_75t_SL g2426 ( 
.A1(n_2410),
.A2(n_2392),
.B1(n_2404),
.B2(n_2409),
.C(n_2408),
.Y(n_2426)
);

NAND4xp25_ASAP7_75t_SL g2427 ( 
.A(n_2415),
.B(n_2395),
.C(n_2396),
.D(n_2403),
.Y(n_2427)
);

NAND3xp33_ASAP7_75t_SL g2428 ( 
.A(n_2411),
.B(n_2392),
.C(n_2397),
.Y(n_2428)
);

AOI221xp5_ASAP7_75t_L g2429 ( 
.A1(n_2412),
.A2(n_2398),
.B1(n_2397),
.B2(n_2387),
.C(n_2401),
.Y(n_2429)
);

AOI211xp5_ASAP7_75t_L g2430 ( 
.A1(n_2413),
.A2(n_2398),
.B(n_2406),
.C(n_2117),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2421),
.Y(n_2431)
);

AOI221xp5_ASAP7_75t_L g2432 ( 
.A1(n_2422),
.A2(n_2424),
.B1(n_2416),
.B2(n_2418),
.C(n_2417),
.Y(n_2432)
);

AOI221x1_ASAP7_75t_L g2433 ( 
.A1(n_2420),
.A2(n_2256),
.B1(n_2195),
.B2(n_2170),
.C(n_2194),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2423),
.Y(n_2434)
);

AO21x1_ASAP7_75t_L g2435 ( 
.A1(n_2419),
.A2(n_2260),
.B(n_2249),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2411),
.B(n_2249),
.Y(n_2436)
);

AOI322xp5_ASAP7_75t_L g2437 ( 
.A1(n_2410),
.A2(n_2012),
.A3(n_1977),
.B1(n_1970),
.B2(n_1983),
.C1(n_2030),
.C2(n_2033),
.Y(n_2437)
);

NOR2x1_ASAP7_75t_L g2438 ( 
.A(n_2428),
.B(n_2061),
.Y(n_2438)
);

NAND2xp33_ASAP7_75t_R g2439 ( 
.A(n_2431),
.B(n_2205),
.Y(n_2439)
);

NOR2xp33_ASAP7_75t_R g2440 ( 
.A(n_2427),
.B(n_2154),
.Y(n_2440)
);

INVx1_ASAP7_75t_SL g2441 ( 
.A(n_2436),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2429),
.Y(n_2442)
);

AOI21xp33_ASAP7_75t_SL g2443 ( 
.A1(n_2425),
.A2(n_2135),
.B(n_2129),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2426),
.B(n_2141),
.Y(n_2444)
);

NOR2xp33_ASAP7_75t_L g2445 ( 
.A(n_2443),
.B(n_2434),
.Y(n_2445)
);

AO22x1_ASAP7_75t_L g2446 ( 
.A1(n_2438),
.A2(n_2430),
.B1(n_2437),
.B2(n_2432),
.Y(n_2446)
);

AND3x4_ASAP7_75t_L g2447 ( 
.A(n_2440),
.B(n_2433),
.C(n_2435),
.Y(n_2447)
);

NOR4xp75_ASAP7_75t_SL g2448 ( 
.A(n_2444),
.B(n_2154),
.C(n_2020),
.D(n_2125),
.Y(n_2448)
);

INVx1_ASAP7_75t_SL g2449 ( 
.A(n_2441),
.Y(n_2449)
);

NOR2xp67_ASAP7_75t_L g2450 ( 
.A(n_2442),
.B(n_2253),
.Y(n_2450)
);

AND3x4_ASAP7_75t_L g2451 ( 
.A(n_2439),
.B(n_2051),
.C(n_2154),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_2438),
.B(n_2141),
.Y(n_2452)
);

NAND3xp33_ASAP7_75t_L g2453 ( 
.A(n_2445),
.B(n_2446),
.C(n_2450),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2449),
.B(n_2156),
.Y(n_2454)
);

AOI22xp5_ASAP7_75t_L g2455 ( 
.A1(n_2451),
.A2(n_2117),
.B1(n_2173),
.B2(n_2019),
.Y(n_2455)
);

AOI32xp33_ASAP7_75t_L g2456 ( 
.A1(n_2452),
.A2(n_2173),
.A3(n_2253),
.B1(n_2175),
.B2(n_2178),
.Y(n_2456)
);

NAND3xp33_ASAP7_75t_L g2457 ( 
.A(n_2448),
.B(n_2117),
.C(n_2180),
.Y(n_2457)
);

NOR4xp25_ASAP7_75t_L g2458 ( 
.A(n_2447),
.B(n_2178),
.C(n_2175),
.D(n_2206),
.Y(n_2458)
);

NOR4xp25_ASAP7_75t_L g2459 ( 
.A(n_2449),
.B(n_2199),
.C(n_2204),
.D(n_2194),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2454),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2453),
.Y(n_2461)
);

CKINVDCx5p33_ASAP7_75t_R g2462 ( 
.A(n_2455),
.Y(n_2462)
);

HB1xp67_ASAP7_75t_L g2463 ( 
.A(n_2458),
.Y(n_2463)
);

XNOR2xp5_ASAP7_75t_L g2464 ( 
.A(n_2461),
.B(n_2457),
.Y(n_2464)
);

XNOR2xp5_ASAP7_75t_L g2465 ( 
.A(n_2463),
.B(n_2462),
.Y(n_2465)
);

XNOR2x1_ASAP7_75t_L g2466 ( 
.A(n_2465),
.B(n_2460),
.Y(n_2466)
);

OAI22xp5_ASAP7_75t_L g2467 ( 
.A1(n_2464),
.A2(n_2460),
.B1(n_2456),
.B2(n_2459),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2466),
.Y(n_2468)
);

AOI22xp33_ASAP7_75t_SL g2469 ( 
.A1(n_2467),
.A2(n_2154),
.B1(n_2117),
.B2(n_2180),
.Y(n_2469)
);

CKINVDCx20_ASAP7_75t_R g2470 ( 
.A(n_2467),
.Y(n_2470)
);

AOI21xp5_ASAP7_75t_L g2471 ( 
.A1(n_2468),
.A2(n_2156),
.B(n_2135),
.Y(n_2471)
);

AOI21xp5_ASAP7_75t_L g2472 ( 
.A1(n_2469),
.A2(n_2129),
.B(n_1993),
.Y(n_2472)
);

OAI21xp5_ASAP7_75t_L g2473 ( 
.A1(n_2471),
.A2(n_2470),
.B(n_1999),
.Y(n_2473)
);

AOI22xp33_ASAP7_75t_SL g2474 ( 
.A1(n_2472),
.A2(n_2051),
.B1(n_1999),
.B2(n_2208),
.Y(n_2474)
);

NAND3xp33_ASAP7_75t_L g2475 ( 
.A(n_2473),
.B(n_2011),
.C(n_2009),
.Y(n_2475)
);

AOI22xp33_ASAP7_75t_L g2476 ( 
.A1(n_2475),
.A2(n_2474),
.B1(n_1974),
.B2(n_1976),
.Y(n_2476)
);

AOI211xp5_ASAP7_75t_L g2477 ( 
.A1(n_2476),
.A2(n_1961),
.B(n_1968),
.C(n_1969),
.Y(n_2477)
);


endmodule