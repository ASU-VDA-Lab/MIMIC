module fake_netlist_6_1622_n_903 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_903);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_903;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_893;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_758;
wire n_525;
wire n_720;
wire n_842;
wire n_611;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_184;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_438;
wire n_267;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_484;
wire n_262;
wire n_613;
wire n_736;
wire n_187;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_176),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_94),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_118),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_51),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_57),
.Y(n_188)
);

NOR2xp67_ASAP7_75t_L g189 ( 
.A(n_114),
.B(n_151),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_15),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_111),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_11),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_59),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_0),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_160),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_169),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_132),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_166),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_106),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_167),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_78),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_52),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_1),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_85),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_12),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_42),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_122),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_127),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_17),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_14),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_39),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_79),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_156),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_7),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_168),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_34),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_124),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_61),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_35),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_50),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_145),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_153),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_30),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_18),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_45),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g229 ( 
.A(n_107),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_89),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_26),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_1),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_110),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_149),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_98),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_55),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_141),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_101),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_178),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_143),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_64),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_100),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_10),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_11),
.B(n_134),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_32),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_135),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_76),
.Y(n_247)
);

BUFx2_ASAP7_75t_SL g248 ( 
.A(n_8),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_40),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_74),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_137),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_66),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_6),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_60),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_87),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_163),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_90),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_65),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_0),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_120),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_125),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_108),
.Y(n_262)
);

NOR2xp67_ASAP7_75t_L g263 ( 
.A(n_129),
.B(n_91),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_146),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_97),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_29),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_67),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_185),
.B(n_2),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_190),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_246),
.Y(n_270)
);

AND2x4_ASAP7_75t_L g271 ( 
.A(n_207),
.B(n_2),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_207),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_205),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_274)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_246),
.Y(n_275)
);

AND2x6_ASAP7_75t_L g276 ( 
.A(n_246),
.B(n_27),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_235),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_208),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_190),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_246),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_243),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_243),
.Y(n_282)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_229),
.Y(n_283)
);

BUFx8_ASAP7_75t_L g284 ( 
.A(n_223),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_243),
.Y(n_285)
);

BUFx8_ASAP7_75t_SL g286 ( 
.A(n_205),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_185),
.B(n_3),
.Y(n_287)
);

AOI22x1_ASAP7_75t_SL g288 ( 
.A1(n_192),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_227),
.Y(n_289)
);

BUFx12f_ASAP7_75t_L g290 ( 
.A(n_229),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_235),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_244),
.B(n_7),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_184),
.Y(n_293)
);

AND2x4_ASAP7_75t_L g294 ( 
.A(n_225),
.B(n_8),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_248),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_253),
.Y(n_296)
);

AND2x4_ASAP7_75t_L g297 ( 
.A(n_225),
.B(n_9),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_208),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_194),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_259),
.Y(n_300)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_229),
.Y(n_301)
);

AND2x2_ASAP7_75t_SL g302 ( 
.A(n_186),
.B(n_13),
.Y(n_302)
);

BUFx12f_ASAP7_75t_L g303 ( 
.A(n_240),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_195),
.Y(n_304)
);

AND2x4_ASAP7_75t_L g305 ( 
.A(n_187),
.B(n_13),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_188),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_191),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_202),
.B(n_211),
.Y(n_308)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_240),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_193),
.Y(n_310)
);

INVx6_ASAP7_75t_L g311 ( 
.A(n_240),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_200),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_203),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_206),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_214),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_216),
.Y(n_316)
);

OAI22x1_ASAP7_75t_L g317 ( 
.A1(n_212),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_196),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_218),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_213),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_220),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_224),
.B(n_16),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_217),
.A2(n_231),
.B1(n_232),
.B2(n_211),
.Y(n_323)
);

AND2x4_ASAP7_75t_L g324 ( 
.A(n_228),
.B(n_17),
.Y(n_324)
);

BUFx10_ASAP7_75t_L g325 ( 
.A(n_283),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_293),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_308),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_272),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_304),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_282),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_281),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_299),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_318),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_286),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_286),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_285),
.Y(n_336)
);

BUFx10_ASAP7_75t_L g337 ( 
.A(n_283),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_284),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_285),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_R g340 ( 
.A(n_320),
.B(n_202),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_270),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_290),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_291),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_284),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_270),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_291),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_291),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_303),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_283),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_323),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_319),
.Y(n_351)
);

NAND2xp33_ASAP7_75t_R g352 ( 
.A(n_320),
.B(n_197),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_307),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_310),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_301),
.B(n_239),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_R g356 ( 
.A(n_308),
.B(n_255),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_311),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_270),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_315),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_270),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_311),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_280),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_311),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_321),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_312),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_279),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_273),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_277),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_301),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_R g370 ( 
.A(n_302),
.B(n_255),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_312),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_301),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_312),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_301),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_309),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_312),
.Y(n_376)
);

BUFx8_ASAP7_75t_L g377 ( 
.A(n_271),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_313),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_353),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_365),
.B(n_275),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_371),
.B(n_275),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_373),
.B(n_275),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_366),
.Y(n_383)
);

XOR2x2_ASAP7_75t_L g384 ( 
.A(n_329),
.B(n_274),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_354),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_341),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_376),
.B(n_275),
.Y(n_387)
);

NAND2xp33_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_292),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_378),
.B(n_305),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_330),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_366),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_367),
.B(n_292),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_340),
.B(n_302),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_359),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_368),
.B(n_309),
.Y(n_395)
);

AND2x6_ASAP7_75t_SL g396 ( 
.A(n_350),
.B(n_322),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_341),
.B(n_305),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_346),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_364),
.B(n_309),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_374),
.B(n_309),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_345),
.B(n_324),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_327),
.B(n_189),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_345),
.B(n_324),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_346),
.B(n_271),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_343),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_349),
.B(n_263),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_347),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_333),
.B(n_269),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_336),
.Y(n_409)
);

NOR3xp33_ASAP7_75t_L g410 ( 
.A(n_326),
.B(n_274),
.C(n_322),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_L g411 ( 
.A(n_332),
.B(n_198),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_331),
.B(n_306),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_325),
.B(n_278),
.Y(n_413)
);

NAND2xp33_ASAP7_75t_L g414 ( 
.A(n_356),
.B(n_276),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_357),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_361),
.B(n_294),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_363),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_355),
.B(n_306),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_330),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_358),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_336),
.Y(n_421)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_325),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_358),
.Y(n_423)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_325),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g425 ( 
.A(n_337),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_360),
.B(n_362),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_360),
.B(n_313),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_352),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_350),
.A2(n_294),
.B1(n_297),
.B2(n_317),
.Y(n_429)
);

AND2x4_ASAP7_75t_SL g430 ( 
.A(n_337),
.B(n_300),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_362),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_328),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_339),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_351),
.B(n_306),
.Y(n_434)
);

NOR2xp67_ASAP7_75t_L g435 ( 
.A(n_369),
.B(n_199),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_372),
.B(n_313),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_337),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_377),
.B(n_297),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_375),
.B(n_313),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_377),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_377),
.B(n_314),
.Y(n_441)
);

OAI22xp33_ASAP7_75t_L g442 ( 
.A1(n_342),
.A2(n_287),
.B1(n_268),
.B2(n_300),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_348),
.Y(n_443)
);

BUFx6f_ASAP7_75t_SL g444 ( 
.A(n_338),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_334),
.B(n_314),
.Y(n_445)
);

NAND2xp33_ASAP7_75t_L g446 ( 
.A(n_335),
.B(n_276),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_379),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_398),
.B(n_289),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_385),
.Y(n_449)
);

NOR2x1_ASAP7_75t_L g450 ( 
.A(n_414),
.B(n_268),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_398),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_404),
.B(n_241),
.Y(n_452)
);

AO22x2_ASAP7_75t_L g453 ( 
.A1(n_393),
.A2(n_288),
.B1(n_295),
.B2(n_287),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_388),
.A2(n_276),
.B1(n_242),
.B2(n_260),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_415),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_394),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_409),
.B(n_296),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_421),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_397),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_437),
.Y(n_460)
);

A2O1A1Ixp33_ASAP7_75t_L g461 ( 
.A1(n_392),
.A2(n_251),
.B(n_250),
.C(n_254),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_437),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_390),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_404),
.B(n_261),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_401),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_413),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_391),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_402),
.B(n_278),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_403),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_392),
.B(n_265),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_389),
.B(n_266),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_405),
.B(n_298),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_418),
.B(n_314),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_432),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_418),
.B(n_314),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_416),
.A2(n_276),
.B(n_201),
.Y(n_476)
);

NAND3xp33_ASAP7_75t_SL g477 ( 
.A(n_410),
.B(n_344),
.C(n_338),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_428),
.B(n_204),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_437),
.B(n_209),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_407),
.B(n_298),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_408),
.Y(n_481)
);

NOR2xp67_ASAP7_75t_L g482 ( 
.A(n_436),
.B(n_28),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_390),
.Y(n_483)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_437),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_408),
.B(n_210),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_439),
.B(n_316),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_393),
.A2(n_247),
.B1(n_219),
.B2(n_221),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_411),
.B(n_395),
.Y(n_488)
);

O2A1O1Ixp5_ASAP7_75t_L g489 ( 
.A1(n_402),
.A2(n_276),
.B(n_316),
.C(n_245),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_416),
.A2(n_249),
.B1(n_222),
.B2(n_226),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_419),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_395),
.B(n_316),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_426),
.A2(n_256),
.B(n_230),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_419),
.Y(n_494)
);

AND2x6_ASAP7_75t_SL g495 ( 
.A(n_443),
.B(n_344),
.Y(n_495)
);

NAND2xp33_ASAP7_75t_SL g496 ( 
.A(n_438),
.B(n_215),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_417),
.B(n_233),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_429),
.A2(n_257),
.B1(n_267),
.B2(n_264),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_433),
.B(n_234),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_430),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_422),
.B(n_236),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_423),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_423),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_400),
.B(n_386),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_431),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_383),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_438),
.B(n_237),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_431),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_420),
.B(n_316),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_427),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_430),
.B(n_238),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_434),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_445),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_442),
.B(n_252),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_434),
.Y(n_515)
);

NAND2x1p5_ASAP7_75t_L g516 ( 
.A(n_424),
.B(n_280),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_481),
.A2(n_425),
.B1(n_441),
.B2(n_440),
.Y(n_517)
);

AND2x2_ASAP7_75t_SL g518 ( 
.A(n_507),
.B(n_446),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_513),
.B(n_406),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_450),
.A2(n_486),
.B(n_484),
.Y(n_520)
);

A2O1A1Ixp33_ASAP7_75t_SL g521 ( 
.A1(n_485),
.A2(n_399),
.B(n_412),
.C(n_387),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_459),
.B(n_406),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_463),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_460),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_483),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_503),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_465),
.B(n_435),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_469),
.A2(n_470),
.B1(n_466),
.B2(n_507),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_460),
.Y(n_529)
);

OA22x2_ASAP7_75t_L g530 ( 
.A1(n_498),
.A2(n_384),
.B1(n_396),
.B2(n_444),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_455),
.B(n_444),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_506),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_460),
.Y(n_533)
);

A2O1A1Ixp33_ASAP7_75t_SL g534 ( 
.A1(n_476),
.A2(n_399),
.B(n_412),
.C(n_382),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_467),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_512),
.B(n_258),
.Y(n_536)
);

INVx3_ASAP7_75t_SL g537 ( 
.A(n_468),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_515),
.B(n_262),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_462),
.B(n_280),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_450),
.A2(n_381),
.B(n_380),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_451),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_472),
.B(n_18),
.Y(n_542)
);

NAND2xp33_ASAP7_75t_SL g543 ( 
.A(n_462),
.B(n_280),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_472),
.B(n_19),
.Y(n_544)
);

NOR2x1_ASAP7_75t_SL g545 ( 
.A(n_462),
.B(n_31),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_484),
.A2(n_103),
.B1(n_182),
.B2(n_180),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_510),
.B(n_471),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_480),
.B(n_448),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_514),
.A2(n_99),
.B1(n_179),
.B2(n_177),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_488),
.A2(n_96),
.B1(n_175),
.B2(n_174),
.Y(n_550)
);

OAI21x1_ASAP7_75t_L g551 ( 
.A1(n_503),
.A2(n_183),
.B(n_93),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_452),
.B(n_19),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_504),
.A2(n_95),
.B(n_172),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_491),
.Y(n_554)
);

BUFx4f_ASAP7_75t_L g555 ( 
.A(n_500),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_448),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_464),
.B(n_20),
.Y(n_557)
);

A2O1A1Ixp33_ASAP7_75t_L g558 ( 
.A1(n_461),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_473),
.A2(n_92),
.B(n_171),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_447),
.B(n_21),
.Y(n_560)
);

O2A1O1Ixp5_ASAP7_75t_L g561 ( 
.A1(n_489),
.A2(n_102),
.B(n_165),
.C(n_164),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_R g562 ( 
.A(n_496),
.B(n_33),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_494),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_449),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_456),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_478),
.B(n_22),
.Y(n_566)
);

OAI21xp33_ASAP7_75t_SL g567 ( 
.A1(n_458),
.A2(n_23),
.B(n_24),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_475),
.A2(n_88),
.B(n_162),
.Y(n_568)
);

OAI21xp33_ASAP7_75t_SL g569 ( 
.A1(n_454),
.A2(n_23),
.B(n_24),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_457),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_487),
.A2(n_104),
.B1(n_161),
.B2(n_36),
.Y(n_571)
);

O2A1O1Ixp33_ASAP7_75t_L g572 ( 
.A1(n_493),
.A2(n_25),
.B(n_26),
.C(n_37),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_457),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_480),
.Y(n_574)
);

BUFx4f_ASAP7_75t_SL g575 ( 
.A(n_497),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_492),
.B(n_474),
.Y(n_576)
);

BUFx4f_ASAP7_75t_SL g577 ( 
.A(n_532),
.Y(n_577)
);

AOI22x1_ASAP7_75t_L g578 ( 
.A1(n_540),
.A2(n_520),
.B1(n_553),
.B2(n_523),
.Y(n_578)
);

AOI22x1_ASAP7_75t_L g579 ( 
.A1(n_525),
.A2(n_502),
.B1(n_508),
.B2(n_516),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_535),
.B(n_477),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_547),
.B(n_511),
.Y(n_581)
);

AOI21x1_ASAP7_75t_L g582 ( 
.A1(n_576),
.A2(n_554),
.B(n_563),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_548),
.Y(n_583)
);

OA21x2_ASAP7_75t_L g584 ( 
.A1(n_561),
.A2(n_509),
.B(n_482),
.Y(n_584)
);

BUFx8_ASAP7_75t_L g585 ( 
.A(n_570),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_524),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_524),
.Y(n_587)
);

CKINVDCx11_ASAP7_75t_R g588 ( 
.A(n_537),
.Y(n_588)
);

OAI21x1_ASAP7_75t_L g589 ( 
.A1(n_551),
.A2(n_505),
.B(n_482),
.Y(n_589)
);

OAI21x1_ASAP7_75t_L g590 ( 
.A1(n_559),
.A2(n_505),
.B(n_479),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_541),
.B(n_499),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_519),
.B(n_499),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_564),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_565),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_574),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_526),
.Y(n_596)
);

AO21x2_ASAP7_75t_L g597 ( 
.A1(n_521),
.A2(n_501),
.B(n_490),
.Y(n_597)
);

AOI21x1_ASAP7_75t_L g598 ( 
.A1(n_527),
.A2(n_453),
.B(n_38),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_560),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_556),
.Y(n_600)
);

OAI21x1_ASAP7_75t_L g601 ( 
.A1(n_568),
.A2(n_112),
.B(n_41),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_524),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_529),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_529),
.Y(n_604)
);

OAI21x1_ASAP7_75t_L g605 ( 
.A1(n_572),
.A2(n_113),
.B(n_43),
.Y(n_605)
);

OAI21x1_ASAP7_75t_L g606 ( 
.A1(n_539),
.A2(n_115),
.B(n_44),
.Y(n_606)
);

OAI21x1_ASAP7_75t_SL g607 ( 
.A1(n_545),
.A2(n_116),
.B(n_46),
.Y(n_607)
);

INVxp67_ASAP7_75t_SL g608 ( 
.A(n_529),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_533),
.Y(n_609)
);

INVx3_ASAP7_75t_SL g610 ( 
.A(n_518),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_533),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_533),
.Y(n_612)
);

OAI21x1_ASAP7_75t_L g613 ( 
.A1(n_550),
.A2(n_117),
.B(n_47),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_522),
.A2(n_453),
.B(n_48),
.Y(n_614)
);

OR2x6_ASAP7_75t_L g615 ( 
.A(n_570),
.B(n_495),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_570),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_542),
.Y(n_617)
);

INVx1_ASAP7_75t_SL g618 ( 
.A(n_544),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_573),
.Y(n_619)
);

INVx5_ASAP7_75t_L g620 ( 
.A(n_573),
.Y(n_620)
);

NAND2x1p5_ASAP7_75t_L g621 ( 
.A(n_573),
.B(n_119),
.Y(n_621)
);

AO21x2_ASAP7_75t_L g622 ( 
.A1(n_534),
.A2(n_109),
.B(n_49),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_575),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_528),
.B(n_121),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_577),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_581),
.B(n_536),
.Y(n_626)
);

AOI21x1_ASAP7_75t_L g627 ( 
.A1(n_582),
.A2(n_552),
.B(n_557),
.Y(n_627)
);

OAI22xp33_ASAP7_75t_L g628 ( 
.A1(n_610),
.A2(n_530),
.B1(n_531),
.B2(n_566),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_599),
.B(n_538),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_614),
.A2(n_567),
.B1(n_569),
.B2(n_571),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_624),
.A2(n_517),
.B1(n_555),
.B2(n_549),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_593),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_624),
.A2(n_567),
.B1(n_569),
.B2(n_562),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_594),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_592),
.B(n_555),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_596),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_624),
.A2(n_546),
.B1(n_558),
.B2(n_543),
.Y(n_637)
);

INVx6_ASAP7_75t_L g638 ( 
.A(n_585),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_577),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_596),
.Y(n_640)
);

CKINVDCx11_ASAP7_75t_R g641 ( 
.A(n_588),
.Y(n_641)
);

AOI21xp33_ASAP7_75t_SL g642 ( 
.A1(n_580),
.A2(n_25),
.B(n_53),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_578),
.A2(n_54),
.B(n_56),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_610),
.A2(n_591),
.B1(n_618),
.B2(n_623),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_604),
.Y(n_645)
);

CKINVDCx11_ASAP7_75t_R g646 ( 
.A(n_588),
.Y(n_646)
);

OA21x2_ASAP7_75t_L g647 ( 
.A1(n_605),
.A2(n_58),
.B(n_62),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_585),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_620),
.A2(n_63),
.B1(n_68),
.B2(n_69),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_583),
.B(n_70),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_583),
.B(n_71),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_601),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_597),
.A2(n_72),
.B1(n_73),
.B2(n_75),
.Y(n_653)
);

OAI22xp33_ASAP7_75t_L g654 ( 
.A1(n_580),
.A2(n_77),
.B1(n_80),
.B2(n_81),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_602),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_604),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_L g657 ( 
.A1(n_590),
.A2(n_82),
.B(n_83),
.Y(n_657)
);

OR2x6_ASAP7_75t_L g658 ( 
.A(n_619),
.B(n_84),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_612),
.Y(n_659)
);

INVx6_ASAP7_75t_L g660 ( 
.A(n_585),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_600),
.Y(n_661)
);

OAI21x1_ASAP7_75t_L g662 ( 
.A1(n_589),
.A2(n_86),
.B(n_105),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_608),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_604),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_616),
.Y(n_665)
);

OAI22xp5_ASAP7_75t_L g666 ( 
.A1(n_620),
.A2(n_123),
.B1(n_126),
.B2(n_128),
.Y(n_666)
);

OAI21xp5_ASAP7_75t_SL g667 ( 
.A1(n_591),
.A2(n_130),
.B(n_131),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_591),
.B(n_173),
.Y(n_668)
);

AOI21x1_ASAP7_75t_L g669 ( 
.A1(n_589),
.A2(n_133),
.B(n_136),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_628),
.A2(n_617),
.B1(n_597),
.B2(n_615),
.Y(n_670)
);

INVxp33_ASAP7_75t_L g671 ( 
.A(n_644),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_668),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_626),
.B(n_598),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_668),
.B(n_661),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_663),
.Y(n_675)
);

NAND2xp33_ASAP7_75t_R g676 ( 
.A(n_635),
.B(n_595),
.Y(n_676)
);

OAI22xp5_ASAP7_75t_L g677 ( 
.A1(n_633),
.A2(n_620),
.B1(n_615),
.B2(n_619),
.Y(n_677)
);

INVxp67_ASAP7_75t_L g678 ( 
.A(n_632),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_638),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_629),
.B(n_628),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_634),
.B(n_615),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_636),
.B(n_615),
.Y(n_682)
);

NOR3xp33_ASAP7_75t_SL g683 ( 
.A(n_667),
.B(n_654),
.C(n_650),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_640),
.B(n_611),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_655),
.Y(n_685)
);

NAND2xp33_ASAP7_75t_R g686 ( 
.A(n_647),
.B(n_613),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_631),
.B(n_620),
.Y(n_687)
);

NAND2xp33_ASAP7_75t_SL g688 ( 
.A(n_625),
.B(n_604),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_633),
.B(n_620),
.Y(n_689)
);

AND2x4_ASAP7_75t_SL g690 ( 
.A(n_639),
.B(n_586),
.Y(n_690)
);

NAND3xp33_ASAP7_75t_L g691 ( 
.A(n_630),
.B(n_579),
.C(n_584),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_630),
.B(n_605),
.Y(n_692)
);

NAND2xp33_ASAP7_75t_R g693 ( 
.A(n_647),
.B(n_613),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_645),
.Y(n_694)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_656),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_659),
.Y(n_696)
);

XOR2xp5_ASAP7_75t_L g697 ( 
.A(n_648),
.B(n_621),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_665),
.Y(n_698)
);

AO31x2_ASAP7_75t_L g699 ( 
.A1(n_652),
.A2(n_622),
.A3(n_584),
.B(n_586),
.Y(n_699)
);

INVxp67_ASAP7_75t_SL g700 ( 
.A(n_664),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_658),
.B(n_603),
.Y(n_701)
);

INVx4_ASAP7_75t_L g702 ( 
.A(n_638),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_654),
.A2(n_637),
.B1(n_653),
.B2(n_638),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_651),
.B(n_648),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_658),
.B(n_603),
.Y(n_705)
);

AND2x4_ASAP7_75t_SL g706 ( 
.A(n_658),
.B(n_586),
.Y(n_706)
);

CKINVDCx16_ASAP7_75t_R g707 ( 
.A(n_641),
.Y(n_707)
);

NOR3xp33_ASAP7_75t_SL g708 ( 
.A(n_649),
.B(n_607),
.C(n_621),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_642),
.B(n_611),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_660),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_641),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_637),
.B(n_609),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_646),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_657),
.B(n_609),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_646),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_652),
.B(n_587),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_627),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_653),
.B(n_587),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_R g719 ( 
.A(n_660),
.B(n_587),
.Y(n_719)
);

NAND2xp33_ASAP7_75t_SL g720 ( 
.A(n_660),
.B(n_622),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_717),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_680),
.B(n_647),
.Y(n_722)
);

INVx4_ASAP7_75t_L g723 ( 
.A(n_712),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_674),
.B(n_643),
.Y(n_724)
);

NOR2x1_ASAP7_75t_R g725 ( 
.A(n_711),
.B(n_713),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_698),
.B(n_606),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_685),
.B(n_606),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_696),
.B(n_662),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_716),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_699),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_675),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_678),
.B(n_601),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_692),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_673),
.B(n_669),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_694),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_710),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_692),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_673),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_671),
.B(n_666),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_691),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_687),
.B(n_670),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_712),
.B(n_590),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_676),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_703),
.A2(n_584),
.B1(n_139),
.B2(n_140),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_716),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_695),
.B(n_138),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_691),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_714),
.B(n_159),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_714),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_677),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_677),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_672),
.B(n_142),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_700),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_681),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_672),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_689),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_684),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_682),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_721),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_731),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_749),
.B(n_702),
.Y(n_761)
);

OA21x2_ASAP7_75t_L g762 ( 
.A1(n_740),
.A2(n_708),
.B(n_718),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_749),
.B(n_704),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_721),
.Y(n_764)
);

OAI221xp5_ASAP7_75t_SL g765 ( 
.A1(n_743),
.A2(n_697),
.B1(n_709),
.B2(n_683),
.C(n_679),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_758),
.B(n_701),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_749),
.B(n_705),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_756),
.B(n_705),
.Y(n_768)
);

OR2x2_ASAP7_75t_L g769 ( 
.A(n_733),
.B(n_720),
.Y(n_769)
);

INVx1_ASAP7_75t_SL g770 ( 
.A(n_731),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_730),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_733),
.B(n_702),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_756),
.B(n_706),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_756),
.B(n_690),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_721),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_758),
.B(n_707),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_738),
.B(n_688),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_738),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_758),
.B(n_715),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_740),
.B(n_144),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_757),
.B(n_719),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_730),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_757),
.B(n_147),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_735),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_737),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_737),
.B(n_693),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_SL g787 ( 
.A1(n_744),
.A2(n_686),
.B(n_152),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_763),
.B(n_747),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_763),
.B(n_747),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_786),
.B(n_747),
.Y(n_790)
);

BUFx2_ASAP7_75t_L g791 ( 
.A(n_760),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_775),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_778),
.Y(n_793)
);

AND2x4_ASAP7_75t_L g794 ( 
.A(n_760),
.B(n_729),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_786),
.B(n_767),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_767),
.B(n_742),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_759),
.B(n_742),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_775),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_784),
.B(n_754),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_770),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_759),
.B(n_722),
.Y(n_801)
);

NAND2x1p5_ASAP7_75t_L g802 ( 
.A(n_762),
.B(n_723),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_759),
.B(n_722),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_779),
.B(n_736),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_766),
.B(n_757),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_764),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_770),
.B(n_741),
.Y(n_807)
);

OR2x6_ASAP7_75t_L g808 ( 
.A(n_802),
.B(n_761),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_792),
.Y(n_809)
);

AOI32xp33_ASAP7_75t_L g810 ( 
.A1(n_790),
.A2(n_776),
.A3(n_780),
.B1(n_748),
.B2(n_768),
.Y(n_810)
);

O2A1O1Ixp5_ASAP7_75t_R g811 ( 
.A1(n_807),
.A2(n_799),
.B(n_777),
.C(n_781),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_792),
.Y(n_812)
);

A2O1A1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_804),
.A2(n_787),
.B(n_765),
.C(n_739),
.Y(n_813)
);

OR2x2_ASAP7_75t_L g814 ( 
.A(n_795),
.B(n_790),
.Y(n_814)
);

NOR3xp33_ASAP7_75t_L g815 ( 
.A(n_800),
.B(n_787),
.C(n_783),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_795),
.B(n_789),
.Y(n_816)
);

OAI31xp33_ASAP7_75t_L g817 ( 
.A1(n_802),
.A2(n_776),
.A3(n_748),
.B(n_780),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_791),
.Y(n_818)
);

NOR2x1p5_ASAP7_75t_SL g819 ( 
.A(n_806),
.B(n_782),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_788),
.B(n_768),
.Y(n_820)
);

OAI21xp33_ASAP7_75t_L g821 ( 
.A1(n_811),
.A2(n_777),
.B(n_805),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_813),
.B(n_725),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_815),
.A2(n_802),
.B(n_793),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_809),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_SL g825 ( 
.A1(n_808),
.A2(n_762),
.B1(n_723),
.B2(n_736),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_SL g826 ( 
.A1(n_808),
.A2(n_762),
.B1(n_723),
.B2(n_736),
.Y(n_826)
);

AOI31xp33_ASAP7_75t_L g827 ( 
.A1(n_814),
.A2(n_725),
.A3(n_818),
.B(n_816),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_822),
.A2(n_817),
.B(n_810),
.C(n_819),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_824),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_SL g830 ( 
.A1(n_823),
.A2(n_762),
.B1(n_827),
.B2(n_723),
.Y(n_830)
);

AOI221xp5_ASAP7_75t_L g831 ( 
.A1(n_821),
.A2(n_812),
.B1(n_809),
.B2(n_788),
.C(n_789),
.Y(n_831)
);

INVx1_ASAP7_75t_SL g832 ( 
.A(n_825),
.Y(n_832)
);

NAND3xp33_ASAP7_75t_L g833 ( 
.A(n_826),
.B(n_772),
.C(n_774),
.Y(n_833)
);

AOI221xp5_ASAP7_75t_L g834 ( 
.A1(n_832),
.A2(n_791),
.B1(n_820),
.B2(n_798),
.C(n_801),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_831),
.B(n_796),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_829),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_833),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_828),
.B(n_796),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_837),
.B(n_830),
.Y(n_839)
);

OA22x2_ASAP7_75t_L g840 ( 
.A1(n_835),
.A2(n_794),
.B1(n_798),
.B2(n_761),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_838),
.A2(n_724),
.B(n_732),
.Y(n_841)
);

NAND4xp25_ASAP7_75t_L g842 ( 
.A(n_839),
.B(n_834),
.C(n_836),
.D(n_741),
.Y(n_842)
);

AOI221xp5_ASAP7_75t_L g843 ( 
.A1(n_841),
.A2(n_785),
.B1(n_794),
.B2(n_750),
.C(n_751),
.Y(n_843)
);

XNOR2xp5_ASAP7_75t_L g844 ( 
.A(n_840),
.B(n_774),
.Y(n_844)
);

OAI211xp5_ASAP7_75t_L g845 ( 
.A1(n_839),
.A2(n_772),
.B(n_746),
.C(n_769),
.Y(n_845)
);

NOR2x1_ASAP7_75t_L g846 ( 
.A(n_842),
.B(n_752),
.Y(n_846)
);

NOR2xp67_ASAP7_75t_L g847 ( 
.A(n_845),
.B(n_844),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_843),
.B(n_797),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_842),
.A2(n_794),
.B1(n_761),
.B2(n_773),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_842),
.B(n_803),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_844),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_843),
.B(n_803),
.Y(n_852)
);

OAI32xp33_ASAP7_75t_L g853 ( 
.A1(n_851),
.A2(n_769),
.A3(n_750),
.B1(n_751),
.B2(n_785),
.Y(n_853)
);

NOR2x1p5_ASAP7_75t_L g854 ( 
.A(n_850),
.B(n_752),
.Y(n_854)
);

NOR2x1p5_ASAP7_75t_L g855 ( 
.A(n_852),
.B(n_752),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_848),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_847),
.Y(n_857)
);

NOR4xp75_ASAP7_75t_SL g858 ( 
.A(n_846),
.B(n_752),
.C(n_746),
.D(n_755),
.Y(n_858)
);

XNOR2x1_ASAP7_75t_L g859 ( 
.A(n_849),
.B(n_148),
.Y(n_859)
);

OAI211xp5_ASAP7_75t_SL g860 ( 
.A1(n_851),
.A2(n_753),
.B(n_778),
.C(n_806),
.Y(n_860)
);

NOR4xp25_ASAP7_75t_L g861 ( 
.A(n_851),
.B(n_753),
.C(n_728),
.D(n_727),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_857),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_856),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_854),
.B(n_797),
.Y(n_864)
);

OAI21xp33_ASAP7_75t_SL g865 ( 
.A1(n_855),
.A2(n_801),
.B(n_773),
.Y(n_865)
);

INVx1_ASAP7_75t_SL g866 ( 
.A(n_859),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_858),
.Y(n_867)
);

INVx1_ASAP7_75t_SL g868 ( 
.A(n_853),
.Y(n_868)
);

CKINVDCx20_ASAP7_75t_R g869 ( 
.A(n_860),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_863),
.Y(n_870)
);

INVxp67_ASAP7_75t_L g871 ( 
.A(n_862),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_869),
.A2(n_866),
.B1(n_868),
.B2(n_867),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_869),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_864),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_865),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_862),
.B(n_861),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_862),
.B(n_761),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_862),
.A2(n_771),
.B1(n_755),
.B2(n_729),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_L g879 ( 
.A1(n_862),
.A2(n_771),
.B1(n_755),
.B2(n_729),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_873),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_875),
.Y(n_881)
);

BUFx2_ASAP7_75t_SL g882 ( 
.A(n_870),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_872),
.B(n_764),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_871),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_874),
.Y(n_885)
);

INVx3_ASAP7_75t_SL g886 ( 
.A(n_877),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_876),
.B(n_764),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_878),
.A2(n_755),
.B1(n_729),
.B2(n_727),
.Y(n_888)
);

AOI31xp33_ASAP7_75t_L g889 ( 
.A1(n_879),
.A2(n_154),
.A3(n_155),
.B(n_157),
.Y(n_889)
);

INVxp67_ASAP7_75t_L g890 ( 
.A(n_880),
.Y(n_890)
);

INVxp67_ASAP7_75t_L g891 ( 
.A(n_882),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_884),
.Y(n_892)
);

XOR2x1_ASAP7_75t_L g893 ( 
.A(n_881),
.B(n_158),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_885),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_883),
.A2(n_887),
.B(n_889),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_892),
.Y(n_896)
);

OAI22x1_ASAP7_75t_L g897 ( 
.A1(n_890),
.A2(n_886),
.B1(n_891),
.B2(n_894),
.Y(n_897)
);

AOI222xp33_ASAP7_75t_L g898 ( 
.A1(n_893),
.A2(n_888),
.B1(n_889),
.B2(n_734),
.C1(n_728),
.C2(n_726),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_896),
.A2(n_895),
.B(n_734),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_897),
.B(n_755),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_SL g901 ( 
.A1(n_900),
.A2(n_898),
.B1(n_755),
.B2(n_726),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_901),
.B(n_899),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_902),
.A2(n_771),
.B1(n_782),
.B2(n_745),
.Y(n_903)
);


endmodule