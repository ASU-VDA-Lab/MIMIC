module fake_jpeg_26631_n_182 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_182);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_182;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_8),
.B(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_34),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_43),
.Y(n_47)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_25),
.B1(n_15),
.B2(n_24),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_49),
.A2(n_15),
.B1(n_18),
.B2(n_36),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_30),
.B1(n_23),
.B2(n_31),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_59),
.B1(n_18),
.B2(n_32),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_38),
.A2(n_30),
.B1(n_23),
.B2(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_34),
.B(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_28),
.Y(n_73)
);

NOR2x1_ASAP7_75t_R g62 ( 
.A(n_45),
.B(n_25),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_20),
.B(n_17),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_37),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_77),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_57),
.A2(n_39),
.B1(n_49),
.B2(n_53),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_64),
.A2(n_69),
.B1(n_58),
.B2(n_3),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_65),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_67),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_21),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_24),
.B1(n_20),
.B2(n_17),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_71),
.A2(n_82),
.B1(n_54),
.B2(n_58),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_48),
.B(n_28),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_72),
.B(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_26),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_78),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_26),
.B1(n_15),
.B2(n_29),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_54),
.C(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_29),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_84),
.B1(n_79),
.B2(n_68),
.Y(n_100)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_35),
.B1(n_42),
.B2(n_15),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_29),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_54),
.B(n_10),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_51),
.A2(n_24),
.B1(n_20),
.B2(n_17),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_85),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_89),
.B(n_96),
.Y(n_114)
);

NOR2x1_ASAP7_75t_SL g118 ( 
.A(n_94),
.B(n_82),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_63),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_97),
.B(n_103),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_101),
.B1(n_69),
.B2(n_80),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_107),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_68),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_123),
.Y(n_139)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_111),
.B(n_116),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_104),
.B(n_88),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_113),
.B(n_124),
.Y(n_130)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_122),
.Y(n_141)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_117),
.B(n_119),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_82),
.B(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_121),
.A2(n_102),
.B1(n_90),
.B2(n_96),
.Y(n_132)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_103),
.B(n_108),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_127),
.A2(n_137),
.B(n_140),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_97),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_121),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_125),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_133),
.Y(n_152)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_62),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_112),
.B(n_71),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_92),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

NOR4xp25_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_74),
.C(n_61),
.D(n_70),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_109),
.C(n_118),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_142),
.B(n_143),
.Y(n_157)
);

HAxp5_ASAP7_75t_SL g143 ( 
.A(n_127),
.B(n_109),
.CON(n_143),
.SN(n_143)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_147),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_132),
.C(n_133),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_149),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_95),
.C(n_9),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_1),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_146),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_154),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_151),
.A2(n_139),
.B1(n_143),
.B2(n_144),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_152),
.B(n_130),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_160),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_150),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_164),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_142),
.C(n_134),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_136),
.C(n_128),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_168),
.C(n_13),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_128),
.C(n_138),
.Y(n_168)
);

A2O1A1O1Ixp25_ASAP7_75t_L g169 ( 
.A1(n_162),
.A2(n_154),
.B(n_159),
.C(n_161),
.D(n_10),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_169),
.A2(n_165),
.B(n_172),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_95),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_171),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_165),
.A2(n_13),
.B1(n_5),
.B2(n_6),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_4),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_174),
.A2(n_175),
.B(n_177),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_173),
.A2(n_4),
.B(n_5),
.Y(n_177)
);

AOI21x1_ASAP7_75t_L g179 ( 
.A1(n_176),
.A2(n_169),
.B(n_170),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_179),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_SL g181 ( 
.A1(n_180),
.A2(n_178),
.B(n_5),
.C(n_6),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_4),
.Y(n_182)
);


endmodule