module fake_jpeg_16689_n_263 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_263);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_263;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_7),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_19),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_50),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_24),
.C(n_20),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_60),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_19),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_27),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_22),
.B1(n_33),
.B2(n_31),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_35),
.A2(n_22),
.B1(n_27),
.B2(n_33),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_28),
.B1(n_23),
.B2(n_16),
.Y(n_77)
);

CKINVDCx9p33_ASAP7_75t_R g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_26),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_18),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_61),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_33),
.B1(n_22),
.B2(n_31),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_64),
.A2(n_32),
.B1(n_29),
.B2(n_52),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_42),
.C(n_21),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_65),
.A2(n_73),
.B1(n_59),
.B2(n_46),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_66),
.B(n_78),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_0),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_68),
.A2(n_77),
.B1(n_0),
.B2(n_1),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_28),
.B1(n_31),
.B2(n_29),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_11),
.C(n_13),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_44),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_50),
.A2(n_32),
.B(n_23),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_79),
.A2(n_32),
.B(n_21),
.Y(n_106)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_83),
.Y(n_89)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_86),
.B(n_87),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_72),
.A2(n_54),
.B1(n_45),
.B2(n_47),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_88),
.A2(n_91),
.B1(n_96),
.B2(n_71),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_59),
.B(n_57),
.C(n_43),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_106),
.B(n_107),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_86),
.A2(n_66),
.B1(n_65),
.B2(n_73),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_70),
.A2(n_28),
.B1(n_45),
.B2(n_47),
.Y(n_94)
);

AO21x1_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_98),
.B(n_99),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_102),
.B1(n_80),
.B2(n_68),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_78),
.A2(n_53),
.B1(n_55),
.B2(n_52),
.Y(n_96)
);

OAI21xp33_ASAP7_75t_SL g98 ( 
.A1(n_79),
.A2(n_26),
.B(n_20),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_70),
.A2(n_24),
.B1(n_55),
.B2(n_29),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_104),
.B(n_68),
.Y(n_115)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

AOI32xp33_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_29),
.A3(n_17),
.B1(n_18),
.B2(n_21),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_109),
.B(n_75),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_67),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_113),
.B(n_123),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_114),
.A2(n_117),
.B1(n_84),
.B2(n_7),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_115),
.B(n_116),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_80),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_80),
.B1(n_77),
.B2(n_68),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_118),
.A2(n_135),
.B1(n_104),
.B2(n_107),
.Y(n_144)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_67),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_92),
.B(n_103),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_132),
.B(n_106),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_82),
.Y(n_126)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_81),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_128),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_75),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_108),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_130),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_97),
.B(n_17),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_97),
.B(n_17),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_133),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_96),
.B(n_85),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_83),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_137),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_88),
.A2(n_52),
.B1(n_84),
.B2(n_74),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_89),
.B(n_21),
.C(n_32),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_32),
.C(n_101),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_90),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_146),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_147),
.C(n_149),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_124),
.B1(n_119),
.B2(n_115),
.Y(n_167)
);

AND2x2_ASAP7_75t_SL g145 ( 
.A(n_127),
.B(n_101),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_2),
.B(n_4),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_93),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_93),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_114),
.A2(n_105),
.B1(n_84),
.B2(n_93),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_148),
.A2(n_159),
.B1(n_160),
.B2(n_123),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_21),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_121),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_154),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_152),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_100),
.C(n_18),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_155),
.A2(n_125),
.B1(n_124),
.B2(n_129),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_158),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_132),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_119),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_163),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_166),
.B(n_168),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_167),
.A2(n_171),
.B(n_172),
.Y(n_201)
);

XNOR2x1_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_117),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_124),
.B(n_122),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_164),
.A2(n_135),
.B1(n_136),
.B2(n_133),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_173),
.A2(n_176),
.B1(n_183),
.B2(n_186),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_164),
.A2(n_136),
.B1(n_112),
.B2(n_120),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_161),
.A2(n_112),
.B(n_120),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_153),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_SL g190 ( 
.A1(n_178),
.A2(n_157),
.B(n_159),
.C(n_160),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_139),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_4),
.Y(n_180)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_145),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_140),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_185),
.Y(n_189)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_146),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_5),
.B1(n_8),
.B2(n_10),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_188),
.A2(n_186),
.B1(n_166),
.B2(n_180),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_190),
.A2(n_207),
.B1(n_183),
.B2(n_188),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_182),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_191),
.B(n_194),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

NOR3xp33_ASAP7_75t_SL g194 ( 
.A(n_172),
.B(n_141),
.C(n_157),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_140),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_196),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_175),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_208),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_139),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_198),
.B(n_204),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_167),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_202),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_170),
.B(n_151),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_147),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_171),
.B1(n_187),
.B2(n_165),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_210),
.A2(n_217),
.B1(n_218),
.B2(n_221),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_189),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_205),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_181),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_201),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_196),
.A2(n_171),
.B1(n_165),
.B2(n_169),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_208),
.A2(n_169),
.B1(n_168),
.B2(n_174),
.Y(n_218)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_219),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_192),
.A2(n_173),
.B1(n_176),
.B2(n_174),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_178),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

BUFx24_ASAP7_75t_SL g224 ( 
.A(n_209),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_224),
.B(n_229),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_223),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_227),
.B(n_228),
.Y(n_236)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_223),
.Y(n_228)
);

FAx1_ASAP7_75t_SL g229 ( 
.A(n_218),
.B(n_202),
.CI(n_194),
.CON(n_229),
.SN(n_229)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_232),
.C(n_234),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_201),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_233),
.A2(n_216),
.B(n_205),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_215),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_226),
.A2(n_213),
.B(n_217),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_190),
.Y(n_248)
);

INVx11_ASAP7_75t_L g238 ( 
.A(n_229),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_238),
.B(n_240),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_225),
.A2(n_222),
.B(n_214),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_210),
.C(n_207),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_231),
.A2(n_214),
.B1(n_221),
.B2(n_220),
.Y(n_240)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_241),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_203),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_238),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_243),
.B(n_206),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_235),
.C(n_148),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_248),
.A2(n_237),
.B1(n_239),
.B2(n_236),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_242),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_250),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_247),
.A2(n_150),
.B1(n_241),
.B2(n_151),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_252),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_253),
.A2(n_244),
.B(n_246),
.Y(n_254)
);

A2O1A1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_252),
.A2(n_248),
.B(n_146),
.C(n_144),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_253),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_257),
.A2(n_8),
.B(n_10),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_256),
.Y(n_260)
);

AOI322xp5_ASAP7_75t_L g261 ( 
.A1(n_260),
.A2(n_11),
.A3(n_12),
.B1(n_15),
.B2(n_258),
.C1(n_254),
.C2(n_257),
.Y(n_261)
);

BUFx24_ASAP7_75t_SL g262 ( 
.A(n_261),
.Y(n_262)
);

BUFx24_ASAP7_75t_SL g263 ( 
.A(n_262),
.Y(n_263)
);


endmodule