module fake_jpeg_29481_n_145 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_145);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_23),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_2),
.B(n_25),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_3),
.B(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_35),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g58 ( 
.A(n_49),
.B(n_1),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_47),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_55),
.Y(n_65)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_56),
.B(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_74),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_67),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_35),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_46),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_75),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_71),
.B(n_36),
.Y(n_81)
);

CKINVDCx6p67_ASAP7_75t_R g72 ( 
.A(n_59),
.Y(n_72)
);

INVxp67_ASAP7_75t_SL g84 ( 
.A(n_72),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_57),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_51),
.Y(n_75)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_81),
.Y(n_99)
);

AO22x2_ASAP7_75t_L g78 ( 
.A1(n_66),
.A2(n_38),
.B1(n_53),
.B2(n_48),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_88),
.Y(n_111)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_73),
.A2(n_70),
.B1(n_76),
.B2(n_38),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_50),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_90),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_69),
.B(n_63),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_89),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_42),
.B1(n_39),
.B2(n_41),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_44),
.B1(n_37),
.B2(n_34),
.Y(n_89)
);

BUFx4f_ASAP7_75t_SL g90 ( 
.A(n_72),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_63),
.A2(n_22),
.B1(n_32),
.B2(n_31),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_93),
.Y(n_100)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_1),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_3),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_6),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_5),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_98),
.B(n_102),
.Y(n_118)
);

AND2x4_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_5),
.Y(n_101)
);

NOR3xp33_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_109),
.C(n_115),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_89),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_6),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_7),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_112),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_SL g109 ( 
.A1(n_78),
.A2(n_90),
.B(n_84),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_33),
.B(n_11),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_110),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_82),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_30),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_114),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_8),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_13),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_119),
.B(n_126),
.Y(n_135)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_121),
.Y(n_132)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_14),
.C(n_15),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_123),
.B(n_101),
.Y(n_131)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_105),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_129),
.A2(n_101),
.B(n_96),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_96),
.B(n_100),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_131),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_117),
.Y(n_138)
);

AO221x1_ASAP7_75t_L g137 ( 
.A1(n_133),
.A2(n_116),
.B1(n_128),
.B2(n_109),
.C(n_117),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_138),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_128),
.B1(n_135),
.B2(n_136),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_132),
.C(n_125),
.Y(n_142)
);

BUFx24_ASAP7_75t_SL g143 ( 
.A(n_142),
.Y(n_143)
);

AOI31xp33_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_127),
.A3(n_122),
.B(n_19),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_18),
.Y(n_145)
);


endmodule