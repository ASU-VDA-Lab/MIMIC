module fake_jpeg_25337_n_170 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_170);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_20),
.Y(n_58)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

CKINVDCx6p67_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_22),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_26),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_25),
.B1(n_19),
.B2(n_17),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_46),
.B1(n_18),
.B2(n_21),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_36),
.B(n_16),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_58),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_19),
.B1(n_17),
.B2(n_27),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_27),
.B(n_15),
.C(n_30),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_21),
.B(n_31),
.C(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_54),
.Y(n_63)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_26),
.C(n_29),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_26),
.C(n_29),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_38),
.B1(n_34),
.B2(n_39),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_45),
.B1(n_73),
.B2(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_58),
.B(n_16),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_64),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_65),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_74),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_15),
.B1(n_30),
.B2(n_22),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_20),
.B1(n_2),
.B2(n_3),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_23),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_72),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_23),
.Y(n_72)
);

AO21x1_ASAP7_75t_SL g89 ( 
.A1(n_73),
.A2(n_1),
.B(n_4),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_50),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_41),
.C(n_29),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_76),
.B1(n_45),
.B2(n_47),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_41),
.B(n_20),
.C(n_40),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_68),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_81),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_48),
.B1(n_45),
.B2(n_55),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_80),
.A2(n_90),
.B1(n_71),
.B2(n_51),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_31),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_74),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_84),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_64),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_50),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_89),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_88),
.A2(n_56),
.B1(n_47),
.B2(n_5),
.Y(n_110)
);

OAI32xp33_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_51),
.A3(n_45),
.B1(n_5),
.B2(n_7),
.Y(n_92)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_66),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_94),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_66),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_62),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_104),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_76),
.B(n_59),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_108),
.B(n_109),
.Y(n_124)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

NOR3xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_75),
.C(n_59),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_107),
.Y(n_113)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_71),
.B1(n_51),
.B2(n_56),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_86),
.B1(n_92),
.B2(n_79),
.Y(n_123)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_112),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_102),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_77),
.Y(n_114)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_85),
.Y(n_115)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_116),
.C(n_118),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_85),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_91),
.C(n_82),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_104),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_120),
.Y(n_135)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_97),
.B(n_82),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_122),
.A2(n_123),
.B(n_101),
.Y(n_126)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_129),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_126),
.A2(n_130),
.B(n_131),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_124),
.A2(n_103),
.B(n_96),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_127),
.B(n_134),
.Y(n_139)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_SL g130 ( 
.A(n_123),
.B(n_101),
.C(n_100),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_96),
.B(n_99),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_110),
.B1(n_91),
.B2(n_79),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_59),
.B1(n_56),
.B2(n_8),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_1),
.B(n_4),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_118),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_140),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_115),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_133),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_142),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_116),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_136),
.B(n_117),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_145),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_47),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_146),
.A2(n_135),
.B(n_132),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_R g147 ( 
.A(n_139),
.B(n_130),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_153),
.B(n_148),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_149),
.A2(n_142),
.B1(n_7),
.B2(n_8),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_144),
.B(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_151),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_132),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_148),
.B(n_137),
.Y(n_154)
);

FAx1_ASAP7_75t_SL g160 ( 
.A(n_154),
.B(n_9),
.CI(n_10),
.CON(n_160),
.SN(n_160)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_138),
.C(n_11),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_157),
.B(n_158),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_140),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_59),
.Y(n_161)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_160),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_162),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_9),
.C(n_10),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_163),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_166),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_160),
.C(n_13),
.Y(n_168)
);

OAI22x1_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_164),
.B1(n_4),
.B2(n_7),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_167),
.Y(n_170)
);


endmodule