module fake_ariane_1750_n_108 (n_8, n_3, n_2, n_11, n_7, n_16, n_5, n_14, n_1, n_0, n_12, n_15, n_6, n_13, n_9, n_17, n_4, n_10, n_108);

input n_8;
input n_3;
input n_2;
input n_11;
input n_7;
input n_16;
input n_5;
input n_14;
input n_1;
input n_0;
input n_12;
input n_15;
input n_6;
input n_13;
input n_9;
input n_17;
input n_4;
input n_10;

output n_108;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_18;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_19;
wire n_40;
wire n_106;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_58;
wire n_37;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_102;
wire n_22;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_35;
wire n_54;
wire n_25;

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVxp33_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVxp33_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_22),
.Y(n_37)
);

OAI21x1_ASAP7_75t_L g38 ( 
.A1(n_26),
.A2(n_6),
.B(n_7),
.Y(n_38)
);

AND2x4_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_24),
.Y(n_42)
);

AND2x4_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_2),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_19),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NAND2x1p5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_19),
.Y(n_52)
);

AND2x4_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_20),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_49),
.B(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_53),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_57),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_58),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_43),
.B1(n_39),
.B2(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

OA21x2_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_38),
.B(n_56),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_43),
.B(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_39),
.B1(n_51),
.B2(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_37),
.B1(n_61),
.B2(n_47),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_68),
.B1(n_52),
.B2(n_44),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_74),
.A2(n_58),
.B1(n_40),
.B2(n_54),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_75),
.B(n_77),
.Y(n_79)
);

AND2x4_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_72),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_71),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_33),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_4),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_4),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

AOI222xp33_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_71),
.B1(n_35),
.B2(n_82),
.C1(n_79),
.C2(n_56),
.Y(n_89)
);

NOR4xp25_ASAP7_75t_SL g90 ( 
.A(n_86),
.B(n_83),
.C(n_66),
.D(n_35),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_35),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_12),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_92),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_88),
.Y(n_95)
);

OAI31xp33_ASAP7_75t_L g96 ( 
.A1(n_94),
.A2(n_84),
.A3(n_86),
.B(n_89),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

AOI222xp33_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_54),
.B1(n_90),
.B2(n_55),
.C1(n_58),
.C2(n_66),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_96),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_98),
.A2(n_66),
.B1(n_16),
.B2(n_13),
.Y(n_101)
);

CKINVDCx5p33_ASAP7_75t_R g102 ( 
.A(n_100),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g103 ( 
.A(n_101),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_54),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_102),
.B(n_55),
.Y(n_108)
);


endmodule