module real_jpeg_18457_n_4 (n_0, n_1, n_2, n_30, n_28, n_29, n_3, n_4);

input n_0;
input n_1;
input n_2;
input n_30;
input n_28;
input n_29;
input n_3;

output n_4;

wire n_17;
wire n_8;
wire n_21;
wire n_10;
wire n_9;
wire n_12;
wire n_24;
wire n_6;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_5;
wire n_26;
wire n_20;
wire n_19;
wire n_16;
wire n_15;
wire n_13;

AND2x2_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_17),
.Y(n_16)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g5 ( 
.A1(n_2),
.A2(n_6),
.B1(n_7),
.B2(n_12),
.Y(n_5)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g4 ( 
.A(n_5),
.B(n_13),
.Y(n_4)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g7 ( 
.A(n_8),
.B(n_11),
.Y(n_7)
);

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_9),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_20),
.C(n_21),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_19),
.Y(n_17)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2x1_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g11 ( 
.A(n_28),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_29),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_30),
.Y(n_23)
);


endmodule