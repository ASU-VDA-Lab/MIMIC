module fake_jpeg_3150_n_203 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_203);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_7),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_10),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

BUFx12f_ASAP7_75t_SL g70 ( 
.A(n_63),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_74),
.Y(n_86)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_68),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_71),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_53),
.Y(n_93)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_70),
.A2(n_66),
.B1(n_52),
.B2(n_63),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_84),
.A2(n_87),
.B1(n_47),
.B2(n_67),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_52),
.B(n_53),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_76),
.A2(n_66),
.B1(n_52),
.B2(n_53),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_51),
.Y(n_92)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_99),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_94),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_46),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_82),
.B(n_55),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_96),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_62),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_49),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_102),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_103),
.B1(n_59),
.B2(n_57),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_49),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_79),
.A2(n_58),
.B1(n_60),
.B2(n_54),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_67),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_107),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_47),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_59),
.C(n_57),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_1),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_78),
.A2(n_61),
.B1(n_64),
.B2(n_59),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_108),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_90),
.B1(n_81),
.B2(n_77),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_114),
.B1(n_126),
.B2(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_100),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_116),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_91),
.A2(n_77),
.B1(n_81),
.B2(n_61),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

BUFx4f_ASAP7_75t_SL g149 ( 
.A(n_119),
.Y(n_149)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_12),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_57),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_31),
.Y(n_144)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_91),
.A2(n_64),
.B1(n_4),
.B2(n_5),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_99),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_9),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_121),
.A2(n_108),
.B1(n_105),
.B2(n_95),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_132),
.A2(n_134),
.B1(n_145),
.B2(n_153),
.Y(n_157)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_135),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_117),
.A2(n_113),
.B1(n_129),
.B2(n_124),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_127),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_115),
.B(n_6),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_141),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_105),
.B(n_97),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_33),
.B(n_40),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_147),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_122),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_11),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

NOR2x1_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_13),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_154),
.Y(n_165)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_125),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_15),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_146),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_155),
.A2(n_145),
.B1(n_153),
.B2(n_143),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_36),
.C(n_43),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_164),
.C(n_167),
.Y(n_177)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_142),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_170),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_34),
.C(n_41),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_169),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_44),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

A2O1A1O1Ixp25_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_32),
.B(n_38),
.C(n_21),
.D(n_23),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

XNOR2x2_ASAP7_75t_SL g171 ( 
.A(n_148),
.B(n_17),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_149),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_132),
.B(n_150),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_174),
.B(n_179),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_161),
.A2(n_149),
.B1(n_138),
.B2(n_19),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_180),
.A2(n_183),
.B1(n_161),
.B2(n_171),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_149),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_184),
.B(n_186),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_167),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_177),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_178),
.A2(n_159),
.B1(n_170),
.B2(n_160),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_175),
.A2(n_165),
.B1(n_157),
.B2(n_172),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_190),
.C(n_176),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_182),
.A2(n_164),
.B1(n_169),
.B2(n_30),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_192),
.B(n_26),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_194),
.Y(n_196)
);

XNOR2x1_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_177),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_191),
.A2(n_188),
.B1(n_187),
.B2(n_186),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_191),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_27),
.C(n_37),
.Y(n_199)
);

BUFx24_ASAP7_75t_SL g200 ( 
.A(n_198),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_200),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_201),
.A2(n_195),
.B1(n_196),
.B2(n_199),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_196),
.Y(n_203)
);


endmodule