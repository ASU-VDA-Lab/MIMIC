module fake_netlist_6_2714_n_171 (n_41, n_16, n_1, n_34, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_27, n_3, n_14, n_38, n_0, n_39, n_32, n_4, n_36, n_22, n_26, n_13, n_35, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_40, n_171);

input n_41;
input n_16;
input n_1;
input n_34;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_27;
input n_3;
input n_14;
input n_38;
input n_0;
input n_39;
input n_32;
input n_4;
input n_36;
input n_22;
input n_26;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;
input n_40;

output n_171;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_163;
wire n_146;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_127;
wire n_125;
wire n_168;
wire n_153;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_140;
wire n_70;
wire n_120;
wire n_67;
wire n_82;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_48;
wire n_65;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_134;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx2_ASAP7_75t_SL g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

INVxp33_ASAP7_75t_SL g47 ( 
.A(n_26),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

INVxp33_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

INVxp33_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_32),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_12),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_62),
.Y(n_74)
);

AOI21x1_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_18),
.B(n_36),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_0),
.Y(n_78)
);

OR2x6_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_0),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_8),
.B1(n_9),
.B2(n_13),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_17),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_19),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_43),
.B(n_23),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_45),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_81),
.B(n_53),
.Y(n_93)
);

CKINVDCx5p33_ASAP7_75t_R g94 ( 
.A(n_90),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_76),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_50),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_84),
.B(n_69),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_44),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_65),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_101),
.B(n_78),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_87),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_84),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_85),
.B(n_82),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

AND2x4_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_79),
.Y(n_120)
);

OAI21x1_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_75),
.B(n_47),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_93),
.B(n_56),
.Y(n_123)
);

NAND2x1p5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_96),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_92),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_100),
.B(n_79),
.Y(n_126)
);

O2A1O1Ixp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_79),
.B(n_94),
.C(n_100),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_120),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_94),
.Y(n_129)
);

AOI221xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_54),
.B1(n_51),
.B2(n_48),
.C(n_46),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_27),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_29),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_40),
.Y(n_135)
);

INVxp67_ASAP7_75t_SL g136 ( 
.A(n_124),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_119),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_125),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_118),
.B1(n_114),
.B2(n_117),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_119),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_113),
.Y(n_145)
);

AND2x4_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_109),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_145),
.A2(n_134),
.B(n_126),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_141),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

AOI21x1_ASAP7_75t_L g153 ( 
.A1(n_147),
.A2(n_121),
.B(n_109),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_130),
.B1(n_142),
.B2(n_144),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_152),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_143),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_157),
.B(n_155),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_156),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_158),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_149),
.B(n_136),
.Y(n_162)
);

OAI211xp5_ASAP7_75t_SL g163 ( 
.A1(n_160),
.A2(n_126),
.B(n_150),
.C(n_148),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_161),
.A2(n_136),
.B(n_142),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_165),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_162),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_164),
.B1(n_143),
.B2(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_168),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_137),
.B(n_153),
.Y(n_170)
);

AOI221xp5_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_33),
.B1(n_35),
.B2(n_146),
.C(n_169),
.Y(n_171)
);


endmodule