module fake_jpeg_17459_n_117 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_117);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_117;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_51),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_52),
.B(n_47),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_55),
.A2(n_43),
.B1(n_45),
.B2(n_48),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_55),
.B(n_49),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_62),
.B1(n_64),
.B2(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_53),
.B(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_63),
.Y(n_79)
);

NOR2x1_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_42),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_50),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_42),
.B1(n_44),
.B2(n_40),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_50),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_72),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_36),
.B1(n_41),
.B2(n_39),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_88)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_75),
.Y(n_91)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_92)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_77),
.Y(n_85)
);

AO22x1_ASAP7_75t_SL g78 ( 
.A1(n_64),
.A2(n_45),
.B1(n_42),
.B2(n_23),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_78),
.A2(n_81),
.B1(n_60),
.B2(n_79),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_38),
.C(n_21),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_0),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_84),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_70),
.Y(n_87)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_90),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_1),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

AOI32xp33_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_81),
.A3(n_78),
.B1(n_73),
.B2(n_8),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_93),
.A2(n_95),
.B(n_89),
.Y(n_99)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_26),
.C(n_35),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_103),
.B(n_5),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_97),
.B(n_94),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_82),
.C(n_85),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_101),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_96),
.B(n_91),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_102),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_95),
.A2(n_92),
.B1(n_71),
.B2(n_7),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_6),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_104),
.C(n_107),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

AOI31xp67_ASAP7_75t_SL g111 ( 
.A1(n_110),
.A2(n_109),
.A3(n_7),
.B(n_13),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_11),
.B(n_15),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_16),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_17),
.B1(n_22),
.B2(n_24),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_114),
.A2(n_25),
.B(n_27),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_115),
.A2(n_33),
.B(n_29),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_28),
.Y(n_117)
);


endmodule