module real_aes_10365_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_769;
wire n_434;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_1343;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_269;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1352;
wire n_1280;
wire n_1323;
wire n_1097;
wire n_1369;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVxp33_ASAP7_75t_L g1335 ( .A(n_0), .Y(n_1335) );
AOI22xp33_ASAP7_75t_L g1359 ( .A1(n_0), .A2(n_248), .B1(n_486), .B2(n_1360), .Y(n_1359) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_1), .A2(n_191), .B1(n_1081), .B2(n_1083), .Y(n_1080) );
AOI22xp33_ASAP7_75t_SL g1114 ( .A1(n_1), .A2(n_4), .B1(n_580), .B2(n_1115), .Y(n_1114) );
AO221x1_ASAP7_75t_L g1179 ( .A1(n_2), .A2(n_136), .B1(n_1150), .B2(n_1180), .C(n_1181), .Y(n_1179) );
OAI221xp5_ASAP7_75t_L g549 ( .A1(n_3), .A2(n_550), .B1(n_553), .B2(n_561), .C(n_564), .Y(n_549) );
AOI21xp33_ASAP7_75t_L g616 ( .A1(n_3), .A2(n_617), .B(n_619), .Y(n_616) );
AOI221xp5_ASAP7_75t_L g1079 ( .A1(n_4), .A2(n_157), .B1(n_286), .B2(n_763), .C(n_1036), .Y(n_1079) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_5), .Y(n_261) );
AND2x2_ASAP7_75t_L g351 ( .A(n_5), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g406 ( .A(n_5), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_5), .B(n_179), .Y(n_413) );
INVx1_ASAP7_75t_L g388 ( .A(n_6), .Y(n_388) );
INVxp67_ASAP7_75t_L g807 ( .A(n_7), .Y(n_807) );
OAI222xp33_ASAP7_75t_L g822 ( .A1(n_7), .A2(n_36), .B1(n_234), .B2(n_313), .C1(n_464), .C2(n_543), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g1171 ( .A1(n_8), .A2(n_97), .B1(n_1126), .B2(n_1150), .Y(n_1171) );
INVxp67_ASAP7_75t_L g1342 ( .A(n_9), .Y(n_1342) );
AOI22xp33_ASAP7_75t_L g1366 ( .A1(n_9), .A2(n_65), .B1(n_486), .B2(n_1067), .Y(n_1366) );
INVx1_ASAP7_75t_L g397 ( .A(n_10), .Y(n_397) );
XNOR2x2_ASAP7_75t_L g1008 ( .A(n_11), .B(n_1009), .Y(n_1008) );
AOI221xp5_ASAP7_75t_L g974 ( .A1(n_12), .A2(n_159), .B1(n_486), .B2(n_975), .C(n_976), .Y(n_974) );
INVx1_ASAP7_75t_L g994 ( .A(n_12), .Y(n_994) );
OAI221xp5_ASAP7_75t_L g569 ( .A1(n_13), .A2(n_20), .B1(n_570), .B2(n_573), .C(n_574), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g627 ( .A(n_13), .Y(n_627) );
AO22x2_ASAP7_75t_L g713 ( .A1(n_14), .A2(n_714), .B1(n_781), .B2(n_782), .Y(n_713) );
CKINVDCx14_ASAP7_75t_R g781 ( .A(n_14), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_15), .A2(n_72), .B1(n_652), .B2(n_861), .Y(n_860) );
OAI22xp5_ASAP7_75t_L g894 ( .A1(n_15), .A2(n_27), .B1(n_350), .B2(n_411), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_16), .A2(n_222), .B1(n_652), .B2(n_831), .Y(n_983) );
INVx1_ASAP7_75t_L g1003 ( .A(n_16), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_17), .A2(n_33), .B1(n_486), .B2(n_1071), .Y(n_1070) );
INVxp33_ASAP7_75t_SL g1104 ( .A(n_17), .Y(n_1104) );
AOI221xp5_ASAP7_75t_L g1382 ( .A1(n_18), .A2(n_233), .B1(n_647), .B2(n_838), .C(n_839), .Y(n_1382) );
INVx1_ASAP7_75t_L g1402 ( .A(n_18), .Y(n_1402) );
AO221x2_ASAP7_75t_L g1201 ( .A1(n_19), .A2(n_158), .B1(n_1180), .B2(n_1202), .C(n_1204), .Y(n_1201) );
CKINVDCx5p33_ASAP7_75t_R g626 ( .A(n_20), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g886 ( .A1(n_21), .A2(n_129), .B1(n_402), .B2(n_887), .C(n_888), .Y(n_886) );
OAI22xp5_ASAP7_75t_L g897 ( .A1(n_21), .A2(n_205), .B1(n_451), .B2(n_538), .Y(n_897) );
INVx2_ASAP7_75t_L g282 ( .A(n_22), .Y(n_282) );
OR2x2_ASAP7_75t_L g441 ( .A(n_22), .B(n_330), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_23), .A2(n_216), .B1(n_665), .B2(n_667), .Y(n_664) );
OAI221xp5_ASAP7_75t_L g685 ( .A1(n_23), .A2(n_216), .B1(n_686), .B2(n_688), .C(n_689), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_24), .A2(n_52), .B1(n_747), .B2(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g880 ( .A(n_24), .Y(n_880) );
INVx1_ASAP7_75t_L g808 ( .A(n_25), .Y(n_808) );
OAI221xp5_ASAP7_75t_L g920 ( .A1(n_26), .A2(n_87), .B1(n_686), .B2(n_688), .C(n_921), .Y(n_920) );
OAI22xp5_ASAP7_75t_L g948 ( .A1(n_26), .A2(n_87), .B1(n_667), .B2(n_818), .Y(n_948) );
OAI222xp33_ASAP7_75t_L g896 ( .A1(n_27), .A2(n_129), .B1(n_135), .B2(n_540), .C1(n_542), .C2(n_674), .Y(n_896) );
BUFx2_ASAP7_75t_L g284 ( .A(n_28), .Y(n_284) );
BUFx2_ASAP7_75t_L g318 ( .A(n_28), .Y(n_318) );
INVx1_ASAP7_75t_L g332 ( .A(n_28), .Y(n_332) );
OR2x2_ASAP7_75t_L g572 ( .A(n_28), .B(n_413), .Y(n_572) );
INVx1_ASAP7_75t_L g717 ( .A(n_29), .Y(n_717) );
AOI21xp33_ASAP7_75t_L g762 ( .A1(n_29), .A2(n_485), .B(n_763), .Y(n_762) );
AOI22xp33_ASAP7_75t_SL g560 ( .A1(n_30), .A2(n_139), .B1(n_414), .B2(n_506), .Y(n_560) );
INVx1_ASAP7_75t_L g607 ( .A(n_30), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g733 ( .A(n_31), .Y(n_733) );
INVx1_ASAP7_75t_L g471 ( .A(n_32), .Y(n_471) );
INVxp33_ASAP7_75t_SL g1099 ( .A(n_33), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_34), .A2(n_75), .B1(n_432), .B2(n_566), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_34), .A2(n_75), .B1(n_590), .B2(n_593), .Y(n_589) );
INVx1_ASAP7_75t_L g795 ( .A(n_35), .Y(n_795) );
INVxp67_ASAP7_75t_L g805 ( .A(n_36), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_37), .A2(n_184), .B1(n_652), .B2(n_654), .Y(n_651) );
INVx1_ASAP7_75t_L g692 ( .A(n_37), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g764 ( .A1(n_38), .A2(n_199), .B1(n_765), .B2(n_767), .C(n_769), .Y(n_764) );
INVx1_ASAP7_75t_L g774 ( .A(n_38), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_39), .A2(n_43), .B1(n_499), .B2(n_1014), .Y(n_1013) );
OAI22xp5_ASAP7_75t_L g1057 ( .A1(n_39), .A2(n_56), .B1(n_451), .B2(n_538), .Y(n_1057) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_40), .Y(n_333) );
INVx1_ASAP7_75t_L g868 ( .A(n_41), .Y(n_868) );
OAI221xp5_ASAP7_75t_L g890 ( .A1(n_41), .A2(n_73), .B1(n_514), .B2(n_891), .C(n_893), .Y(n_890) );
INVx1_ASAP7_75t_L g1182 ( .A(n_42), .Y(n_1182) );
INVxp67_ASAP7_75t_SL g1055 ( .A(n_43), .Y(n_1055) );
INVx1_ASAP7_75t_L g556 ( .A(n_44), .Y(n_556) );
AOI21xp33_ASAP7_75t_L g603 ( .A1(n_44), .A2(n_604), .B(n_605), .Y(n_603) );
INVx1_ASAP7_75t_L g1028 ( .A(n_45), .Y(n_1028) );
CKINVDCx5p33_ASAP7_75t_R g978 ( .A(n_46), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_47), .A2(n_173), .B1(n_473), .B2(n_475), .Y(n_472) );
INVxp67_ASAP7_75t_SL g525 ( .A(n_47), .Y(n_525) );
INVx1_ASAP7_75t_L g940 ( .A(n_48), .Y(n_940) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_49), .Y(n_533) );
AOI221xp5_ASAP7_75t_L g646 ( .A1(n_50), .A2(n_58), .B1(n_604), .B2(n_647), .C(n_649), .Y(n_646) );
INVxp67_ASAP7_75t_SL g695 ( .A(n_50), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_51), .A2(n_177), .B1(n_311), .B2(n_312), .Y(n_310) );
OAI22xp33_ASAP7_75t_L g346 ( .A1(n_51), .A2(n_244), .B1(n_347), .B2(n_357), .Y(n_346) );
INVx1_ASAP7_75t_L g878 ( .A(n_52), .Y(n_878) );
AO221x1_ASAP7_75t_L g1154 ( .A1(n_53), .A2(n_68), .B1(n_1126), .B2(n_1150), .C(n_1155), .Y(n_1154) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_54), .Y(n_340) );
INVx1_ASAP7_75t_L g1183 ( .A(n_55), .Y(n_1183) );
AOI221xp5_ASAP7_75t_L g1016 ( .A1(n_56), .A2(n_169), .B1(n_402), .B2(n_1017), .C(n_1019), .Y(n_1016) );
INVxp33_ASAP7_75t_SL g926 ( .A(n_57), .Y(n_926) );
AOI221xp5_ASAP7_75t_L g954 ( .A1(n_57), .A2(n_83), .B1(n_955), .B2(n_956), .C(n_958), .Y(n_954) );
INVxp67_ASAP7_75t_SL g697 ( .A(n_58), .Y(n_697) );
INVxp67_ASAP7_75t_L g1340 ( .A(n_59), .Y(n_1340) );
AOI221xp5_ASAP7_75t_L g1363 ( .A1(n_59), .A2(n_160), .B1(n_649), .B2(n_1364), .C(n_1365), .Y(n_1363) );
INVxp33_ASAP7_75t_SL g1092 ( .A(n_60), .Y(n_1092) );
AOI22xp33_ASAP7_75t_SL g1118 ( .A1(n_60), .A2(n_96), .B1(n_1112), .B2(n_1119), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g1383 ( .A1(n_61), .A2(n_214), .B1(n_474), .B2(n_486), .Y(n_1383) );
INVx1_ASAP7_75t_L g1403 ( .A(n_61), .Y(n_1403) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_62), .Y(n_559) );
AO221x1_ASAP7_75t_L g1160 ( .A1(n_63), .A2(n_103), .B1(n_1126), .B2(n_1150), .C(n_1161), .Y(n_1160) );
INVx1_ASAP7_75t_L g1207 ( .A(n_64), .Y(n_1207) );
INVxp67_ASAP7_75t_L g1344 ( .A(n_65), .Y(n_1344) );
INVxp33_ASAP7_75t_L g912 ( .A(n_66), .Y(n_912) );
AOI221xp5_ASAP7_75t_L g949 ( .A1(n_66), .A2(n_246), .B1(n_486), .B2(n_950), .C(n_951), .Y(n_949) );
AOI221xp5_ASAP7_75t_L g835 ( .A1(n_67), .A2(n_124), .B1(n_836), .B2(n_838), .C(n_839), .Y(n_835) );
OAI221xp5_ASAP7_75t_L g842 ( .A1(n_67), .A2(n_144), .B1(n_843), .B2(n_844), .C(n_847), .Y(n_842) );
INVx1_ASAP7_75t_L g1158 ( .A(n_69), .Y(n_1158) );
INVx1_ASAP7_75t_L g281 ( .A(n_70), .Y(n_281) );
INVx1_ASAP7_75t_L g330 ( .A(n_70), .Y(n_330) );
INVx1_ASAP7_75t_L g641 ( .A(n_71), .Y(n_641) );
INVx1_ASAP7_75t_L g889 ( .A(n_72), .Y(n_889) );
INVx1_ASAP7_75t_L g867 ( .A(n_73), .Y(n_867) );
INVxp33_ASAP7_75t_L g1093 ( .A(n_74), .Y(n_1093) );
AOI22xp33_ASAP7_75t_SL g1116 ( .A1(n_74), .A2(n_186), .B1(n_580), .B2(n_1117), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_76), .A2(n_114), .B1(n_484), .B2(n_486), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_76), .A2(n_114), .B1(n_347), .B2(n_430), .Y(n_529) );
OAI221xp5_ASAP7_75t_L g1336 ( .A1(n_77), .A2(n_106), .B1(n_790), .B2(n_921), .C(n_1337), .Y(n_1336) );
OAI22xp5_ASAP7_75t_L g1361 ( .A1(n_77), .A2(n_106), .B1(n_667), .B2(n_765), .Y(n_1361) );
OAI22xp33_ASAP7_75t_L g584 ( .A1(n_78), .A2(n_130), .B1(n_585), .B2(n_587), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_78), .A2(n_189), .B1(n_288), .B2(n_611), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g1074 ( .A1(n_79), .A2(n_225), .B1(n_1075), .B2(n_1076), .Y(n_1074) );
INVxp67_ASAP7_75t_SL g1096 ( .A(n_79), .Y(n_1096) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_80), .A2(n_189), .B1(n_578), .B2(n_581), .Y(n_577) );
INVx1_ASAP7_75t_L g613 ( .A(n_80), .Y(n_613) );
XNOR2xp5_ASAP7_75t_L g785 ( .A(n_81), .B(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g1030 ( .A(n_82), .Y(n_1030) );
AOI221xp5_ASAP7_75t_L g1035 ( .A1(n_82), .A2(n_239), .B1(n_1036), .B2(n_1038), .C(n_1039), .Y(n_1035) );
INVxp67_ASAP7_75t_SL g929 ( .A(n_83), .Y(n_929) );
CKINVDCx5p33_ASAP7_75t_R g1393 ( .A(n_84), .Y(n_1393) );
INVxp67_ASAP7_75t_L g793 ( .A(n_85), .Y(n_793) );
AOI221xp5_ASAP7_75t_L g825 ( .A1(n_85), .A2(n_142), .B1(n_604), .B2(n_649), .C(n_749), .Y(n_825) );
AOI22xp33_ASAP7_75t_SL g858 ( .A1(n_86), .A2(n_105), .B1(n_838), .B2(n_859), .Y(n_858) );
AOI21xp33_ASAP7_75t_L g876 ( .A1(n_86), .A2(n_414), .B(n_562), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g1176 ( .A1(n_88), .A2(n_198), .B1(n_1126), .B2(n_1150), .Y(n_1176) );
AOI221xp5_ASAP7_75t_L g1388 ( .A1(n_89), .A2(n_203), .B1(n_605), .B2(n_647), .C(n_955), .Y(n_1388) );
INVx1_ASAP7_75t_L g1412 ( .A(n_89), .Y(n_1412) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_90), .A2(n_209), .B1(n_661), .B2(n_662), .Y(n_660) );
INVx1_ASAP7_75t_L g684 ( .A(n_90), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_91), .A2(n_190), .B1(n_299), .B2(n_647), .C(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g681 ( .A(n_91), .Y(n_681) );
OAI22xp33_ASAP7_75t_L g489 ( .A1(n_92), .A2(n_215), .B1(n_323), .B2(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g512 ( .A(n_92), .Y(n_512) );
INVx1_ASAP7_75t_L g1163 ( .A(n_93), .Y(n_1163) );
INVx1_ASAP7_75t_L g253 ( .A(n_94), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g985 ( .A(n_95), .Y(n_985) );
INVxp67_ASAP7_75t_SL g1087 ( .A(n_96), .Y(n_1087) );
CKINVDCx5p33_ASAP7_75t_R g1395 ( .A(n_98), .Y(n_1395) );
XOR2x2_ASAP7_75t_L g458 ( .A(n_99), .B(n_459), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g1139 ( .A1(n_99), .A2(n_181), .B1(n_1140), .B2(n_1146), .Y(n_1139) );
INVx1_ASAP7_75t_L g480 ( .A(n_100), .Y(n_480) );
OAI221xp5_ASAP7_75t_L g515 ( .A1(n_100), .A2(n_427), .B1(n_516), .B2(n_522), .C(n_527), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g730 ( .A(n_101), .Y(n_730) );
CKINVDCx5p33_ASAP7_75t_R g1063 ( .A(n_102), .Y(n_1063) );
AOI222xp33_ASAP7_75t_L g1324 ( .A1(n_103), .A2(n_1325), .B1(n_1369), .B2(n_1373), .C1(n_1420), .C2(n_1424), .Y(n_1324) );
XNOR2x1_ASAP7_75t_L g1326 ( .A(n_103), .B(n_1327), .Y(n_1326) );
INVx1_ASAP7_75t_L g1162 ( .A(n_104), .Y(n_1162) );
INVx1_ASAP7_75t_L g875 ( .A(n_105), .Y(n_875) );
INVx1_ASAP7_75t_L g1348 ( .A(n_107), .Y(n_1348) );
XOR2xp5_ASAP7_75t_L g546 ( .A(n_108), .B(n_547), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g1149 ( .A1(n_109), .A2(n_163), .B1(n_1126), .B2(n_1150), .Y(n_1149) );
AOI22xp5_ASAP7_75t_L g1177 ( .A1(n_110), .A2(n_247), .B1(n_1140), .B2(n_1146), .Y(n_1177) );
AOI221xp5_ASAP7_75t_L g503 ( .A1(n_111), .A2(n_170), .B1(n_504), .B2(n_505), .C(n_507), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_111), .A2(n_151), .B1(n_451), .B2(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g941 ( .A(n_112), .Y(n_941) );
OAI222xp33_ASAP7_75t_L g788 ( .A1(n_113), .A2(n_143), .B1(n_238), .B2(n_587), .C1(n_789), .C2(n_790), .Y(n_788) );
INVx1_ASAP7_75t_L g816 ( .A(n_113), .Y(n_816) );
INVx1_ASAP7_75t_L g1033 ( .A(n_115), .Y(n_1033) );
INVx1_ASAP7_75t_L g497 ( .A(n_116), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_116), .A2(n_170), .B1(n_540), .B2(n_542), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g736 ( .A(n_117), .Y(n_736) );
INVx1_ASAP7_75t_L g1205 ( .A(n_118), .Y(n_1205) );
XNOR2xp5_ASAP7_75t_L g849 ( .A(n_119), .B(n_850), .Y(n_849) );
CKINVDCx5p33_ASAP7_75t_R g1394 ( .A(n_120), .Y(n_1394) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_121), .A2(n_229), .B1(n_286), .B2(n_291), .Y(n_285) );
INVx1_ASAP7_75t_L g370 ( .A(n_121), .Y(n_370) );
INVx1_ASAP7_75t_L g934 ( .A(n_122), .Y(n_934) );
AOI221xp5_ASAP7_75t_L g981 ( .A1(n_123), .A2(n_241), .B1(n_604), .B2(n_958), .C(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g1002 ( .A(n_123), .Y(n_1002) );
OAI332xp33_ASAP7_75t_L g791 ( .A1(n_124), .A2(n_561), .A3(n_707), .B1(n_741), .B2(n_792), .B3(n_797), .C1(n_800), .C2(n_806), .Y(n_791) );
INVx1_ASAP7_75t_L g720 ( .A(n_125), .Y(n_720) );
AOI22xp33_ASAP7_75t_SL g760 ( .A1(n_125), .A2(n_174), .B1(n_487), .B2(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g1353 ( .A(n_126), .Y(n_1353) );
CKINVDCx5p33_ASAP7_75t_R g971 ( .A(n_127), .Y(n_971) );
OAI22xp5_ASAP7_75t_L g1021 ( .A1(n_128), .A2(n_153), .B1(n_514), .B2(n_891), .Y(n_1021) );
OAI221xp5_ASAP7_75t_L g1049 ( .A1(n_128), .A2(n_153), .B1(n_1050), .B2(n_1052), .C(n_1053), .Y(n_1049) );
INVx1_ASAP7_75t_L g621 ( .A(n_130), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g1374 ( .A1(n_131), .A2(n_1375), .B1(n_1376), .B2(n_1419), .Y(n_1374) );
CKINVDCx5p33_ASAP7_75t_R g1375 ( .A(n_131), .Y(n_1375) );
INVx1_ASAP7_75t_L g645 ( .A(n_132), .Y(n_645) );
XNOR2xp5_ASAP7_75t_L g966 ( .A(n_133), .B(n_967), .Y(n_966) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_134), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_135), .A2(n_205), .B1(n_884), .B2(n_885), .Y(n_883) );
AOI22xp33_ASAP7_75t_SL g862 ( .A1(n_137), .A2(n_148), .B1(n_292), .B2(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g871 ( .A(n_137), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_138), .A2(n_244), .B1(n_298), .B2(n_304), .Y(n_309) );
OAI22xp33_ASAP7_75t_L g426 ( .A1(n_138), .A2(n_177), .B1(n_427), .B2(n_430), .Y(n_426) );
INVx1_ASAP7_75t_L g602 ( .A(n_139), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_140), .A2(n_168), .B1(n_740), .B2(n_741), .Y(n_739) );
INVx1_ASAP7_75t_L g753 ( .A(n_140), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_141), .A2(n_196), .B1(n_585), .B2(n_587), .Y(n_742) );
AOI22xp33_ASAP7_75t_SL g756 ( .A1(n_141), .A2(n_168), .B1(n_485), .B2(n_487), .Y(n_756) );
INVx1_ASAP7_75t_L g798 ( .A(n_142), .Y(n_798) );
INVx1_ASAP7_75t_L g829 ( .A(n_143), .Y(n_829) );
INVx1_ASAP7_75t_L g834 ( .A(n_144), .Y(n_834) );
CKINVDCx5p33_ASAP7_75t_R g731 ( .A(n_145), .Y(n_731) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_146), .Y(n_255) );
AND3x2_ASAP7_75t_L g1129 ( .A(n_146), .B(n_253), .C(n_1130), .Y(n_1129) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_146), .B(n_253), .Y(n_1145) );
OA332x1_ASAP7_75t_L g715 ( .A1(n_147), .A2(n_550), .A3(n_561), .B1(n_716), .B2(n_723), .B3(n_729), .C1(n_732), .C2(n_737), .Y(n_715) );
AOI21xp5_ASAP7_75t_L g757 ( .A1(n_147), .A2(n_659), .B(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g872 ( .A(n_148), .Y(n_872) );
INVxp33_ASAP7_75t_L g924 ( .A(n_149), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_149), .A2(n_175), .B1(n_960), .B2(n_961), .Y(n_959) );
INVx1_ASAP7_75t_L g963 ( .A(n_150), .Y(n_963) );
INVx1_ASAP7_75t_L g502 ( .A(n_151), .Y(n_502) );
OAI22xp33_ASAP7_75t_SL g972 ( .A1(n_152), .A2(n_164), .B1(n_818), .B2(n_973), .Y(n_972) );
OAI221xp5_ASAP7_75t_L g996 ( .A1(n_152), .A2(n_164), .B1(n_686), .B2(n_688), .C(n_921), .Y(n_996) );
INVx2_ASAP7_75t_L g266 ( .A(n_154), .Y(n_266) );
INVx1_ASAP7_75t_L g671 ( .A(n_155), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g1066 ( .A1(n_156), .A2(n_220), .B1(n_304), .B2(n_1067), .C(n_1068), .Y(n_1066) );
INVxp33_ASAP7_75t_SL g1101 ( .A(n_156), .Y(n_1101) );
AOI22xp33_ASAP7_75t_SL g1109 ( .A1(n_157), .A2(n_191), .B1(n_1110), .B2(n_1112), .Y(n_1109) );
INVx1_ASAP7_75t_L g991 ( .A(n_159), .Y(n_991) );
INVxp33_ASAP7_75t_L g1346 ( .A(n_160), .Y(n_1346) );
AOI22xp33_ASAP7_75t_L g1389 ( .A1(n_161), .A2(n_224), .B1(n_838), .B2(n_1390), .Y(n_1389) );
INVx1_ASAP7_75t_L g1409 ( .A(n_161), .Y(n_1409) );
CKINVDCx5p33_ASAP7_75t_R g1391 ( .A(n_162), .Y(n_1391) );
INVx1_ASAP7_75t_L g1349 ( .A(n_165), .Y(n_1349) );
INVx1_ASAP7_75t_L g1027 ( .A(n_166), .Y(n_1027) );
INVx1_ASAP7_75t_L g1130 ( .A(n_167), .Y(n_1130) );
INVxp67_ASAP7_75t_SL g1056 ( .A(n_169), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_171), .A2(n_237), .B1(n_414), .B2(n_506), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_171), .A2(n_237), .B1(n_596), .B2(n_597), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_172), .A2(n_218), .B1(n_298), .B2(n_304), .Y(n_297) );
INVx1_ASAP7_75t_L g382 ( .A(n_172), .Y(n_382) );
INVxp67_ASAP7_75t_SL g523 ( .A(n_173), .Y(n_523) );
INVx1_ASAP7_75t_L g724 ( .A(n_174), .Y(n_724) );
INVxp67_ASAP7_75t_SL g931 ( .A(n_175), .Y(n_931) );
OAI211xp5_ASAP7_75t_L g1011 ( .A1(n_176), .A2(n_357), .B(n_1012), .C(n_1022), .Y(n_1011) );
AOI221xp5_ASAP7_75t_L g1041 ( .A1(n_176), .A2(n_183), .B1(n_298), .B2(n_1042), .C(n_1044), .Y(n_1041) );
CKINVDCx20_ASAP7_75t_R g1059 ( .A(n_178), .Y(n_1059) );
INVx1_ASAP7_75t_L g268 ( .A(n_179), .Y(n_268) );
INVx2_ASAP7_75t_L g352 ( .A(n_179), .Y(n_352) );
INVx1_ASAP7_75t_L g1023 ( .A(n_180), .Y(n_1023) );
AOI22xp5_ASAP7_75t_L g1170 ( .A1(n_182), .A2(n_200), .B1(n_1140), .B2(n_1146), .Y(n_1170) );
OAI221xp5_ASAP7_75t_L g1025 ( .A1(n_183), .A2(n_427), .B1(n_527), .B2(n_1026), .C(n_1029), .Y(n_1025) );
INVx1_ASAP7_75t_L g699 ( .A(n_184), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_185), .A2(n_635), .B1(n_710), .B2(n_711), .Y(n_634) );
INVx1_ASAP7_75t_L g711 ( .A(n_185), .Y(n_711) );
INVxp67_ASAP7_75t_SL g1073 ( .A(n_186), .Y(n_1073) );
INVx1_ASAP7_75t_L g938 ( .A(n_187), .Y(n_938) );
INVxp33_ASAP7_75t_L g1334 ( .A(n_188), .Y(n_1334) );
AOI221xp5_ASAP7_75t_L g1358 ( .A1(n_188), .A2(n_192), .B1(n_619), .B2(n_749), .C(n_960), .Y(n_1358) );
INVx1_ASAP7_75t_L g679 ( .A(n_190), .Y(n_679) );
INVxp33_ASAP7_75t_L g1332 ( .A(n_192), .Y(n_1332) );
CKINVDCx5p33_ASAP7_75t_R g980 ( .A(n_193), .Y(n_980) );
INVx1_ASAP7_75t_L g917 ( .A(n_194), .Y(n_917) );
INVx1_ASAP7_75t_L g467 ( .A(n_195), .Y(n_467) );
INVx1_ASAP7_75t_L g770 ( .A(n_196), .Y(n_770) );
INVx1_ASAP7_75t_L g417 ( .A(n_197), .Y(n_417) );
INVx1_ASAP7_75t_L g778 ( .A(n_199), .Y(n_778) );
XOR2xp5_ASAP7_75t_L g273 ( .A(n_200), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g907 ( .A(n_201), .Y(n_907) );
CKINVDCx5p33_ASAP7_75t_R g1384 ( .A(n_202), .Y(n_1384) );
INVx1_ASAP7_75t_L g1410 ( .A(n_203), .Y(n_1410) );
INVx1_ASAP7_75t_L g393 ( .A(n_204), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g986 ( .A(n_206), .Y(n_986) );
OAI22xp5_ASAP7_75t_L g1385 ( .A1(n_207), .A2(n_212), .B1(n_667), .B2(n_1386), .Y(n_1385) );
OAI221xp5_ASAP7_75t_L g1404 ( .A1(n_207), .A2(n_212), .B1(n_688), .B2(n_689), .C(n_1405), .Y(n_1404) );
INVx1_ASAP7_75t_L g1351 ( .A(n_208), .Y(n_1351) );
INVx1_ASAP7_75t_L g678 ( .A(n_209), .Y(n_678) );
INVx1_ASAP7_75t_L g1128 ( .A(n_210), .Y(n_1128) );
NAND2xp5_ASAP7_75t_L g1148 ( .A(n_210), .B(n_1143), .Y(n_1148) );
INVx1_ASAP7_75t_L g819 ( .A(n_211), .Y(n_819) );
INVx1_ASAP7_75t_L g657 ( .A(n_213), .Y(n_657) );
INVx1_ASAP7_75t_L g1399 ( .A(n_214), .Y(n_1399) );
INVx1_ASAP7_75t_L g509 ( .A(n_215), .Y(n_509) );
INVx1_ASAP7_75t_L g799 ( .A(n_217), .Y(n_799) );
INVx1_ASAP7_75t_L g378 ( .A(n_218), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g977 ( .A(n_219), .Y(n_977) );
INVxp33_ASAP7_75t_L g1103 ( .A(n_220), .Y(n_1103) );
CKINVDCx5p33_ASAP7_75t_R g1355 ( .A(n_221), .Y(n_1355) );
INVx1_ASAP7_75t_L g999 ( .A(n_222), .Y(n_999) );
AO22x1_ASAP7_75t_L g1195 ( .A1(n_223), .A2(n_231), .B1(n_1126), .B2(n_1196), .Y(n_1195) );
INVx1_ASAP7_75t_L g1414 ( .A(n_224), .Y(n_1414) );
INVxp67_ASAP7_75t_SL g1097 ( .A(n_225), .Y(n_1097) );
INVx2_ASAP7_75t_L g265 ( .A(n_226), .Y(n_265) );
INVx1_ASAP7_75t_L g482 ( .A(n_227), .Y(n_482) );
OAI211xp5_ASAP7_75t_SL g492 ( .A1(n_227), .A2(n_357), .B(n_493), .C(n_508), .Y(n_492) );
AO22x1_ASAP7_75t_L g1197 ( .A1(n_228), .A2(n_240), .B1(n_1140), .B2(n_1146), .Y(n_1197) );
INVx1_ASAP7_75t_L g364 ( .A(n_229), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g727 ( .A(n_230), .Y(n_727) );
INVx1_ASAP7_75t_L g1024 ( .A(n_232), .Y(n_1024) );
INVx1_ASAP7_75t_L g1400 ( .A(n_233), .Y(n_1400) );
INVxp67_ASAP7_75t_L g801 ( .A(n_234), .Y(n_801) );
INVx1_ASAP7_75t_L g914 ( .A(n_235), .Y(n_914) );
INVx1_ASAP7_75t_L g987 ( .A(n_236), .Y(n_987) );
INVx1_ASAP7_75t_L g820 ( .A(n_238), .Y(n_820) );
AOI21xp33_ASAP7_75t_L g1031 ( .A1(n_239), .A2(n_562), .B(n_1017), .Y(n_1031) );
INVx1_ASAP7_75t_L g1000 ( .A(n_241), .Y(n_1000) );
BUFx3_ASAP7_75t_L g290 ( .A(n_242), .Y(n_290) );
INVx1_ASAP7_75t_L g296 ( .A(n_242), .Y(n_296) );
INVx1_ASAP7_75t_L g289 ( .A(n_243), .Y(n_289) );
BUFx3_ASAP7_75t_L g295 ( .A(n_243), .Y(n_295) );
INVx1_ASAP7_75t_L g639 ( .A(n_245), .Y(n_639) );
INVxp33_ASAP7_75t_L g918 ( .A(n_246), .Y(n_918) );
INVxp33_ASAP7_75t_L g1331 ( .A(n_248), .Y(n_1331) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_269), .B(n_1122), .Y(n_249) );
AND2x4_ASAP7_75t_L g250 ( .A(n_251), .B(n_256), .Y(n_250) );
AND2x4_ASAP7_75t_L g1372 ( .A(n_251), .B(n_257), .Y(n_1372) );
NOR2xp33_ASAP7_75t_SL g251 ( .A(n_252), .B(n_254), .Y(n_251) );
INVx1_ASAP7_75t_SL g1423 ( .A(n_252), .Y(n_1423) );
NAND2xp5_ASAP7_75t_L g1429 ( .A(n_252), .B(n_254), .Y(n_1429) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g1422 ( .A(n_254), .B(n_1423), .Y(n_1422) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_258), .B(n_262), .Y(n_257) );
INVxp67_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g385 ( .A(n_260), .B(n_268), .Y(n_385) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g562 ( .A(n_261), .B(n_563), .Y(n_562) );
OR2x6_ASAP7_75t_L g262 ( .A(n_263), .B(n_267), .Y(n_262) );
BUFx2_ASAP7_75t_L g381 ( .A(n_263), .Y(n_381) );
INVx1_ASAP7_75t_L g399 ( .A(n_263), .Y(n_399) );
INVx2_ASAP7_75t_SL g520 ( .A(n_263), .Y(n_520) );
OR2x2_ASAP7_75t_L g587 ( .A(n_263), .B(n_572), .Y(n_587) );
BUFx6f_ASAP7_75t_L g705 ( .A(n_263), .Y(n_705) );
INVx2_ASAP7_75t_SL g726 ( .A(n_263), .Y(n_726) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
AND2x4_ASAP7_75t_L g355 ( .A(n_265), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g361 ( .A(n_265), .Y(n_361) );
INVx2_ASAP7_75t_L g369 ( .A(n_265), .Y(n_369) );
INVx1_ASAP7_75t_L g377 ( .A(n_265), .Y(n_377) );
AND2x2_ASAP7_75t_L g416 ( .A(n_265), .B(n_266), .Y(n_416) );
INVx2_ASAP7_75t_L g356 ( .A(n_266), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_266), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g376 ( .A(n_266), .Y(n_376) );
INVx1_ASAP7_75t_L g423 ( .A(n_266), .Y(n_423) );
INVx1_ASAP7_75t_L g434 ( .A(n_266), .Y(n_434) );
INVx2_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
XNOR2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_902), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_631), .B1(n_900), .B2(n_901), .Y(n_270) );
INVx1_ASAP7_75t_L g900 ( .A(n_271), .Y(n_900) );
XNOR2x1_ASAP7_75t_SL g271 ( .A(n_272), .B(n_456), .Y(n_271) );
BUFx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND4xp75_ASAP7_75t_L g274 ( .A(n_275), .B(n_345), .C(n_437), .D(n_446), .Y(n_274) );
AND2x2_ASAP7_75t_SL g275 ( .A(n_276), .B(n_321), .Y(n_275) );
AOI33xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_285), .A3(n_297), .B1(n_309), .B2(n_310), .B3(n_315), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_278), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_278), .A2(n_316), .B1(n_462), .B2(n_477), .Y(n_461) );
INVx2_ASAP7_75t_L g1040 ( .A(n_278), .Y(n_1040) );
OR2x6_ASAP7_75t_L g278 ( .A(n_279), .B(n_283), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx2_ASAP7_75t_SL g605 ( .A(n_280), .Y(n_605) );
BUFx3_ASAP7_75t_L g650 ( .A(n_280), .Y(n_650) );
INVx1_ASAP7_75t_L g763 ( .A(n_280), .Y(n_763) );
INVx1_ASAP7_75t_L g855 ( .A(n_280), .Y(n_855) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
AND2x4_ASAP7_75t_L g319 ( .A(n_281), .B(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_282), .Y(n_320) );
INVx2_ASAP7_75t_L g531 ( .A(n_283), .Y(n_531) );
AND2x2_ASAP7_75t_L g568 ( .A(n_283), .B(n_403), .Y(n_568) );
BUFx2_ASAP7_75t_L g670 ( .A(n_283), .Y(n_670) );
OR2x2_ASAP7_75t_L g854 ( .A(n_283), .B(n_855), .Y(n_854) );
AND2x4_ASAP7_75t_L g1108 ( .A(n_283), .B(n_385), .Y(n_1108) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx2_ASAP7_75t_L g436 ( .A(n_284), .Y(n_436) );
OR2x6_ASAP7_75t_L g561 ( .A(n_284), .B(n_562), .Y(n_561) );
BUFx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
BUFx3_ASAP7_75t_L g311 ( .A(n_287), .Y(n_311) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_SL g449 ( .A(n_288), .Y(n_449) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_288), .Y(n_474) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_288), .Y(n_485) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_288), .Y(n_604) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_288), .Y(n_661) );
BUFx3_ASAP7_75t_L g863 ( .A(n_288), .Y(n_863) );
BUFx2_ASAP7_75t_L g955 ( .A(n_288), .Y(n_955) );
HB1xp67_ASAP7_75t_L g975 ( .A(n_288), .Y(n_975) );
BUFx2_ASAP7_75t_L g1364 ( .A(n_288), .Y(n_1364) );
AND2x4_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx1_ASAP7_75t_L g455 ( .A(n_289), .Y(n_455) );
INVx2_ASAP7_75t_L g302 ( .A(n_290), .Y(n_302) );
AND2x2_ASAP7_75t_L g308 ( .A(n_290), .B(n_295), .Y(n_308) );
BUFx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OR2x6_ASAP7_75t_L g443 ( .A(n_293), .B(n_440), .Y(n_443) );
OR2x2_ASAP7_75t_L g538 ( .A(n_293), .B(n_440), .Y(n_538) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_294), .Y(n_314) );
INVx1_ASAP7_75t_L g476 ( .A(n_294), .Y(n_476) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_294), .Y(n_487) );
INVx2_ASAP7_75t_L g594 ( .A(n_294), .Y(n_594) );
AND2x4_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx2_ASAP7_75t_L g303 ( .A(n_295), .Y(n_303) );
INVx1_ASAP7_75t_L g454 ( .A(n_296), .Y(n_454) );
BUFx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g438 ( .A(n_299), .B(n_439), .Y(n_438) );
A2O1A1Ixp33_ASAP7_75t_L g620 ( .A1(n_299), .A2(n_621), .B(n_622), .C(n_628), .Y(n_620) );
INVx2_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g758 ( .A(n_300), .Y(n_758) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g445 ( .A(n_301), .B(n_328), .Y(n_445) );
INVx6_ASAP7_75t_L g618 ( .A(n_301), .Y(n_618) );
AND2x4_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g326 ( .A(n_302), .Y(n_326) );
INVx1_ASAP7_75t_L g338 ( .A(n_303), .Y(n_338) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g1037 ( .A(n_306), .Y(n_1037) );
AND2x4_ASAP7_75t_L g1088 ( .A(n_306), .B(n_1089), .Y(n_1088) );
BUFx6f_ASAP7_75t_L g1365 ( .A(n_306), .Y(n_1365) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g343 ( .A(n_307), .Y(n_343) );
INVx2_ASAP7_75t_L g648 ( .A(n_307), .Y(n_648) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_308), .Y(n_599) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_314), .Y(n_654) );
INVx1_ASAP7_75t_L g663 ( .A(n_314), .Y(n_663) );
BUFx6f_ASAP7_75t_L g747 ( .A(n_314), .Y(n_747) );
INVx1_ASAP7_75t_L g824 ( .A(n_314), .Y(n_824) );
BUFx6f_ASAP7_75t_L g1085 ( .A(n_314), .Y(n_1085) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx4_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AOI221xp5_ASAP7_75t_L g1034 ( .A1(n_317), .A2(n_1035), .B1(n_1040), .B2(n_1041), .C(n_1049), .Y(n_1034) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AND2x4_ASAP7_75t_L g444 ( .A(n_318), .B(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g864 ( .A(n_318), .B(n_319), .Y(n_864) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_319), .Y(n_619) );
INVx2_ASAP7_75t_SL g659 ( .A(n_319), .Y(n_659) );
INVx1_ASAP7_75t_L g839 ( .A(n_319), .Y(n_839) );
OAI221xp5_ASAP7_75t_L g951 ( .A1(n_319), .A2(n_541), .B1(n_623), .B2(n_914), .C(n_917), .Y(n_951) );
OAI221xp5_ASAP7_75t_L g976 ( .A1(n_319), .A2(n_541), .B1(n_623), .B2(n_977), .C(n_978), .Y(n_976) );
INVx2_ASAP7_75t_L g1069 ( .A(n_319), .Y(n_1069) );
AND2x4_ASAP7_75t_L g328 ( .A(n_320), .B(n_329), .Y(n_328) );
AOI221xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_333), .B1(n_334), .B2(n_340), .C(n_341), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g865 ( .A1(n_322), .A2(n_341), .B1(n_866), .B2(n_867), .C(n_868), .Y(n_865) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x6_ASAP7_75t_L g323 ( .A(n_324), .B(n_327), .Y(n_323) );
OR2x2_ASAP7_75t_L g1052 ( .A(n_324), .B(n_327), .Y(n_1052) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_325), .A2(n_625), .B1(n_626), .B2(n_627), .Y(n_624) );
AND2x4_ASAP7_75t_L g668 ( .A(n_325), .B(n_328), .Y(n_668) );
AND2x2_ASAP7_75t_L g768 ( .A(n_325), .B(n_328), .Y(n_768) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_325), .B(n_328), .Y(n_1077) );
BUFx3_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_SL g339 ( .A(n_327), .Y(n_339) );
INVx1_ASAP7_75t_L g344 ( .A(n_327), .Y(n_344) );
NAND2x1p5_ASAP7_75t_L g327 ( .A(n_328), .B(n_331), .Y(n_327) );
BUFx2_ASAP7_75t_L g629 ( .A(n_328), .Y(n_629) );
AND2x4_ASAP7_75t_L g666 ( .A(n_328), .B(n_625), .Y(n_666) );
AND2x4_ASAP7_75t_L g766 ( .A(n_328), .B(n_625), .Y(n_766) );
INVx1_ASAP7_75t_L g1090 ( .A(n_328), .Y(n_1090) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x6_ASAP7_75t_L g709 ( .A(n_331), .B(n_404), .Y(n_709) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g440 ( .A(n_332), .B(n_441), .Y(n_440) );
AND2x4_ASAP7_75t_L g552 ( .A(n_332), .B(n_351), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_333), .A2(n_340), .B1(n_421), .B2(n_424), .Y(n_420) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_335), .Y(n_490) );
INVx2_ASAP7_75t_L g866 ( .A(n_335), .Y(n_866) );
INVx2_ASAP7_75t_L g1051 ( .A(n_335), .Y(n_1051) );
NAND2x1p5_ASAP7_75t_L g335 ( .A(n_336), .B(n_339), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g625 ( .A(n_337), .Y(n_625) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
BUFx2_ASAP7_75t_L g488 ( .A(n_341), .Y(n_488) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_344), .B(n_859), .Y(n_1053) );
OAI31xp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_362), .A3(n_426), .B(n_435), .Y(n_345) );
INVx3_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AOI221x1_ASAP7_75t_L g870 ( .A1(n_348), .A2(n_431), .B1(n_871), .B2(n_872), .C(n_873), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_348), .A2(n_431), .B1(n_1023), .B2(n_1024), .Y(n_1022) );
AND2x4_ASAP7_75t_L g348 ( .A(n_349), .B(n_353), .Y(n_348) );
AND2x4_ASAP7_75t_L g358 ( .A(n_349), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x4_ASAP7_75t_L g428 ( .A(n_351), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g431 ( .A(n_351), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g405 ( .A(n_352), .Y(n_405) );
INVx1_ASAP7_75t_L g563 ( .A(n_352), .Y(n_563) );
INVx1_ASAP7_75t_L g879 ( .A(n_353), .Y(n_879) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g566 ( .A(n_354), .Y(n_566) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_355), .Y(n_372) );
INVx3_ASAP7_75t_L g392 ( .A(n_355), .Y(n_392) );
AND2x4_ASAP7_75t_L g360 ( .A(n_356), .B(n_361), .Y(n_360) );
INVx8_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AOI221xp5_ASAP7_75t_SL g882 ( .A1(n_358), .A2(n_883), .B1(n_886), .B2(n_889), .C(n_890), .Y(n_882) );
BUFx6f_ASAP7_75t_L g888 ( .A(n_359), .Y(n_888) );
BUFx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_360), .Y(n_506) );
BUFx3_ASAP7_75t_L g575 ( .A(n_360), .Y(n_575) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_360), .Y(n_583) );
BUFx2_ASAP7_75t_L g780 ( .A(n_360), .Y(n_780) );
OAI221xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_373), .B1(n_386), .B2(n_394), .C(n_407), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B1(n_370), .B2(n_371), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_365), .A2(n_697), .B1(n_698), .B2(n_699), .Y(n_696) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_SL g387 ( .A(n_366), .Y(n_387) );
INVx2_ASAP7_75t_L g794 ( .A(n_366), .Y(n_794) );
BUFx3_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g496 ( .A(n_367), .Y(n_496) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g555 ( .A(n_368), .Y(n_555) );
BUFx2_ASAP7_75t_L g719 ( .A(n_368), .Y(n_719) );
INVx1_ASAP7_75t_L g425 ( .A(n_369), .Y(n_425) );
AND2x4_ASAP7_75t_L g432 ( .A(n_369), .B(n_433), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_371), .A2(n_733), .B1(n_734), .B2(n_736), .Y(n_732) );
INVx2_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_SL g526 ( .A(n_372), .Y(n_526) );
INVx4_ASAP7_75t_L g796 ( .A(n_372), .Y(n_796) );
BUFx3_ASAP7_75t_L g1115 ( .A(n_372), .Y(n_1115) );
OAI221xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_378), .B1(n_379), .B2(n_382), .C(n_383), .Y(n_373) );
OAI22xp33_ASAP7_75t_L g1006 ( .A1(n_374), .A2(n_705), .B1(n_980), .B2(n_985), .Y(n_1006) );
OAI21xp5_ASAP7_75t_SL g1029 ( .A1(n_374), .A2(n_1030), .B(n_1031), .Y(n_1029) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx3_ASAP7_75t_L g419 ( .A(n_375), .Y(n_419) );
BUFx2_ASAP7_75t_L g518 ( .A(n_375), .Y(n_518) );
INVx2_ASAP7_75t_L g528 ( .A(n_375), .Y(n_528) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_376), .B(n_377), .Y(n_396) );
INVx1_ASAP7_75t_L g777 ( .A(n_377), .Y(n_777) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g925 ( .A(n_380), .Y(n_925) );
INVx2_ASAP7_75t_SL g1408 ( .A(n_380), .Y(n_1408) );
INVx2_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx2_ASAP7_75t_SL g521 ( .A(n_385), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B1(n_389), .B2(n_393), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_388), .A2(n_397), .B1(n_447), .B2(n_450), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g928 ( .A1(n_389), .A2(n_929), .B1(n_930), .B2(n_931), .Y(n_928) );
OAI22xp5_ASAP7_75t_L g1001 ( .A1(n_389), .A2(n_930), .B1(n_1002), .B2(n_1003), .Y(n_1001) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g885 ( .A(n_391), .Y(n_885) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx3_ASAP7_75t_L g501 ( .A(n_392), .Y(n_501) );
INVx3_ASAP7_75t_L g558 ( .A(n_392), .Y(n_558) );
AOI222xp33_ASAP7_75t_L g437 ( .A1(n_393), .A2(n_400), .B1(n_417), .B2(n_438), .C1(n_442), .C2(n_444), .Y(n_437) );
OAI221xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_397), .B1(n_398), .B2(n_400), .C(n_401), .Y(n_394) );
BUFx3_ASAP7_75t_L g706 ( .A(n_395), .Y(n_706) );
BUFx3_ASAP7_75t_L g728 ( .A(n_395), .Y(n_728) );
OAI22xp33_ASAP7_75t_L g729 ( .A1(n_395), .A2(n_705), .B1(n_730), .B2(n_731), .Y(n_729) );
INVx2_ASAP7_75t_L g810 ( .A(n_395), .Y(n_810) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI22xp5_ASAP7_75t_SL g806 ( .A1(n_398), .A2(n_807), .B1(n_808), .B2(n_809), .Y(n_806) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx2_ASAP7_75t_L g507 ( .A(n_404), .Y(n_507) );
NAND2x1p5_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_417), .B(n_418), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NOR2xp67_ASAP7_75t_L g535 ( .A(n_409), .B(n_531), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_414), .Y(n_409) );
AND2x2_ASAP7_75t_L g510 ( .A(n_410), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI21xp33_ASAP7_75t_L g418 ( .A1(n_411), .A2(n_419), .B(n_420), .Y(n_418) );
OR2x6_ASAP7_75t_L g514 ( .A(n_411), .B(n_425), .Y(n_514) );
OR2x2_ASAP7_75t_L g527 ( .A(n_411), .B(n_528), .Y(n_527) );
OR2x6_ASAP7_75t_L g881 ( .A(n_411), .B(n_528), .Y(n_881) );
INVx1_ASAP7_75t_L g892 ( .A(n_411), .Y(n_892) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
BUFx2_ASAP7_75t_L g504 ( .A(n_414), .Y(n_504) );
AND2x2_ASAP7_75t_L g551 ( .A(n_414), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_SL g683 ( .A(n_415), .Y(n_683) );
INVx2_ASAP7_75t_L g895 ( .A(n_415), .Y(n_895) );
INVx3_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_416), .Y(n_429) );
OAI21xp5_ASAP7_75t_SL g874 ( .A1(n_419), .A2(n_875), .B(n_876), .Y(n_874) );
BUFx2_ASAP7_75t_L g1352 ( .A(n_419), .Y(n_1352) );
NAND2x1_ASAP7_75t_SL g570 ( .A(n_421), .B(n_571), .Y(n_570) );
NAND2x1p5_ASAP7_75t_L g891 ( .A(n_421), .B(n_892), .Y(n_891) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_423), .Y(n_511) );
NAND2x1p5_ASAP7_75t_L g573 ( .A(n_424), .B(n_571), .Y(n_573) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
CKINVDCx6p67_ASAP7_75t_R g427 ( .A(n_428), .Y(n_427) );
BUFx2_ASAP7_75t_L g887 ( .A(n_429), .Y(n_887) );
INVx3_ASAP7_75t_L g1111 ( .A(n_429), .Y(n_1111) );
INVx3_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_432), .Y(n_580) );
BUFx6f_ASAP7_75t_L g884 ( .A(n_432), .Y(n_884) );
INVx1_ASAP7_75t_L g1015 ( .A(n_432), .Y(n_1015) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g630 ( .A(n_435), .Y(n_630) );
BUFx8_ASAP7_75t_SL g1368 ( .A(n_435), .Y(n_1368) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g771 ( .A(n_436), .Y(n_771) );
AOI221xp5_ASAP7_75t_L g1054 ( .A1(n_438), .A2(n_447), .B1(n_1055), .B2(n_1056), .C(n_1057), .Y(n_1054) );
AND2x2_ASAP7_75t_L g447 ( .A(n_439), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OR2x6_ASAP7_75t_L g451 ( .A(n_440), .B(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g540 ( .A(n_440), .B(n_541), .Y(n_540) );
OR2x2_ASAP7_75t_L g542 ( .A(n_440), .B(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g592 ( .A(n_441), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_441), .B(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g596 ( .A(n_441), .B(n_466), .Y(n_596) );
A2O1A1Ixp33_ASAP7_75t_L g744 ( .A1(n_441), .A2(n_745), .B(n_748), .C(n_750), .Y(n_744) );
CKINVDCx6p67_ASAP7_75t_R g442 ( .A(n_443), .Y(n_442) );
OR2x6_ASAP7_75t_L g534 ( .A(n_444), .B(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g674 ( .A(n_444), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_445), .B(n_770), .Y(n_769) );
INVx2_ASAP7_75t_L g815 ( .A(n_445), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_448), .A2(n_731), .B1(n_733), .B2(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_SL g857 ( .A(n_449), .Y(n_857) );
INVx1_ASAP7_75t_L g950 ( .A(n_449), .Y(n_950) );
OAI22xp5_ASAP7_75t_L g1039 ( .A1(n_449), .A2(n_663), .B1(n_1027), .B2(n_1028), .Y(n_1039) );
CKINVDCx6p67_ASAP7_75t_R g450 ( .A(n_451), .Y(n_450) );
OAI21xp33_ASAP7_75t_L g601 ( .A1(n_452), .A2(n_602), .B(n_603), .Y(n_601) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx4f_ASAP7_75t_L g470 ( .A(n_453), .Y(n_470) );
INVx1_ASAP7_75t_L g614 ( .A(n_453), .Y(n_614) );
INVx1_ASAP7_75t_L g623 ( .A(n_453), .Y(n_623) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
OR2x2_ASAP7_75t_L g466 ( .A(n_454), .B(n_455), .Y(n_466) );
AO22x2_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_458), .B1(n_544), .B2(n_545), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND4x1_ASAP7_75t_L g459 ( .A(n_460), .B(n_491), .C(n_532), .D(n_536), .Y(n_459) );
NOR3xp33_ASAP7_75t_L g460 ( .A(n_461), .B(n_488), .C(n_489), .Y(n_460) );
OAI221xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_467), .B1(n_468), .B2(n_471), .C(n_472), .Y(n_462) );
BUFx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OAI221xp5_ASAP7_75t_SL g823 ( .A1(n_464), .A2(n_795), .B1(n_799), .B2(n_824), .C(n_825), .Y(n_823) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g479 ( .A(n_466), .Y(n_479) );
INVx1_ASAP7_75t_L g609 ( .A(n_466), .Y(n_609) );
OAI221xp5_ASAP7_75t_L g516 ( .A1(n_467), .A2(n_471), .B1(n_517), .B2(n_519), .C(n_521), .Y(n_516) );
BUFx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OAI211xp5_ASAP7_75t_L g759 ( .A1(n_469), .A2(n_727), .B(n_760), .C(n_762), .Y(n_759) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g481 ( .A(n_470), .Y(n_481) );
BUFx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g543 ( .A(n_474), .Y(n_543) );
AND2x2_ASAP7_75t_L g591 ( .A(n_474), .B(n_592), .Y(n_591) );
BUFx4f_ASAP7_75t_L g1046 ( .A(n_474), .Y(n_1046) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OAI221xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_480), .B1(n_481), .B2(n_482), .C(n_483), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g541 ( .A(n_479), .Y(n_541) );
BUFx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x4_ASAP7_75t_L g947 ( .A(n_485), .B(n_592), .Y(n_947) );
INVx2_ASAP7_75t_SL g1072 ( .A(n_485), .Y(n_1072) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OAI31xp33_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_515), .A3(n_529), .B(n_530), .Y(n_491) );
OAI221xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_497), .B1(n_498), .B2(n_502), .C(n_503), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g524 ( .A(n_495), .Y(n_524) );
INVx1_ASAP7_75t_L g933 ( .A(n_495), .Y(n_933) );
INVx2_ASAP7_75t_L g1005 ( .A(n_495), .Y(n_1005) );
INVx2_ASAP7_75t_L g1341 ( .A(n_495), .Y(n_1341) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_496), .A2(n_878), .B1(n_879), .B2(n_880), .Y(n_877) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g1347 ( .A1(n_500), .A2(n_1341), .B1(n_1348), .B2(n_1349), .Y(n_1347) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g586 ( .A(n_501), .B(n_552), .Y(n_586) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_501), .Y(n_722) );
INVx1_ASAP7_75t_L g804 ( .A(n_501), .Y(n_804) );
INVx2_ASAP7_75t_L g937 ( .A(n_501), .Y(n_937) );
INVx2_ASAP7_75t_L g1413 ( .A(n_501), .Y(n_1413) );
BUFx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_SL g1020 ( .A(n_506), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B1(n_512), .B2(n_513), .Y(n_508) );
AND2x4_ASAP7_75t_L g773 ( .A(n_511), .B(n_571), .Y(n_773) );
CKINVDCx11_ASAP7_75t_R g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g927 ( .A(n_518), .Y(n_927) );
OAI22xp33_ASAP7_75t_L g691 ( .A1(n_519), .A2(n_692), .B1(n_693), .B2(n_695), .Y(n_691) );
OAI22xp33_ASAP7_75t_L g1343 ( .A1(n_519), .A2(n_1344), .B1(n_1345), .B2(n_1346), .Y(n_1343) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OAI22xp5_ASAP7_75t_SL g522 ( .A1(n_523), .A2(n_524), .B1(n_525), .B2(n_526), .Y(n_522) );
INVx1_ASAP7_75t_L g694 ( .A(n_528), .Y(n_694) );
OAI22xp33_ASAP7_75t_L g797 ( .A1(n_528), .A2(n_725), .B1(n_798), .B2(n_799), .Y(n_797) );
AOI31xp33_ASAP7_75t_L g1064 ( .A1(n_530), .A2(n_1065), .A3(n_1078), .B(n_1091), .Y(n_1064) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g968 ( .A1(n_531), .A2(n_964), .B1(n_969), .B2(n_987), .Y(n_968) );
AOI22xp5_ASAP7_75t_L g1379 ( .A1(n_531), .A2(n_672), .B1(n_1380), .B2(n_1395), .Y(n_1379) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g1032 ( .A(n_534), .B(n_1033), .Y(n_1032) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .Y(n_536) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND3xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_576), .C(n_588), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_569), .Y(n_548) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g579 ( .A(n_552), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g582 ( .A(n_552), .B(n_583), .Y(n_582) );
AND2x4_ASAP7_75t_L g682 ( .A(n_552), .B(n_683), .Y(n_682) );
AND2x4_ASAP7_75t_L g846 ( .A(n_552), .B(n_558), .Y(n_846) );
AND2x6_ASAP7_75t_L g915 ( .A(n_552), .B(n_575), .Y(n_915) );
AND2x2_ASAP7_75t_L g919 ( .A(n_552), .B(n_580), .Y(n_919) );
AND2x2_ASAP7_75t_L g995 ( .A(n_552), .B(n_580), .Y(n_995) );
OAI221xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_556), .B1(n_557), .B2(n_559), .C(n_560), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_555), .Y(n_702) );
INVx1_ASAP7_75t_L g735 ( .A(n_555), .Y(n_735) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g698 ( .A(n_558), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_559), .A2(n_607), .B1(n_608), .B2(n_610), .Y(n_606) );
OAI33xp33_ASAP7_75t_L g690 ( .A1(n_561), .A2(n_691), .A3(n_696), .B1(n_700), .B2(n_704), .B3(n_707), .Y(n_690) );
OAI33xp33_ASAP7_75t_L g922 ( .A1(n_561), .A2(n_923), .A3(n_928), .B1(n_932), .B2(n_939), .B3(n_942), .Y(n_922) );
OAI33xp33_ASAP7_75t_L g997 ( .A1(n_561), .A2(n_942), .A3(n_998), .B1(n_1001), .B2(n_1004), .B3(n_1006), .Y(n_997) );
OAI33xp33_ASAP7_75t_L g1338 ( .A1(n_561), .A2(n_942), .A3(n_1339), .B1(n_1343), .B2(n_1347), .B3(n_1350), .Y(n_1338) );
OAI33xp33_ASAP7_75t_L g1406 ( .A1(n_561), .A2(n_942), .A3(n_1407), .B1(n_1411), .B2(n_1415), .B3(n_1418), .Y(n_1406) );
NAND3xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .C(n_568), .Y(n_564) );
INVx1_ASAP7_75t_L g703 ( .A(n_566), .Y(n_703) );
INVx2_ASAP7_75t_L g687 ( .A(n_570), .Y(n_687) );
HB1xp67_ASAP7_75t_L g1405 ( .A(n_570), .Y(n_1405) );
NAND2x1p5_ASAP7_75t_L g574 ( .A(n_571), .B(n_575), .Y(n_574) );
AND2x4_ASAP7_75t_L g775 ( .A(n_571), .B(n_776), .Y(n_775) );
AND2x4_ASAP7_75t_L g779 ( .A(n_571), .B(n_780), .Y(n_779) );
INVx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
BUFx4f_ASAP7_75t_L g688 ( .A(n_573), .Y(n_688) );
BUFx4f_ASAP7_75t_L g790 ( .A(n_573), .Y(n_790) );
BUFx3_ASAP7_75t_L g689 ( .A(n_574), .Y(n_689) );
BUFx2_ASAP7_75t_L g921 ( .A(n_574), .Y(n_921) );
NOR2xp33_ASAP7_75t_SL g576 ( .A(n_577), .B(n_584), .Y(n_576) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_579), .A2(n_681), .B1(n_682), .B2(n_684), .Y(n_680) );
INVx1_ASAP7_75t_L g740 ( .A(n_579), .Y(n_740) );
INVx1_ASAP7_75t_L g789 ( .A(n_579), .Y(n_789) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_582), .A2(n_586), .B1(n_678), .B2(n_679), .Y(n_677) );
INVxp67_ASAP7_75t_L g741 ( .A(n_582), .Y(n_741) );
INVx2_ASAP7_75t_SL g1113 ( .A(n_583), .Y(n_1113) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x4_ASAP7_75t_L g673 ( .A(n_587), .B(n_674), .Y(n_673) );
OAI31xp33_ASAP7_75t_SL g588 ( .A1(n_589), .A2(n_595), .A3(n_600), .B(n_630), .Y(n_588) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_591), .A2(n_657), .B1(n_658), .B2(n_660), .C(n_664), .Y(n_656) );
AOI221xp5_ASAP7_75t_L g1381 ( .A1(n_591), .A2(n_1382), .B1(n_1383), .B2(n_1384), .C(n_1385), .Y(n_1381) );
AND2x4_ASAP7_75t_L g598 ( .A(n_592), .B(n_599), .Y(n_598) );
AOI221xp5_ASAP7_75t_L g821 ( .A1(n_592), .A2(n_598), .B1(n_655), .B2(n_808), .C(n_822), .Y(n_821) );
INVx4_ASAP7_75t_L g642 ( .A(n_593), .Y(n_642) );
INVx1_ASAP7_75t_L g611 ( .A(n_594), .Y(n_611) );
INVx2_ASAP7_75t_L g833 ( .A(n_594), .Y(n_833) );
INVx6_ASAP7_75t_L g640 ( .A(n_596), .Y(n_640) );
INVx1_ASAP7_75t_L g644 ( .A(n_597), .Y(n_644) );
INVx2_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
HB1xp67_ASAP7_75t_L g953 ( .A(n_598), .Y(n_953) );
AOI221xp5_ASAP7_75t_L g979 ( .A1(n_598), .A2(n_655), .B1(n_980), .B2(n_981), .C(n_983), .Y(n_979) );
BUFx6f_ASAP7_75t_L g1086 ( .A(n_598), .Y(n_1086) );
AOI221xp5_ASAP7_75t_L g1387 ( .A1(n_598), .A2(n_655), .B1(n_1388), .B2(n_1389), .C(n_1391), .Y(n_1387) );
AND2x4_ASAP7_75t_L g655 ( .A(n_599), .B(n_629), .Y(n_655) );
BUFx4f_ASAP7_75t_L g749 ( .A(n_599), .Y(n_749) );
INVx1_ASAP7_75t_L g837 ( .A(n_599), .Y(n_837) );
BUFx6f_ASAP7_75t_L g859 ( .A(n_599), .Y(n_859) );
INVx2_ASAP7_75t_SL g957 ( .A(n_599), .Y(n_957) );
OAI211xp5_ASAP7_75t_SL g600 ( .A1(n_601), .A2(n_606), .B(n_612), .C(n_620), .Y(n_600) );
BUFx3_ASAP7_75t_L g828 ( .A(n_604), .Y(n_828) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OAI211xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_614), .B(n_615), .C(n_616), .Y(n_612) );
BUFx6f_ASAP7_75t_L g960 ( .A(n_617), .Y(n_960) );
INVx1_ASAP7_75t_L g1082 ( .A(n_617), .Y(n_1082) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_618), .Y(n_653) );
INVx2_ASAP7_75t_L g746 ( .A(n_618), .Y(n_746) );
INVx1_ASAP7_75t_L g761 ( .A(n_618), .Y(n_761) );
INVx1_ASAP7_75t_L g838 ( .A(n_618), .Y(n_838) );
NAND2xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx1_ASAP7_75t_L g755 ( .A(n_623), .Y(n_755) );
BUFx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g944 ( .A1(n_630), .A2(n_945), .B1(n_963), .B2(n_964), .Y(n_944) );
INVx1_ASAP7_75t_L g901 ( .A(n_631), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_783), .B1(n_784), .B2(n_899), .Y(n_631) );
INVx1_ASAP7_75t_L g899 ( .A(n_632), .Y(n_899) );
XNOR2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_712), .Y(n_632) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g710 ( .A(n_635), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_675), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_669), .B1(n_671), .B2(n_672), .Y(n_636) );
NAND3xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_643), .C(n_656), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_640), .B1(n_641), .B2(n_642), .Y(n_638) );
OAI22xp33_ASAP7_75t_L g704 ( .A1(n_639), .A2(n_645), .B1(n_705), .B2(n_706), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_640), .A2(n_642), .B1(n_938), .B2(n_940), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_640), .A2(n_642), .B1(n_985), .B2(n_986), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_640), .A2(n_642), .B1(n_1092), .B2(n_1093), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g1367 ( .A1(n_640), .A2(n_642), .B1(n_1349), .B2(n_1351), .Y(n_1367) );
AOI22xp33_ASAP7_75t_L g1392 ( .A1(n_640), .A2(n_642), .B1(n_1393), .B2(n_1394), .Y(n_1392) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_641), .A2(n_657), .B1(n_701), .B2(n_703), .Y(n_700) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .B1(n_646), .B2(n_651), .C(n_655), .Y(n_643) );
INVx3_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g861 ( .A(n_648), .Y(n_861) );
INVx3_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVxp67_ASAP7_75t_L g958 ( .A(n_650), .Y(n_958) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx4_ASAP7_75t_L g1067 ( .A(n_653), .Y(n_1067) );
INVx1_ASAP7_75t_L g750 ( .A(n_655), .Y(n_750) );
AOI221xp5_ASAP7_75t_L g952 ( .A1(n_655), .A2(n_941), .B1(n_953), .B2(n_954), .C(n_959), .Y(n_952) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g961 ( .A(n_663), .Y(n_961) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
INVx4_ASAP7_75t_L g818 ( .A(n_666), .Y(n_818) );
INVx2_ASAP7_75t_L g1386 ( .A(n_666), .Y(n_1386) );
INVx2_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
AOI222xp33_ASAP7_75t_SL g813 ( .A1(n_668), .A2(n_814), .B1(n_816), .B2(n_817), .C1(n_819), .C2(n_820), .Y(n_813) );
INVx2_ASAP7_75t_L g973 ( .A(n_668), .Y(n_973) );
CKINVDCx8_ASAP7_75t_R g669 ( .A(n_670), .Y(n_669) );
OAI21xp5_ASAP7_75t_SL g1010 ( .A1(n_670), .A2(n_1011), .B(n_1025), .Y(n_1010) );
INVx2_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g964 ( .A(n_673), .Y(n_964) );
INVx5_ASAP7_75t_L g1062 ( .A(n_673), .Y(n_1062) );
NOR3xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_685), .C(n_690), .Y(n_675) );
NAND2xp5_ASAP7_75t_SL g676 ( .A(n_677), .B(n_680), .Y(n_676) );
INVx1_ASAP7_75t_L g843 ( .A(n_682), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_682), .A2(n_917), .B1(n_918), .B2(n_919), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_682), .A2(n_978), .B1(n_994), .B2(n_995), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_682), .A2(n_919), .B1(n_1103), .B2(n_1104), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g1333 ( .A1(n_682), .A2(n_919), .B1(n_1334), .B2(n_1335), .Y(n_1333) );
AOI22xp33_ASAP7_75t_L g1401 ( .A1(n_682), .A2(n_995), .B1(n_1402), .B2(n_1403), .Y(n_1401) );
INVx1_ASAP7_75t_L g1018 ( .A(n_683), .Y(n_1018) );
BUFx3_ASAP7_75t_L g1119 ( .A(n_683), .Y(n_1119) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx2_ASAP7_75t_SL g1337 ( .A(n_687), .Y(n_1337) );
OAI22xp33_ASAP7_75t_L g1418 ( .A1(n_693), .A2(n_1391), .B1(n_1393), .B2(n_1408), .Y(n_1418) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g1026 ( .A1(n_698), .A2(n_701), .B1(n_1027), .B2(n_1028), .Y(n_1026) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g737 ( .A(n_708), .Y(n_737) );
AOI33xp33_ASAP7_75t_L g1105 ( .A1(n_708), .A2(n_1106), .A3(n_1109), .B1(n_1114), .B2(n_1116), .B3(n_1118), .Y(n_1105) );
INVx6_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx5_ASAP7_75t_L g943 ( .A(n_709), .Y(n_943) );
OAI22xp33_ASAP7_75t_L g1155 ( .A1(n_711), .A2(n_1156), .B1(n_1158), .B2(n_1159), .Y(n_1155) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_SL g782 ( .A(n_714), .Y(n_782) );
NAND4xp75_ASAP7_75t_L g714 ( .A(n_715), .B(n_738), .C(n_743), .D(n_772), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B1(n_720), .B2(n_721), .Y(n_716) );
BUFx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g803 ( .A(n_719), .Y(n_803) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OAI22xp33_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_725), .B1(n_727), .B2(n_728), .Y(n_723) );
OAI22xp33_ASAP7_75t_L g1350 ( .A1(n_725), .A2(n_1351), .B1(n_1352), .B2(n_1353), .Y(n_1350) );
INVx3_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OAI22xp33_ASAP7_75t_L g998 ( .A1(n_728), .A2(n_925), .B1(n_999), .B2(n_1000), .Y(n_998) );
OAI22xp33_ASAP7_75t_L g1407 ( .A1(n_728), .A2(n_1408), .B1(n_1409), .B2(n_1410), .Y(n_1407) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_730), .A2(n_736), .B1(n_746), .B2(n_747), .Y(n_745) );
BUFx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
BUFx2_ASAP7_75t_L g930 ( .A(n_735), .Y(n_930) );
NOR2x1_ASAP7_75t_L g738 ( .A(n_739), .B(n_742), .Y(n_738) );
OAI31xp33_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_751), .A3(n_764), .B(n_771), .Y(n_743) );
HB1xp67_ASAP7_75t_L g1038 ( .A(n_746), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_759), .Y(n_751) );
OAI211xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_754), .B(n_756), .C(n_757), .Y(n_752) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g1075 ( .A(n_766), .Y(n_1075) );
INVx3_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g841 ( .A(n_771), .Y(n_841) );
AOI21x1_ASAP7_75t_L g869 ( .A1(n_771), .A2(n_870), .B(n_882), .Y(n_869) );
AOI221xp5_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_774), .B1(n_775), .B2(n_778), .C(n_779), .Y(n_772) );
AOI21xp5_ASAP7_75t_L g847 ( .A1(n_773), .A2(n_779), .B(n_819), .Y(n_847) );
AOI221xp5_ASAP7_75t_L g1095 ( .A1(n_773), .A2(n_775), .B1(n_779), .B2(n_1096), .C(n_1097), .Y(n_1095) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
AO22x2_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_848), .B1(n_849), .B2(n_898), .Y(n_784) );
INVx1_ASAP7_75t_L g898 ( .A(n_785), .Y(n_898) );
AND2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_811), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_791), .Y(n_787) );
OAI22xp33_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_794), .B1(n_795), .B2(n_796), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g1004 ( .A1(n_796), .A2(n_971), .B1(n_986), .B2(n_1005), .Y(n_1004) );
INVx2_ASAP7_75t_SL g1117 ( .A(n_796), .Y(n_1117) );
OAI22xp5_ASAP7_75t_L g1339 ( .A1(n_796), .A2(n_1340), .B1(n_1341), .B2(n_1342), .Y(n_1339) );
OAI22xp5_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_802), .B1(n_804), .B2(n_805), .Y(n_800) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
OAI22xp33_ASAP7_75t_L g939 ( .A1(n_809), .A2(n_925), .B1(n_940), .B2(n_941), .Y(n_939) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g1345 ( .A(n_810), .Y(n_1345) );
AOI21xp5_ASAP7_75t_SL g811 ( .A1(n_812), .A2(n_840), .B(n_842), .Y(n_811) );
NAND4xp25_ASAP7_75t_SL g812 ( .A(n_813), .B(n_821), .C(n_823), .D(n_826), .Y(n_812) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g1048 ( .A(n_824), .Y(n_1048) );
OAI221xp5_ASAP7_75t_L g826 ( .A1(n_827), .A2(n_829), .B1(n_830), .B2(n_834), .C(n_835), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx2_ASAP7_75t_SL g1390 ( .A(n_832), .Y(n_1390) );
INVx2_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
BUFx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
BUFx2_ASAP7_75t_L g913 ( .A(n_846), .Y(n_913) );
BUFx2_ASAP7_75t_L g992 ( .A(n_846), .Y(n_992) );
BUFx2_ASAP7_75t_L g1100 ( .A(n_846), .Y(n_1100) );
AOI22xp33_ASAP7_75t_L g1330 ( .A1(n_846), .A2(n_915), .B1(n_1331), .B2(n_1332), .Y(n_1330) );
AOI22xp33_ASAP7_75t_L g1398 ( .A1(n_846), .A2(n_915), .B1(n_1399), .B2(n_1400), .Y(n_1398) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
NOR4xp75_ASAP7_75t_L g850 ( .A(n_851), .B(n_869), .C(n_896), .D(n_897), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_852), .B(n_865), .Y(n_851) );
AOI33xp33_ASAP7_75t_L g852 ( .A1(n_853), .A2(n_856), .A3(n_858), .B1(n_860), .B2(n_862), .B3(n_864), .Y(n_852) );
INVx3_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g1043 ( .A(n_859), .Y(n_1043) );
OAI21xp5_ASAP7_75t_L g873 ( .A1(n_874), .A2(n_877), .B(n_881), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_894), .B(n_895), .Y(n_893) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
XNOR2xp5_ASAP7_75t_L g903 ( .A(n_904), .B(n_1007), .Y(n_903) );
AO22x2_ASAP7_75t_L g904 ( .A1(n_905), .A2(n_906), .B1(n_965), .B2(n_966), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
XNOR2xp5_ASAP7_75t_L g906 ( .A(n_907), .B(n_908), .Y(n_906) );
AND2x2_ASAP7_75t_L g908 ( .A(n_909), .B(n_944), .Y(n_908) );
NOR3xp33_ASAP7_75t_L g909 ( .A(n_910), .B(n_920), .C(n_922), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_911), .B(n_916), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_912), .A2(n_913), .B1(n_914), .B2(n_915), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_915), .A2(n_977), .B1(n_991), .B2(n_992), .Y(n_990) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_915), .A2(n_1099), .B1(n_1100), .B2(n_1101), .Y(n_1098) );
OAI22xp33_ASAP7_75t_L g923 ( .A1(n_924), .A2(n_925), .B1(n_926), .B2(n_927), .Y(n_923) );
OAI22xp5_ASAP7_75t_L g1411 ( .A1(n_930), .A2(n_1412), .B1(n_1413), .B2(n_1414), .Y(n_1411) );
OAI22xp5_ASAP7_75t_L g1415 ( .A1(n_930), .A2(n_1384), .B1(n_1394), .B2(n_1416), .Y(n_1415) );
OAI22xp5_ASAP7_75t_L g932 ( .A1(n_933), .A2(n_934), .B1(n_935), .B2(n_938), .Y(n_932) );
AOI211xp5_ASAP7_75t_SL g946 ( .A1(n_934), .A2(n_947), .B(n_948), .C(n_949), .Y(n_946) );
INVx1_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
INVx2_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g1417 ( .A(n_937), .Y(n_1417) );
CKINVDCx8_ASAP7_75t_R g942 ( .A(n_943), .Y(n_942) );
NAND3xp33_ASAP7_75t_L g945 ( .A(n_946), .B(n_952), .C(n_962), .Y(n_945) );
AOI211xp5_ASAP7_75t_SL g970 ( .A1(n_947), .A2(n_971), .B(n_972), .C(n_974), .Y(n_970) );
AOI221xp5_ASAP7_75t_L g1065 ( .A1(n_947), .A2(n_1066), .B1(n_1070), .B2(n_1073), .C(n_1074), .Y(n_1065) );
AOI221xp5_ASAP7_75t_L g1357 ( .A1(n_947), .A2(n_1348), .B1(n_1358), .B2(n_1359), .C(n_1361), .Y(n_1357) );
INVx1_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
INVx1_ASAP7_75t_L g982 ( .A(n_957), .Y(n_982) );
INVx1_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
AND2x2_ASAP7_75t_L g967 ( .A(n_968), .B(n_988), .Y(n_967) );
NAND3xp33_ASAP7_75t_L g969 ( .A(n_970), .B(n_979), .C(n_984), .Y(n_969) );
NOR3xp33_ASAP7_75t_SL g988 ( .A(n_989), .B(n_996), .C(n_997), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_990), .B(n_993), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_1008), .A2(n_1058), .B1(n_1120), .B2(n_1121), .Y(n_1007) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1008), .Y(n_1120) );
NAND4xp25_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1032), .C(n_1034), .D(n_1054), .Y(n_1009) );
AOI21xp5_ASAP7_75t_L g1012 ( .A1(n_1013), .A2(n_1016), .B(n_1021), .Y(n_1012) );
INVx2_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
INVx2_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
OAI22xp5_ASAP7_75t_L g1044 ( .A1(n_1023), .A2(n_1024), .B1(n_1045), .B2(n_1047), .Y(n_1044) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
INVx1_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
INVx1_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
INVxp67_ASAP7_75t_SL g1121 ( .A(n_1058), .Y(n_1121) );
XNOR2x1_ASAP7_75t_SL g1058 ( .A(n_1059), .B(n_1060), .Y(n_1058) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1094), .Y(n_1060) );
AOI21xp5_ASAP7_75t_L g1061 ( .A1(n_1062), .A2(n_1063), .B(n_1064), .Y(n_1061) );
AOI21xp33_ASAP7_75t_SL g1354 ( .A1(n_1062), .A2(n_1355), .B(n_1356), .Y(n_1354) );
BUFx2_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1072), .Y(n_1360) );
INVx2_ASAP7_75t_SL g1076 ( .A(n_1077), .Y(n_1076) );
AOI221xp5_ASAP7_75t_L g1078 ( .A1(n_1079), .A2(n_1080), .B1(n_1086), .B2(n_1087), .C(n_1088), .Y(n_1078) );
INVx2_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
INVx1_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
AOI221xp5_ASAP7_75t_L g1362 ( .A1(n_1086), .A2(n_1088), .B1(n_1353), .B2(n_1363), .C(n_1366), .Y(n_1362) );
INVx1_ASAP7_75t_SL g1089 ( .A(n_1090), .Y(n_1089) );
AND4x1_ASAP7_75t_L g1094 ( .A(n_1095), .B(n_1098), .C(n_1102), .D(n_1105), .Y(n_1094) );
INVx2_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
INVx2_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
INVx2_ASAP7_75t_SL g1110 ( .A(n_1111), .Y(n_1110) );
INVx2_ASAP7_75t_SL g1112 ( .A(n_1113), .Y(n_1112) );
OAI21xp33_ASAP7_75t_L g1122 ( .A1(n_1123), .A2(n_1131), .B(n_1324), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
INVx2_ASAP7_75t_L g1180 ( .A(n_1125), .Y(n_1180) );
INVx2_ASAP7_75t_L g1125 ( .A(n_1126), .Y(n_1125) );
AND2x4_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1129), .Y(n_1126) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1127), .Y(n_1151) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1142 ( .A(n_1128), .B(n_1143), .Y(n_1142) );
AND2x4_ASAP7_75t_L g1150 ( .A(n_1129), .B(n_1151), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1129), .B(n_1151), .Y(n_1196) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1130), .Y(n_1143) );
NOR3xp33_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1264), .C(n_1302), .Y(n_1131) );
AOI22xp5_ASAP7_75t_L g1132 ( .A1(n_1133), .A2(n_1200), .B1(n_1245), .B2(n_1253), .Y(n_1132) );
NOR3xp33_ASAP7_75t_SL g1133 ( .A(n_1134), .B(n_1210), .C(n_1213), .Y(n_1133) );
A2O1A1Ixp33_ASAP7_75t_L g1134 ( .A1(n_1135), .A2(n_1164), .B(n_1172), .C(n_1185), .Y(n_1134) );
O2A1O1Ixp33_ASAP7_75t_L g1320 ( .A1(n_1135), .A2(n_1137), .B(n_1321), .C(n_1322), .Y(n_1320) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1136), .B(n_1168), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1137), .B(n_1152), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1137), .B(n_1190), .Y(n_1256) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1137), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1137), .B(n_1219), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1137), .B(n_1223), .Y(n_1281) );
NOR2xp33_ASAP7_75t_L g1317 ( .A(n_1137), .B(n_1178), .Y(n_1317) );
INVx4_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
OR2x2_ASAP7_75t_L g1188 ( .A(n_1138), .B(n_1175), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1138), .B(n_1166), .Y(n_1212) );
INVx3_ASAP7_75t_L g1221 ( .A(n_1138), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1227 ( .A(n_1138), .B(n_1217), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1238 ( .A(n_1138), .B(n_1152), .Y(n_1238) );
NOR2xp67_ASAP7_75t_SL g1240 ( .A(n_1138), .B(n_1199), .Y(n_1240) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1138), .B(n_1168), .Y(n_1271) );
NAND3xp33_ASAP7_75t_L g1300 ( .A(n_1138), .B(n_1289), .C(n_1298), .Y(n_1300) );
AOI211xp5_ASAP7_75t_L g1304 ( .A1(n_1138), .A2(n_1232), .B(n_1305), .C(n_1306), .Y(n_1304) );
AND2x4_ASAP7_75t_L g1138 ( .A(n_1139), .B(n_1149), .Y(n_1138) );
AND2x4_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1144), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
OR2x2_ASAP7_75t_L g1157 ( .A(n_1142), .B(n_1145), .Y(n_1157) );
HB1xp67_ASAP7_75t_L g1428 ( .A(n_1143), .Y(n_1428) );
AND2x4_ASAP7_75t_L g1146 ( .A(n_1144), .B(n_1147), .Y(n_1146) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
OR2x2_ASAP7_75t_L g1159 ( .A(n_1145), .B(n_1148), .Y(n_1159) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1150), .Y(n_1203) );
HB1xp67_ASAP7_75t_L g1426 ( .A(n_1151), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1152), .B(n_1169), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1152), .B(n_1256), .Y(n_1279) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1152), .B(n_1271), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1153), .B(n_1160), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1217 ( .A(n_1153), .B(n_1167), .Y(n_1217) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1154), .B(n_1167), .Y(n_1166) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1154), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_1154), .B(n_1160), .Y(n_1244) );
OAI22xp5_ASAP7_75t_L g1161 ( .A1(n_1156), .A2(n_1159), .B1(n_1162), .B2(n_1163), .Y(n_1161) );
OAI22xp33_ASAP7_75t_L g1181 ( .A1(n_1156), .A2(n_1182), .B1(n_1183), .B2(n_1184), .Y(n_1181) );
BUFx3_ASAP7_75t_L g1206 ( .A(n_1156), .Y(n_1206) );
BUFx6f_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
HB1xp67_ASAP7_75t_L g1184 ( .A(n_1159), .Y(n_1184) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1159), .Y(n_1209) );
INVx2_ASAP7_75t_L g1167 ( .A(n_1160), .Y(n_1167) );
NOR2xp33_ASAP7_75t_L g1323 ( .A(n_1164), .B(n_1230), .Y(n_1323) );
OR2x2_ASAP7_75t_L g1164 ( .A(n_1165), .B(n_1168), .Y(n_1164) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
NAND2xp5_ASAP7_75t_L g1255 ( .A(n_1166), .B(n_1256), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1166), .B(n_1271), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1167), .B(n_1190), .Y(n_1189) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1167), .B(n_1168), .Y(n_1199) );
INVx2_ASAP7_75t_L g1301 ( .A(n_1167), .Y(n_1301) );
OAI322xp33_ASAP7_75t_L g1315 ( .A1(n_1167), .A2(n_1192), .A3(n_1199), .B1(n_1223), .B2(n_1316), .C1(n_1318), .C2(n_1319), .Y(n_1315) );
OR2x2_ASAP7_75t_L g1211 ( .A(n_1168), .B(n_1212), .Y(n_1211) );
OR2x2_ASAP7_75t_L g1233 ( .A(n_1168), .B(n_1224), .Y(n_1233) );
BUFx3_ASAP7_75t_L g1168 ( .A(n_1169), .Y(n_1168) );
INVx2_ASAP7_75t_L g1190 ( .A(n_1169), .Y(n_1190) );
AOI222xp33_ASAP7_75t_L g1239 ( .A1(n_1169), .A2(n_1194), .B1(n_1219), .B2(n_1240), .C1(n_1241), .C2(n_1243), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1169), .B(n_1217), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1169), .B(n_1244), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1171), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1172 ( .A(n_1173), .B(n_1178), .Y(n_1172) );
AOI22xp5_ASAP7_75t_L g1214 ( .A1(n_1173), .A2(n_1215), .B1(n_1218), .B2(n_1220), .Y(n_1214) );
A2O1A1Ixp33_ASAP7_75t_L g1253 ( .A1(n_1173), .A2(n_1254), .B(n_1257), .C(n_1263), .Y(n_1253) );
OR2x2_ASAP7_75t_L g1290 ( .A(n_1173), .B(n_1179), .Y(n_1290) );
OR2x2_ASAP7_75t_L g1309 ( .A(n_1173), .B(n_1310), .Y(n_1309) );
INVx3_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
NOR2xp33_ASAP7_75t_L g1210 ( .A(n_1174), .B(n_1211), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1174), .B(n_1193), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1174), .B(n_1231), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1174), .B(n_1252), .Y(n_1251) );
CKINVDCx5p33_ASAP7_75t_R g1174 ( .A(n_1175), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1175), .B(n_1194), .Y(n_1219) );
INVx1_ASAP7_75t_SL g1237 ( .A(n_1175), .Y(n_1237) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1175), .Y(n_1277) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1175), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1175), .B(n_1193), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1177), .Y(n_1175) );
OR2x2_ASAP7_75t_L g1192 ( .A(n_1178), .B(n_1193), .Y(n_1192) );
AND2x4_ASAP7_75t_SL g1231 ( .A(n_1178), .B(n_1193), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1178), .B(n_1194), .Y(n_1282) );
INVx2_ASAP7_75t_SL g1178 ( .A(n_1179), .Y(n_1178) );
INVx2_ASAP7_75t_L g1187 ( .A(n_1179), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1179), .B(n_1193), .Y(n_1263) );
AOI221xp5_ASAP7_75t_L g1185 ( .A1(n_1186), .A2(n_1189), .B1(n_1191), .B2(n_1198), .C(n_1200), .Y(n_1185) );
NOR2xp33_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1188), .Y(n_1186) );
OAI211xp5_ASAP7_75t_SL g1213 ( .A1(n_1187), .A2(n_1214), .B(n_1225), .C(n_1239), .Y(n_1213) );
INVx2_ASAP7_75t_L g1242 ( .A(n_1187), .Y(n_1242) );
INVx2_ASAP7_75t_L g1249 ( .A(n_1187), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1187), .B(n_1201), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1187), .B(n_1219), .Y(n_1306) );
O2A1O1Ixp33_ASAP7_75t_L g1307 ( .A1(n_1187), .A2(n_1308), .B(n_1311), .C(n_1312), .Y(n_1307) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1188), .Y(n_1286) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1189), .Y(n_1321) );
NAND2xp5_ASAP7_75t_L g1216 ( .A(n_1190), .B(n_1217), .Y(n_1216) );
NOR2x1_ASAP7_75t_L g1223 ( .A(n_1190), .B(n_1224), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1190), .B(n_1244), .Y(n_1243) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1193), .B(n_1258), .Y(n_1297) );
CKINVDCx6p67_ASAP7_75t_R g1193 ( .A(n_1194), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1194), .B(n_1237), .Y(n_1236) );
OR2x6_ASAP7_75t_L g1194 ( .A(n_1195), .B(n_1197), .Y(n_1194) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
BUFx3_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
OAI31xp33_ASAP7_75t_L g1265 ( .A1(n_1201), .A2(n_1266), .A3(n_1275), .B(n_1287), .Y(n_1265) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
OAI22xp33_ASAP7_75t_L g1204 ( .A1(n_1205), .A2(n_1206), .B1(n_1207), .B2(n_1208), .Y(n_1204) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1211), .Y(n_1311) );
OAI31xp33_ASAP7_75t_SL g1273 ( .A1(n_1215), .A2(n_1268), .A3(n_1270), .B(n_1274), .Y(n_1273) );
OAI21xp5_ASAP7_75t_L g1280 ( .A1(n_1215), .A2(n_1281), .B(n_1282), .Y(n_1280) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1216), .Y(n_1215) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1217), .Y(n_1295) );
OAI22xp5_ASAP7_75t_L g1246 ( .A1(n_1218), .A2(n_1221), .B1(n_1247), .B2(n_1249), .Y(n_1246) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1219), .B(n_1317), .Y(n_1316) );
NOR2xp33_ASAP7_75t_L g1220 ( .A(n_1221), .B(n_1222), .Y(n_1220) );
INVx2_ASAP7_75t_L g1248 ( .A(n_1221), .Y(n_1248) );
AOI22xp5_ASAP7_75t_L g1257 ( .A1(n_1221), .A2(n_1258), .B1(n_1259), .B2(n_1261), .Y(n_1257) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_1221), .B(n_1260), .Y(n_1291) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1224), .Y(n_1250) );
AOI221xp5_ASAP7_75t_L g1225 ( .A1(n_1226), .A2(n_1228), .B1(n_1229), .B2(n_1232), .C(n_1234), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
NAND2xp5_ASAP7_75t_L g1247 ( .A(n_1228), .B(n_1248), .Y(n_1247) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1228), .Y(n_1272) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1231), .Y(n_1303) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
NOR2xp33_ASAP7_75t_L g1234 ( .A(n_1235), .B(n_1238), .Y(n_1234) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1236), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1241 ( .A(n_1236), .B(n_1242), .Y(n_1241) );
OAI21xp5_ASAP7_75t_SL g1313 ( .A1(n_1236), .A2(n_1260), .B(n_1281), .Y(n_1313) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1240), .Y(n_1318) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1241), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1243), .B(n_1248), .Y(n_1252) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1244), .Y(n_1296) );
AOI21xp33_ASAP7_75t_L g1245 ( .A1(n_1246), .A2(n_1250), .B(n_1251), .Y(n_1245) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1262), .Y(n_1261) );
OAI21xp33_ASAP7_75t_L g1283 ( .A1(n_1262), .A2(n_1284), .B(n_1286), .Y(n_1283) );
NAND2xp5_ASAP7_75t_SL g1264 ( .A(n_1265), .B(n_1292), .Y(n_1264) );
A2O1A1Ixp33_ASAP7_75t_L g1266 ( .A1(n_1267), .A2(n_1269), .B(n_1272), .C(n_1273), .Y(n_1266) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
A2O1A1Ixp33_ASAP7_75t_L g1312 ( .A1(n_1272), .A2(n_1278), .B(n_1310), .C(n_1313), .Y(n_1312) );
OAI211xp5_ASAP7_75t_SL g1275 ( .A1(n_1276), .A2(n_1278), .B(n_1280), .C(n_1283), .Y(n_1275) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1282), .B(n_1285), .Y(n_1284) );
AOI21xp33_ASAP7_75t_L g1287 ( .A1(n_1288), .A2(n_1290), .B(n_1291), .Y(n_1287) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
AOI32xp33_ASAP7_75t_L g1292 ( .A1(n_1293), .A2(n_1297), .A3(n_1298), .B1(n_1299), .B2(n_1301), .Y(n_1292) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
NAND2xp5_ASAP7_75t_L g1294 ( .A(n_1295), .B(n_1296), .Y(n_1294) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
OAI211xp5_ASAP7_75t_SL g1302 ( .A1(n_1303), .A2(n_1304), .B(n_1307), .C(n_1314), .Y(n_1302) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1306), .Y(n_1322) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1309), .Y(n_1308) );
NOR3xp33_ASAP7_75t_L g1314 ( .A(n_1315), .B(n_1320), .C(n_1323), .Y(n_1314) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1328), .B(n_1354), .Y(n_1327) );
NOR3xp33_ASAP7_75t_L g1328 ( .A(n_1329), .B(n_1336), .C(n_1338), .Y(n_1328) );
NAND2xp5_ASAP7_75t_L g1329 ( .A(n_1330), .B(n_1333), .Y(n_1329) );
AOI31xp33_ASAP7_75t_L g1356 ( .A1(n_1357), .A2(n_1362), .A3(n_1367), .B(n_1368), .Y(n_1356) );
BUFx2_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
INVxp67_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1376), .Y(n_1419) );
HB1xp67_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
NAND2xp5_ASAP7_75t_L g1378 ( .A(n_1379), .B(n_1396), .Y(n_1378) );
NAND3xp33_ASAP7_75t_L g1380 ( .A(n_1381), .B(n_1387), .C(n_1392), .Y(n_1380) );
NOR3xp33_ASAP7_75t_L g1396 ( .A(n_1397), .B(n_1404), .C(n_1406), .Y(n_1396) );
NAND2xp5_ASAP7_75t_L g1397 ( .A(n_1398), .B(n_1401), .Y(n_1397) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1421), .Y(n_1420) );
CKINVDCx5p33_ASAP7_75t_R g1421 ( .A(n_1422), .Y(n_1421) );
A2O1A1Ixp33_ASAP7_75t_L g1424 ( .A1(n_1423), .A2(n_1425), .B(n_1427), .C(n_1429), .Y(n_1424) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
endmodule