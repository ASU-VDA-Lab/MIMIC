module fake_aes_10416_n_647 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_647);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_647;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g87 ( .A(n_51), .Y(n_87) );
CKINVDCx16_ASAP7_75t_R g88 ( .A(n_67), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_19), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_13), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_27), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_66), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_25), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_2), .Y(n_94) );
INVxp67_ASAP7_75t_L g95 ( .A(n_12), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_82), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_24), .Y(n_97) );
HB1xp67_ASAP7_75t_L g98 ( .A(n_69), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_59), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_84), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_56), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_55), .Y(n_102) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_33), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_3), .Y(n_104) );
OR2x2_ASAP7_75t_L g105 ( .A(n_48), .B(n_37), .Y(n_105) );
CKINVDCx14_ASAP7_75t_R g106 ( .A(n_64), .Y(n_106) );
BUFx10_ASAP7_75t_L g107 ( .A(n_32), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_18), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_63), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_31), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_2), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_72), .Y(n_112) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_46), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_26), .Y(n_114) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_57), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_61), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_15), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_68), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_70), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_83), .Y(n_120) );
INVx1_ASAP7_75t_SL g121 ( .A(n_76), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_36), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_8), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_58), .Y(n_124) );
INVx1_ASAP7_75t_SL g125 ( .A(n_74), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_20), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_7), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_77), .Y(n_128) );
INVxp67_ASAP7_75t_SL g129 ( .A(n_45), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_43), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_87), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_111), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_98), .B(n_0), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_115), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_91), .B(n_0), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_107), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_87), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_96), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_96), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_107), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_115), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_97), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_107), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_103), .B(n_1), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_115), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_115), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_97), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_88), .B(n_1), .Y(n_148) );
BUFx3_ASAP7_75t_L g149 ( .A(n_91), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_115), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_118), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_101), .B(n_113), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_118), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_106), .B(n_3), .Y(n_154) );
INVxp33_ASAP7_75t_SL g155 ( .A(n_89), .Y(n_155) );
NOR2x1_ASAP7_75t_L g156 ( .A(n_99), .B(n_4), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_136), .B(n_93), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_136), .B(n_122), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_136), .B(n_123), .Y(n_159) );
NAND3xp33_ASAP7_75t_L g160 ( .A(n_131), .B(n_138), .C(n_147), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_153), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_153), .Y(n_162) );
AND2x6_ASAP7_75t_SL g163 ( .A(n_152), .B(n_90), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_153), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_151), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_151), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_136), .B(n_119), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_136), .B(n_99), .Y(n_168) );
AOI22xp33_ASAP7_75t_L g169 ( .A1(n_135), .A2(n_90), .B1(n_94), .B2(n_104), .Y(n_169) );
OR2x2_ASAP7_75t_L g170 ( .A(n_152), .B(n_133), .Y(n_170) );
AND2x6_ASAP7_75t_L g171 ( .A(n_135), .B(n_100), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_140), .B(n_94), .Y(n_172) );
AND2x6_ASAP7_75t_L g173 ( .A(n_135), .B(n_100), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_155), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_152), .B(n_104), .Y(n_175) );
INVx1_ASAP7_75t_SL g176 ( .A(n_155), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_140), .B(n_126), .Y(n_177) );
OAI21xp33_ASAP7_75t_L g178 ( .A1(n_131), .A2(n_130), .B(n_102), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_151), .Y(n_179) );
INVx2_ASAP7_75t_SL g180 ( .A(n_140), .Y(n_180) );
INVx5_ASAP7_75t_L g181 ( .A(n_135), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_135), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_140), .B(n_143), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_140), .B(n_143), .Y(n_184) );
AND2x4_ASAP7_75t_L g185 ( .A(n_143), .B(n_117), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_143), .B(n_119), .Y(n_186) );
BUFx10_ASAP7_75t_L g187 ( .A(n_135), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_151), .Y(n_188) );
OAI22xp33_ASAP7_75t_L g189 ( .A1(n_176), .A2(n_144), .B1(n_133), .B2(n_148), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_183), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_183), .B(n_143), .Y(n_191) );
INVx2_ASAP7_75t_SL g192 ( .A(n_187), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_165), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_187), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_170), .B(n_159), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_184), .B(n_154), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_172), .Y(n_197) );
BUFx8_ASAP7_75t_L g198 ( .A(n_171), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_170), .A2(n_148), .B1(n_154), .B2(n_144), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_187), .B(n_154), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_172), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_172), .Y(n_202) );
NOR2xp33_ASAP7_75t_R g203 ( .A(n_174), .B(n_132), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_184), .B(n_148), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_184), .B(n_137), .Y(n_205) );
INVx2_ASAP7_75t_SL g206 ( .A(n_184), .Y(n_206) );
INVx2_ASAP7_75t_SL g207 ( .A(n_187), .Y(n_207) );
INVxp67_ASAP7_75t_L g208 ( .A(n_177), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_172), .B(n_137), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_185), .B(n_138), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_163), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_185), .B(n_139), .Y(n_212) );
BUFx8_ASAP7_75t_L g213 ( .A(n_171), .Y(n_213) );
OAI221xp5_ASAP7_75t_L g214 ( .A1(n_169), .A2(n_139), .B1(n_142), .B2(n_147), .C(n_95), .Y(n_214) );
INVxp67_ASAP7_75t_L g215 ( .A(n_175), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_185), .B(n_142), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_185), .Y(n_217) );
BUFx12f_ASAP7_75t_L g218 ( .A(n_163), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_181), .B(n_105), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_171), .B(n_149), .Y(n_220) );
AND2x4_ASAP7_75t_L g221 ( .A(n_175), .B(n_156), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_171), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_180), .A2(n_124), .B(n_112), .Y(n_223) );
NOR2x1_ASAP7_75t_R g224 ( .A(n_157), .B(n_129), .Y(n_224) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_171), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_165), .Y(n_226) );
AND2x6_ASAP7_75t_SL g227 ( .A(n_167), .B(n_132), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_158), .B(n_121), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_181), .B(n_156), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_166), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_219), .A2(n_180), .B(n_182), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_195), .B(n_182), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_208), .A2(n_182), .B(n_160), .C(n_186), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_219), .A2(n_182), .B(n_168), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_193), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_199), .B(n_171), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_193), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_189), .B(n_181), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_226), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_190), .B(n_181), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_230), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_191), .A2(n_160), .B(n_178), .C(n_179), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_204), .B(n_171), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_222), .A2(n_181), .B1(n_92), .B2(n_114), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_197), .Y(n_245) );
INVx3_ASAP7_75t_L g246 ( .A(n_194), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_201), .Y(n_247) );
AND2x4_ASAP7_75t_L g248 ( .A(n_202), .B(n_181), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_198), .Y(n_249) );
AND2x4_ASAP7_75t_SL g250 ( .A(n_194), .B(n_166), .Y(n_250) );
NOR2xp67_ASAP7_75t_R g251 ( .A(n_198), .B(n_179), .Y(n_251) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_194), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_L g253 ( .A1(n_215), .A2(n_178), .B(n_188), .C(n_108), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_217), .Y(n_254) );
INVx4_ASAP7_75t_L g255 ( .A(n_222), .Y(n_255) );
AND2x4_ASAP7_75t_L g256 ( .A(n_221), .B(n_173), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_192), .B(n_188), .Y(n_257) );
BUFx3_ASAP7_75t_L g258 ( .A(n_198), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_206), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_221), .B(n_173), .Y(n_260) );
INVx2_ASAP7_75t_SL g261 ( .A(n_213), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_229), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_203), .Y(n_263) );
BUFx8_ASAP7_75t_L g264 ( .A(n_218), .Y(n_264) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_192), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g266 ( .A1(n_196), .A2(n_173), .B1(n_149), .B2(n_117), .Y(n_266) );
INVx4_ASAP7_75t_L g267 ( .A(n_207), .Y(n_267) );
AND2x4_ASAP7_75t_L g268 ( .A(n_221), .B(n_173), .Y(n_268) );
INVx5_ASAP7_75t_L g269 ( .A(n_207), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_229), .Y(n_270) );
AO21x1_ASAP7_75t_L g271 ( .A1(n_223), .A2(n_134), .B(n_141), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_200), .B(n_173), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g273 ( .A1(n_244), .A2(n_211), .B1(n_218), .B2(n_213), .Y(n_273) );
BUFx2_ASAP7_75t_L g274 ( .A(n_249), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_235), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_256), .B(n_211), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_262), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_262), .Y(n_278) );
A2O1A1Ixp33_ASAP7_75t_L g279 ( .A1(n_233), .A2(n_229), .B(n_216), .C(n_209), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_264), .Y(n_280) );
AO21x2_ASAP7_75t_L g281 ( .A1(n_271), .A2(n_231), .B(n_242), .Y(n_281) );
INVx3_ASAP7_75t_L g282 ( .A(n_267), .Y(n_282) );
OR2x6_ASAP7_75t_L g283 ( .A(n_249), .B(n_225), .Y(n_283) );
OAI21x1_ASAP7_75t_L g284 ( .A1(n_271), .A2(n_220), .B(n_161), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_232), .B(n_200), .Y(n_285) );
AND2x4_ASAP7_75t_L g286 ( .A(n_256), .B(n_205), .Y(n_286) );
OAI21x1_ASAP7_75t_L g287 ( .A1(n_234), .A2(n_161), .B(n_164), .Y(n_287) );
BUFx10_ASAP7_75t_L g288 ( .A(n_250), .Y(n_288) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_236), .A2(n_210), .B1(n_212), .B2(n_214), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g290 ( .A(n_264), .Y(n_290) );
BUFx2_ASAP7_75t_SL g291 ( .A(n_249), .Y(n_291) );
OAI21x1_ASAP7_75t_L g292 ( .A1(n_239), .A2(n_161), .B(n_164), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_256), .A2(n_173), .B1(n_213), .B2(n_203), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_260), .A2(n_173), .B1(n_228), .B2(n_227), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_256), .B(n_127), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_235), .Y(n_296) );
OAI21x1_ASAP7_75t_L g297 ( .A1(n_239), .A2(n_105), .B(n_102), .Y(n_297) );
AND2x4_ASAP7_75t_L g298 ( .A(n_268), .B(n_149), .Y(n_298) );
NOR2xp67_ASAP7_75t_L g299 ( .A(n_263), .B(n_4), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_270), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_237), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_237), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_268), .A2(n_149), .B1(n_127), .B2(n_109), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_258), .Y(n_304) );
OAI21x1_ASAP7_75t_L g305 ( .A1(n_241), .A2(n_109), .B(n_112), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g306 ( .A1(n_241), .A2(n_110), .B1(n_116), .B2(n_130), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_245), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_295), .B(n_263), .Y(n_308) );
AO31x2_ASAP7_75t_L g309 ( .A1(n_279), .A2(n_238), .A3(n_266), .B(n_134), .Y(n_309) );
OAI21xp33_ASAP7_75t_SL g310 ( .A1(n_275), .A2(n_267), .B(n_232), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_294), .B(n_268), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_295), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_288), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_289), .A2(n_270), .B1(n_247), .B2(n_254), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_275), .B(n_268), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_296), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_296), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_280), .B(n_261), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_281), .A2(n_287), .B(n_301), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_290), .A2(n_261), .B1(n_258), .B2(n_259), .Y(n_320) );
OAI211xp5_ASAP7_75t_L g321 ( .A1(n_273), .A2(n_253), .B(n_272), .C(n_259), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_306), .A2(n_254), .B1(n_247), .B2(n_245), .C(n_240), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_307), .Y(n_323) );
OR2x6_ASAP7_75t_L g324 ( .A(n_291), .B(n_258), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_285), .A2(n_240), .B1(n_243), .B2(n_264), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_298), .B(n_240), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_307), .Y(n_327) );
AOI221xp5_ASAP7_75t_L g328 ( .A1(n_303), .A2(n_240), .B1(n_248), .B2(n_153), .C(n_116), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_286), .A2(n_264), .B1(n_252), .B2(n_246), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_301), .B(n_250), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_302), .B(n_250), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_286), .A2(n_252), .B1(n_246), .B2(n_248), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_302), .B(n_248), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_298), .B(n_248), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_277), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_286), .B(n_224), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_316), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_317), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_323), .B(n_278), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_327), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_333), .B(n_281), .Y(n_341) );
BUFx3_ASAP7_75t_L g342 ( .A(n_313), .Y(n_342) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_310), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_309), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_314), .B(n_281), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_333), .B(n_297), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_314), .B(n_297), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_335), .B(n_305), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_312), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_309), .B(n_330), .Y(n_350) );
INVxp67_ASAP7_75t_L g351 ( .A(n_330), .Y(n_351) );
AND2x4_ASAP7_75t_L g352 ( .A(n_324), .B(n_282), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_309), .B(n_331), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_319), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_331), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_309), .Y(n_356) );
INVx4_ASAP7_75t_L g357 ( .A(n_324), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_315), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_324), .B(n_282), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_311), .Y(n_360) );
OR2x2_ASAP7_75t_SL g361 ( .A(n_313), .B(n_290), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_313), .B(n_305), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_313), .B(n_300), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_325), .B(n_298), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_341), .B(n_110), .Y(n_365) );
INVxp67_ASAP7_75t_L g366 ( .A(n_363), .Y(n_366) );
INVx1_ASAP7_75t_SL g367 ( .A(n_361), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_340), .Y(n_368) );
AOI21x1_ASAP7_75t_L g369 ( .A1(n_347), .A2(n_287), .B(n_284), .Y(n_369) );
NAND4xp25_ASAP7_75t_L g370 ( .A(n_364), .B(n_329), .C(n_299), .D(n_325), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_341), .B(n_120), .Y(n_371) );
INVxp67_ASAP7_75t_SL g372 ( .A(n_362), .Y(n_372) );
INVx4_ASAP7_75t_L g373 ( .A(n_357), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_341), .B(n_308), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_360), .B(n_318), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_349), .B(n_329), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_340), .Y(n_377) );
OAI33xp33_ASAP7_75t_L g378 ( .A1(n_349), .A2(n_120), .A3(n_124), .B1(n_128), .B2(n_336), .B3(n_146), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_337), .B(n_326), .Y(n_379) );
OAI33xp33_ASAP7_75t_L g380 ( .A1(n_337), .A2(n_128), .A3(n_150), .B1(n_146), .B2(n_145), .B3(n_141), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_350), .B(n_332), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_364), .A2(n_291), .B1(n_274), .B2(n_304), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_340), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_340), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_350), .B(n_353), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_363), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_338), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_338), .Y(n_388) );
AOI211x1_ASAP7_75t_L g389 ( .A1(n_360), .A2(n_321), .B(n_6), .C(n_7), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_361), .B(n_332), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_348), .Y(n_391) );
AO21x2_ASAP7_75t_L g392 ( .A1(n_345), .A2(n_284), .B(n_292), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_350), .B(n_134), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_348), .Y(n_394) );
BUFx3_ASAP7_75t_L g395 ( .A(n_342), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_361), .B(n_334), .Y(n_396) );
INVx4_ASAP7_75t_L g397 ( .A(n_357), .Y(n_397) );
AND2x4_ASAP7_75t_SL g398 ( .A(n_357), .B(n_288), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_385), .B(n_353), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_385), .B(n_353), .Y(n_400) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_367), .B(n_357), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_391), .B(n_344), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_368), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_386), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_391), .B(n_344), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_368), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_394), .B(n_344), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_394), .B(n_345), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_377), .Y(n_409) );
NAND5xp2_ASAP7_75t_SL g410 ( .A(n_382), .B(n_346), .C(n_320), .D(n_347), .E(n_363), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_381), .B(n_344), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_377), .Y(n_412) );
INVxp67_ASAP7_75t_SL g413 ( .A(n_372), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_374), .B(n_356), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_383), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_383), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_375), .B(n_276), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_381), .B(n_356), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_393), .B(n_356), .Y(n_419) );
INVx1_ASAP7_75t_SL g420 ( .A(n_395), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_384), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_384), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_393), .Y(n_423) );
NOR2x1_ASAP7_75t_L g424 ( .A(n_373), .B(n_357), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_365), .B(n_343), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_373), .B(n_343), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_365), .B(n_347), .Y(n_427) );
INVx1_ASAP7_75t_SL g428 ( .A(n_395), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_374), .B(n_354), .Y(n_429) );
NAND3xp33_ASAP7_75t_L g430 ( .A(n_389), .B(n_362), .C(n_348), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_371), .B(n_346), .Y(n_431) );
INVx6_ASAP7_75t_L g432 ( .A(n_373), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_371), .B(n_346), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_375), .B(n_358), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_366), .B(n_354), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_388), .B(n_387), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_387), .B(n_362), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_369), .B(n_355), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_369), .B(n_355), .Y(n_439) );
INVxp67_ASAP7_75t_L g440 ( .A(n_396), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_379), .B(n_358), .Y(n_441) );
AND2x4_ASAP7_75t_L g442 ( .A(n_397), .B(n_352), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_392), .B(n_358), .Y(n_443) );
BUFx2_ASAP7_75t_SL g444 ( .A(n_397), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_392), .B(n_351), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_392), .B(n_351), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_376), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_436), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_404), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_423), .B(n_390), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_447), .B(n_390), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_399), .B(n_397), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_399), .B(n_396), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_433), .B(n_339), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_400), .B(n_134), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_447), .B(n_370), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_433), .B(n_339), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_431), .B(n_339), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_400), .B(n_342), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_440), .B(n_378), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_413), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_403), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_437), .B(n_352), .Y(n_463) );
NAND4xp25_ASAP7_75t_L g464 ( .A(n_417), .B(n_293), .C(n_328), .D(n_359), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_434), .B(n_380), .Y(n_465) );
NOR2xp33_ASAP7_75t_SL g466 ( .A(n_444), .B(n_342), .Y(n_466) );
INVxp67_ASAP7_75t_L g467 ( .A(n_444), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_403), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_437), .B(n_352), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_411), .B(n_141), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_406), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_406), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_409), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_409), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_427), .B(n_352), .Y(n_475) );
NAND3xp33_ASAP7_75t_SL g476 ( .A(n_420), .B(n_274), .C(n_322), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_412), .Y(n_477) );
NOR2x1_ASAP7_75t_L g478 ( .A(n_424), .B(n_342), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_412), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_429), .B(n_352), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_429), .B(n_359), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g482 ( .A1(n_410), .A2(n_141), .B(n_145), .C(n_146), .Y(n_482) );
NOR2x1_ASAP7_75t_L g483 ( .A(n_424), .B(n_359), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_411), .B(n_145), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_415), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_425), .A2(n_359), .B1(n_398), .B2(n_304), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_415), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_418), .B(n_145), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_427), .B(n_359), .Y(n_489) );
NAND3xp33_ASAP7_75t_SL g490 ( .A(n_420), .B(n_125), .C(n_146), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_416), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_416), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_410), .A2(n_398), .B(n_251), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_421), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_421), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_414), .B(n_5), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_425), .B(n_5), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_418), .B(n_150), .Y(n_498) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_422), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_438), .B(n_150), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_414), .B(n_6), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_422), .Y(n_502) );
BUFx2_ASAP7_75t_L g503 ( .A(n_432), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_441), .B(n_8), .Y(n_504) );
BUFx2_ASAP7_75t_L g505 ( .A(n_432), .Y(n_505) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_490), .A2(n_430), .B(n_426), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_467), .A2(n_432), .B1(n_426), .B2(n_442), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_499), .Y(n_508) );
OAI211xp5_ASAP7_75t_SL g509 ( .A1(n_456), .A2(n_497), .B(n_504), .C(n_449), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_499), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_454), .B(n_408), .Y(n_511) );
NAND3xp33_ASAP7_75t_L g512 ( .A(n_460), .B(n_430), .C(n_438), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_460), .A2(n_426), .B1(n_445), .B2(n_446), .Y(n_513) );
OAI21xp33_ASAP7_75t_L g514 ( .A1(n_453), .A2(n_439), .B(n_408), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_493), .A2(n_426), .B(n_442), .C(n_428), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_455), .B(n_445), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_461), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_461), .Y(n_518) );
AOI32xp33_ASAP7_75t_L g519 ( .A1(n_452), .A2(n_442), .A3(n_428), .B1(n_446), .B2(n_439), .Y(n_519) );
AOI221xp5_ASAP7_75t_L g520 ( .A1(n_448), .A2(n_443), .B1(n_405), .B2(n_402), .C(n_407), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_455), .Y(n_521) );
AOI21xp33_ASAP7_75t_L g522 ( .A1(n_465), .A2(n_496), .B(n_501), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_451), .B(n_443), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_462), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_468), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_453), .B(n_435), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_471), .Y(n_527) );
OAI221xp5_ASAP7_75t_SL g528 ( .A1(n_486), .A2(n_435), .B1(n_419), .B2(n_405), .C(n_407), .Y(n_528) );
INVxp67_ASAP7_75t_L g529 ( .A(n_503), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_457), .B(n_419), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_473), .Y(n_531) );
INVx2_ASAP7_75t_SL g532 ( .A(n_459), .Y(n_532) );
NOR4xp25_ASAP7_75t_L g533 ( .A(n_476), .B(n_401), .C(n_402), .D(n_150), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_500), .Y(n_534) );
O2A1O1Ixp33_ASAP7_75t_L g535 ( .A1(n_465), .A2(n_442), .B(n_283), .C(n_282), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_500), .B(n_432), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_466), .A2(n_251), .B(n_283), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_488), .B(n_153), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_474), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_452), .B(n_153), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_485), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_505), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_480), .A2(n_283), .B1(n_269), .B2(n_246), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_488), .B(n_498), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_487), .Y(n_545) );
AOI31xp33_ASAP7_75t_L g546 ( .A1(n_483), .A2(n_9), .A3(n_10), .B(n_11), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_491), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_492), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_494), .Y(n_549) );
AO22x1_ASAP7_75t_L g550 ( .A1(n_478), .A2(n_153), .B1(n_269), .B2(n_11), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_480), .B(n_153), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_472), .Y(n_552) );
AOI222xp33_ASAP7_75t_L g553 ( .A1(n_502), .A2(n_470), .B1(n_484), .B2(n_498), .C1(n_489), .C2(n_475), .Y(n_553) );
INVxp67_ASAP7_75t_SL g554 ( .A(n_470), .Y(n_554) );
INVxp67_ASAP7_75t_L g555 ( .A(n_484), .Y(n_555) );
NAND3xp33_ASAP7_75t_L g556 ( .A(n_482), .B(n_162), .C(n_283), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_464), .A2(n_288), .B1(n_162), .B2(n_252), .Y(n_557) );
NAND2xp33_ASAP7_75t_SL g558 ( .A(n_507), .B(n_481), .Y(n_558) );
OAI222xp33_ASAP7_75t_L g559 ( .A1(n_519), .A2(n_450), .B1(n_469), .B2(n_463), .C1(n_458), .C2(n_479), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_542), .Y(n_560) );
OAI21xp33_ASAP7_75t_L g561 ( .A1(n_513), .A2(n_495), .B(n_479), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_520), .B(n_495), .Y(n_562) );
A2O1A1Ixp33_ASAP7_75t_L g563 ( .A1(n_535), .A2(n_477), .B(n_472), .C(n_12), .Y(n_563) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_517), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_553), .B(n_477), .Y(n_565) );
OAI221xp5_ASAP7_75t_L g566 ( .A1(n_506), .A2(n_9), .B1(n_10), .B2(n_13), .C(n_14), .Y(n_566) );
OAI221xp5_ASAP7_75t_L g567 ( .A1(n_506), .A2(n_14), .B1(n_15), .B2(n_16), .C(n_17), .Y(n_567) );
OAI321xp33_ASAP7_75t_L g568 ( .A1(n_512), .A2(n_162), .A3(n_17), .B1(n_18), .B2(n_19), .C(n_20), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_518), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_508), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_553), .B(n_16), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_510), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_524), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_514), .B(n_21), .Y(n_574) );
O2A1O1Ixp33_ASAP7_75t_L g575 ( .A1(n_546), .A2(n_509), .B(n_522), .C(n_533), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_526), .B(n_516), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_525), .Y(n_577) );
NOR2x1_ASAP7_75t_L g578 ( .A(n_515), .B(n_546), .Y(n_578) );
NOR3xp33_ASAP7_75t_L g579 ( .A(n_550), .B(n_267), .C(n_255), .Y(n_579) );
NOR3xp33_ASAP7_75t_L g580 ( .A(n_551), .B(n_267), .C(n_255), .Y(n_580) );
NAND2x1_ASAP7_75t_L g581 ( .A(n_532), .B(n_21), .Y(n_581) );
AOI22x1_ASAP7_75t_L g582 ( .A1(n_542), .A2(n_22), .B1(n_255), .B2(n_265), .Y(n_582) );
AOI21xp33_ASAP7_75t_SL g583 ( .A1(n_528), .A2(n_529), .B(n_556), .Y(n_583) );
INVxp67_ASAP7_75t_L g584 ( .A(n_540), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_523), .B(n_22), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_537), .B(n_269), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_527), .Y(n_587) );
INVxp33_ASAP7_75t_L g588 ( .A(n_557), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_552), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_531), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_539), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_541), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_511), .B(n_162), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_564), .Y(n_594) );
BUFx3_ASAP7_75t_L g595 ( .A(n_560), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_565), .B(n_554), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_562), .B(n_549), .Y(n_597) );
OAI21xp5_ASAP7_75t_L g598 ( .A1(n_578), .A2(n_543), .B(n_555), .Y(n_598) );
AOI321xp33_ASAP7_75t_L g599 ( .A1(n_575), .A2(n_521), .A3(n_543), .B1(n_544), .B2(n_536), .C(n_534), .Y(n_599) );
AOI31xp33_ASAP7_75t_L g600 ( .A1(n_583), .A2(n_530), .A3(n_538), .B(n_545), .Y(n_600) );
OAI211xp5_ASAP7_75t_L g601 ( .A1(n_581), .A2(n_548), .B(n_547), .C(n_269), .Y(n_601) );
A2O1A1Ixp33_ASAP7_75t_L g602 ( .A1(n_558), .A2(n_292), .B(n_269), .C(n_252), .Y(n_602) );
OAI221xp5_ASAP7_75t_L g603 ( .A1(n_558), .A2(n_255), .B1(n_162), .B2(n_269), .C(n_252), .Y(n_603) );
OAI221xp5_ASAP7_75t_SL g604 ( .A1(n_563), .A2(n_571), .B1(n_566), .B2(n_567), .C(n_561), .Y(n_604) );
OAI221xp5_ASAP7_75t_L g605 ( .A1(n_563), .A2(n_162), .B1(n_265), .B2(n_257), .C(n_30), .Y(n_605) );
OAI22xp33_ASAP7_75t_SL g606 ( .A1(n_586), .A2(n_23), .B1(n_28), .B2(n_29), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_570), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g608 ( .A1(n_586), .A2(n_34), .B(n_35), .Y(n_608) );
AOI22xp33_ASAP7_75t_SL g609 ( .A1(n_582), .A2(n_265), .B1(n_39), .B2(n_40), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_572), .Y(n_610) );
NOR4xp75_ASAP7_75t_L g611 ( .A(n_574), .B(n_38), .C(n_41), .D(n_42), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_573), .Y(n_612) );
OAI21xp33_ASAP7_75t_SL g613 ( .A1(n_576), .A2(n_44), .B(n_47), .Y(n_613) );
OA22x2_ASAP7_75t_L g614 ( .A1(n_584), .A2(n_49), .B1(n_50), .B2(n_52), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_577), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_595), .B(n_588), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_L g617 ( .A1(n_600), .A2(n_568), .B(n_588), .C(n_585), .Y(n_617) );
OAI22xp5_ASAP7_75t_SL g618 ( .A1(n_598), .A2(n_559), .B1(n_592), .B2(n_591), .Y(n_618) );
O2A1O1Ixp33_ASAP7_75t_L g619 ( .A1(n_604), .A2(n_593), .B(n_569), .C(n_579), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_596), .A2(n_593), .B1(n_580), .B2(n_587), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_612), .Y(n_621) );
AOI211xp5_ASAP7_75t_SL g622 ( .A1(n_604), .A2(n_590), .B(n_589), .C(n_60), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_597), .A2(n_589), .B1(n_265), .B2(n_62), .Y(n_623) );
AO22x2_ASAP7_75t_L g624 ( .A1(n_594), .A2(n_53), .B1(n_54), .B2(n_65), .Y(n_624) );
AOI21xp5_ASAP7_75t_L g625 ( .A1(n_601), .A2(n_265), .B(n_73), .Y(n_625) );
AOI221x1_ASAP7_75t_L g626 ( .A1(n_606), .A2(n_71), .B1(n_75), .B2(n_78), .C(n_79), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_615), .A2(n_80), .B1(n_81), .B2(n_85), .C(n_86), .Y(n_627) );
NOR3xp33_ASAP7_75t_L g628 ( .A(n_618), .B(n_601), .C(n_613), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_616), .B(n_607), .Y(n_629) );
INVx2_ASAP7_75t_SL g630 ( .A(n_621), .Y(n_630) );
CKINVDCx5p33_ASAP7_75t_R g631 ( .A(n_620), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_619), .B(n_599), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_623), .B(n_610), .Y(n_633) );
NOR2x1_ASAP7_75t_L g634 ( .A(n_617), .B(n_608), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_632), .B(n_622), .Y(n_635) );
AND5x1_ASAP7_75t_L g636 ( .A(n_628), .B(n_625), .C(n_627), .D(n_602), .E(n_611), .Y(n_636) );
AND3x4_ASAP7_75t_L g637 ( .A(n_634), .B(n_603), .C(n_624), .Y(n_637) );
OAI221xp5_ASAP7_75t_L g638 ( .A1(n_631), .A2(n_609), .B1(n_605), .B2(n_614), .C(n_624), .Y(n_638) );
NAND2xp33_ASAP7_75t_R g639 ( .A(n_635), .B(n_629), .Y(n_639) );
XNOR2xp5_ASAP7_75t_L g640 ( .A(n_637), .B(n_630), .Y(n_640) );
INVxp67_ASAP7_75t_L g641 ( .A(n_638), .Y(n_641) );
INVx3_ASAP7_75t_L g642 ( .A(n_639), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_641), .Y(n_643) );
AO22x2_ASAP7_75t_L g644 ( .A1(n_642), .A2(n_640), .B1(n_633), .B2(n_626), .Y(n_644) );
OAI21xp5_ASAP7_75t_L g645 ( .A1(n_644), .A2(n_642), .B(n_643), .Y(n_645) );
OR2x2_ASAP7_75t_L g646 ( .A(n_645), .B(n_642), .Y(n_646) );
OAI221xp5_ASAP7_75t_L g647 ( .A1(n_646), .A2(n_642), .B1(n_643), .B2(n_636), .C(n_614), .Y(n_647) );
endmodule