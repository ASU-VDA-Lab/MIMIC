module fake_jpeg_30846_n_222 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_222);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_222;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_4),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

AOI21xp33_ASAP7_75t_L g34 ( 
.A1(n_18),
.A2(n_0),
.B(n_1),
.Y(n_34)
);

OR2x2_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_16),
.Y(n_49)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_1),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_36),
.B(n_41),
.Y(n_73)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_1),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_23),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_44),
.B(n_46),
.Y(n_51)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_2),
.Y(n_46)
);

NOR2x1_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_32),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_25),
.B1(n_27),
.B2(n_31),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_50),
.A2(n_55),
.B1(n_69),
.B2(n_32),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_60),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_21),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_54),
.B(n_33),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_30),
.B1(n_25),
.B2(n_26),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_30),
.C(n_25),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_63),
.C(n_70),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_26),
.B1(n_25),
.B2(n_27),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_66),
.B1(n_55),
.B2(n_56),
.Y(n_87)
);

CKINVDCx12_ASAP7_75t_R g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_37),
.B(n_42),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_17),
.Y(n_76)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_38),
.A2(n_31),
.B1(n_24),
.B2(n_28),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_38),
.A2(n_22),
.B1(n_17),
.B2(n_5),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_35),
.A2(n_24),
.B1(n_22),
.B2(n_29),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_72),
.A2(n_70),
.B1(n_20),
.B2(n_68),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_74),
.B(n_81),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_82),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_51),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_84),
.Y(n_113)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_33),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_22),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_87),
.B1(n_64),
.B2(n_48),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_21),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_86),
.B(n_90),
.Y(n_127)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_49),
.B(n_29),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_91),
.A2(n_62),
.B1(n_48),
.B2(n_71),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_57),
.B(n_20),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_95),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_14),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_72),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_98),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_63),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_12),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_10),
.Y(n_118)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_104),
.A2(n_94),
.B1(n_101),
.B2(n_102),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

BUFx24_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_107),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_103),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_2),
.B(n_3),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_124),
.B(n_78),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_118),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_13),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_121),
.Y(n_128)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_3),
.B(n_5),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_108),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_108),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_136),
.A2(n_147),
.B(n_109),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_96),
.B(n_85),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_137),
.A2(n_116),
.B(n_104),
.Y(n_155)
);

CKINVDCx12_ASAP7_75t_R g138 ( 
.A(n_106),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_138),
.Y(n_159)
);

NOR4xp25_ASAP7_75t_SL g141 ( 
.A(n_116),
.B(n_96),
.C(n_82),
.D(n_93),
.Y(n_141)
);

AOI221xp5_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_128),
.B1(n_130),
.B2(n_133),
.C(n_150),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_88),
.B1(n_83),
.B2(n_93),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_145),
.Y(n_167)
);

AND2x6_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_113),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_144),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_124),
.A2(n_103),
.B1(n_79),
.B2(n_100),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_79),
.C(n_77),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_150),
.C(n_109),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_3),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_136),
.B(n_117),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_151),
.B(n_152),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_130),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_114),
.B(n_119),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_158),
.Y(n_170)
);

OAI321xp33_ASAP7_75t_L g157 ( 
.A1(n_143),
.A2(n_127),
.A3(n_120),
.B1(n_123),
.B2(n_114),
.C(n_119),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_161),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_130),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_162),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_107),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_140),
.C(n_122),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_165),
.Y(n_180)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_163),
.B(n_159),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_175),
.Y(n_190)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_166),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_160),
.A2(n_147),
.B1(n_145),
.B2(n_142),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_177),
.A2(n_182),
.B1(n_167),
.B2(n_152),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_131),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_181),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_153),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_160),
.A2(n_147),
.B1(n_132),
.B2(n_139),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_161),
.C(n_165),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_164),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_178),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_172),
.B(n_157),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_187),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_186),
.A2(n_176),
.B1(n_177),
.B2(n_182),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_172),
.B(n_162),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_191),
.C(n_151),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_170),
.C(n_180),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_180),
.A2(n_168),
.B1(n_153),
.B2(n_139),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_193),
.A2(n_175),
.B1(n_167),
.B2(n_140),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_155),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_174),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_195),
.B(n_199),
.Y(n_206)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_189),
.A2(n_176),
.B1(n_173),
.B2(n_169),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_198),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_184),
.B(n_156),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_202),
.C(n_203),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_122),
.C(n_111),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_201),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_209),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_203),
.A2(n_191),
.B(n_190),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_207),
.A2(n_193),
.B1(n_192),
.B2(n_202),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_211),
.A2(n_212),
.B(n_6),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_205),
.A2(n_195),
.B(n_199),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_204),
.A2(n_111),
.B1(n_126),
.B2(n_9),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_213),
.B(n_214),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_208),
.B(n_6),
.Y(n_214)
);

OAI21x1_ASAP7_75t_SL g215 ( 
.A1(n_211),
.A2(n_206),
.B(n_8),
.Y(n_215)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_8),
.Y(n_218)
);

NOR3xp33_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_216),
.C(n_9),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_219),
.C(n_210),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_8),
.Y(n_222)
);


endmodule