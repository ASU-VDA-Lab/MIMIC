module fake_jpeg_309_n_58 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

BUFx10_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx8_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_5),
.B(n_6),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_1),
.B(n_6),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_5),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_5),
.B(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_12),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_0),
.Y(n_20)
);

A2O1A1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_11),
.A2(n_0),
.B(n_1),
.C(n_3),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_21),
.A2(n_15),
.B(n_8),
.Y(n_31)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_25),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_16),
.Y(n_25)
);

AOI21xp33_ASAP7_75t_L g26 ( 
.A1(n_8),
.A2(n_4),
.B(n_10),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_8),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_23),
.A2(n_10),
.B1(n_9),
.B2(n_13),
.Y(n_27)
);

AO221x1_ASAP7_75t_L g43 ( 
.A1(n_27),
.A2(n_29),
.B1(n_9),
.B2(n_13),
.C(n_22),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_25),
.A2(n_20),
.B(n_21),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_33),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_19),
.A2(n_15),
.B(n_8),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_22),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_17),
.A2(n_9),
.B1(n_13),
.B2(n_18),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_38),
.A2(n_17),
.B1(n_18),
.B2(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

NAND3xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_41),
.C(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

XNOR2x1_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_44),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_47),
.B(n_38),
.Y(n_53)
);

OAI321xp33_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_31),
.A3(n_33),
.B1(n_29),
.B2(n_32),
.C(n_30),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_34),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_44),
.C(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_52),
.Y(n_54)
);

BUFx24_ASAP7_75t_SL g51 ( 
.A(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_53),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_36),
.C(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_49),
.Y(n_57)
);

OAI321xp33_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_42),
.A3(n_54),
.B1(n_55),
.B2(n_56),
.C(n_49),
.Y(n_58)
);


endmodule