module fake_jpeg_30944_n_291 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_291);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_291;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_152;
wire n_73;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_265;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_10),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_6),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_7),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_47),
.Y(n_51)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_25),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_20),
.B1(n_23),
.B2(n_32),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_52),
.A2(n_65),
.B1(n_67),
.B2(n_78),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_47),
.Y(n_53)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_32),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_60),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_35),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_61),
.Y(n_127)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_35),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_64),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_23),
.B1(n_31),
.B2(n_27),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_38),
.B1(n_49),
.B2(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_42),
.B(n_26),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_26),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_75),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_23),
.C(n_20),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_93),
.C(n_96),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_29),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_30),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_44),
.A2(n_31),
.B1(n_27),
.B2(n_34),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_41),
.B(n_25),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_84),
.Y(n_107)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_29),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_45),
.Y(n_85)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_36),
.B(n_30),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_88),
.Y(n_123)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_36),
.B(n_33),
.Y(n_90)
);

BUFx24_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_37),
.A2(n_17),
.B1(n_18),
.B2(n_28),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_15),
.B1(n_89),
.B2(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_36),
.B(n_33),
.Y(n_93)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

AO22x1_ASAP7_75t_L g128 ( 
.A1(n_95),
.A2(n_98),
.B1(n_0),
.B2(n_1),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_37),
.A2(n_28),
.B1(n_17),
.B2(n_18),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_44),
.A2(n_31),
.B1(n_27),
.B2(n_34),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_99),
.B(n_100),
.C(n_0),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_44),
.A2(n_31),
.B1(n_34),
.B2(n_16),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_44),
.A2(n_31),
.B1(n_16),
.B2(n_15),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_105),
.A2(n_116),
.B1(n_100),
.B2(n_65),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_96),
.A2(n_19),
.B1(n_25),
.B2(n_8),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_108),
.A2(n_117),
.B1(n_94),
.B2(n_70),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_57),
.A2(n_19),
.B1(n_25),
.B2(n_8),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_55),
.A2(n_19),
.B1(n_25),
.B2(n_9),
.Y(n_117)
);

AO21x1_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_128),
.B(n_82),
.Y(n_148)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_132),
.A2(n_138),
.B1(n_148),
.B2(n_160),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_51),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_71),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_137),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_54),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_142),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_72),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_102),
.A2(n_97),
.B1(n_78),
.B2(n_99),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_72),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_139),
.B(n_144),
.Y(n_187)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_63),
.B1(n_58),
.B2(n_55),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_141),
.A2(n_152),
.B1(n_76),
.B2(n_115),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_123),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_146),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_82),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_107),
.B(n_121),
.C(n_110),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_154),
.C(n_158),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_79),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_125),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_147),
.B(n_157),
.Y(n_185)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_150),
.Y(n_176)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_127),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_153),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_58),
.B1(n_76),
.B2(n_98),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_82),
.Y(n_154)
);

HAxp5_ASAP7_75t_SL g155 ( 
.A(n_128),
.B(n_66),
.CON(n_155),
.SN(n_155)
);

MAJIxp5_ASAP7_75t_SL g191 ( 
.A(n_155),
.B(n_106),
.C(n_3),
.Y(n_191)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_62),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_126),
.A2(n_95),
.B(n_91),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_56),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_159),
.B(n_161),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_103),
.B(n_56),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_103),
.B(n_14),
.Y(n_162)
);

AOI21xp33_ASAP7_75t_L g175 ( 
.A1(n_162),
.A2(n_11),
.B(n_13),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_62),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_163),
.B(n_106),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_119),
.B(n_120),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_165),
.A2(n_2),
.B(n_4),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_137),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_171),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_158),
.A2(n_118),
.B1(n_94),
.B2(n_106),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_170),
.A2(n_191),
.B(n_156),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_103),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_174),
.A2(n_177),
.B1(n_183),
.B2(n_190),
.Y(n_206)
);

AOI322xp5_ASAP7_75t_SL g205 ( 
.A1(n_175),
.A2(n_192),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_134),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_135),
.A2(n_67),
.B1(n_115),
.B2(n_120),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_163),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_186),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_138),
.A2(n_70),
.B1(n_73),
.B2(n_118),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_180),
.A2(n_193),
.B1(n_157),
.B2(n_131),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_148),
.A2(n_73),
.B1(n_106),
.B2(n_11),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_151),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_189),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_139),
.B(n_133),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_148),
.A2(n_144),
.B1(n_142),
.B2(n_145),
.Y(n_190)
);

NAND3xp33_ASAP7_75t_L g192 ( 
.A(n_146),
.B(n_13),
.C(n_14),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_132),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_133),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_197),
.B(n_198),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_154),
.C(n_161),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_204),
.C(n_189),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_169),
.B(n_154),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_207),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_176),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_201),
.B(n_202),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_164),
.B(n_162),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_173),
.C(n_172),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_212),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_130),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_208),
.B(n_209),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_140),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_149),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_210),
.B(n_211),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_150),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_153),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_143),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_209),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_215),
.A2(n_181),
.B(n_164),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_179),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_216),
.A2(n_193),
.B1(n_188),
.B2(n_184),
.Y(n_233)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_217),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_173),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_220),
.C(n_226),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_200),
.A2(n_182),
.B(n_191),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_219),
.B(n_233),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_221),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_222),
.B(n_234),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_179),
.C(n_165),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_186),
.C(n_180),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_232),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_177),
.C(n_166),
.Y(n_232)
);

INVxp33_ASAP7_75t_SL g237 ( 
.A(n_196),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_237),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_230),
.B(n_196),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_244),
.Y(n_255)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_236),
.Y(n_241)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_241),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_225),
.A2(n_206),
.B1(n_200),
.B2(n_208),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_242),
.A2(n_234),
.B1(n_207),
.B2(n_233),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_201),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_198),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_218),
.Y(n_254)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_236),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_250),
.Y(n_259)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_231),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_212),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_251),
.B(n_221),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_254),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_220),
.C(n_226),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_257),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_229),
.C(n_227),
.Y(n_257)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_258),
.Y(n_265)
);

AOI31xp67_ASAP7_75t_L g260 ( 
.A1(n_247),
.A2(n_219),
.A3(n_228),
.B(n_225),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_260),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_249),
.A2(n_206),
.B1(n_227),
.B2(n_235),
.Y(n_261)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_261),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_240),
.B(n_195),
.Y(n_262)
);

BUFx24_ASAP7_75t_SL g270 ( 
.A(n_262),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_260),
.A2(n_242),
.B(n_195),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_211),
.Y(n_275)
);

OA21x2_ASAP7_75t_SL g266 ( 
.A1(n_255),
.A2(n_213),
.B(n_202),
.Y(n_266)
);

OAI221xp5_ASAP7_75t_L g278 ( 
.A1(n_266),
.A2(n_199),
.B1(n_223),
.B2(n_210),
.C(n_259),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_261),
.A2(n_214),
.B(n_206),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_268),
.A2(n_258),
.B(n_257),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_243),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_275),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_276),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_271),
.A2(n_216),
.B1(n_253),
.B2(n_183),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_278),
.B(n_268),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_243),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_263),
.B(n_270),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_277),
.B(n_256),
.Y(n_282)
);

OAI21xp33_ASAP7_75t_L g281 ( 
.A1(n_275),
.A2(n_265),
.B(n_264),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_281),
.B(n_282),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_283),
.A2(n_246),
.B(n_241),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_254),
.C(n_274),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_245),
.C(n_248),
.Y(n_288)
);

NAND3xp33_ASAP7_75t_SL g287 ( 
.A(n_286),
.B(n_166),
.C(n_280),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_287),
.A2(n_288),
.B(n_285),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_250),
.C(n_194),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_176),
.Y(n_291)
);


endmodule