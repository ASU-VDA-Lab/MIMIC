module real_aes_9134_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_720, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_720;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_527;
wire n_434;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g173 ( .A1(n_0), .A2(n_174), .B(n_175), .C(n_179), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_1), .B(n_168), .Y(n_181) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_3), .B(n_153), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_4), .A2(n_142), .B(n_159), .C(n_470), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_5), .A2(n_162), .B(n_491), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_6), .A2(n_162), .B(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_7), .B(n_168), .Y(n_497) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_8), .A2(n_134), .B(n_221), .Y(n_220) );
AND2x6_ASAP7_75t_L g159 ( .A(n_9), .B(n_160), .Y(n_159) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_10), .A2(n_142), .B(n_159), .C(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g462 ( .A(n_11), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_12), .B(n_115), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_12), .B(n_40), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_13), .B(n_178), .Y(n_472) );
INVx1_ASAP7_75t_L g139 ( .A(n_14), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_15), .B(n_153), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_16), .A2(n_154), .B(n_481), .C(n_483), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_17), .B(n_168), .Y(n_484) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_18), .A2(n_66), .B1(n_125), .B2(n_126), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_18), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_19), .B(n_211), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_20), .A2(n_142), .B(n_205), .C(n_210), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g451 ( .A1(n_21), .A2(n_177), .B(n_229), .C(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_22), .B(n_178), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_23), .B(n_178), .Y(n_513) );
CKINVDCx16_ASAP7_75t_R g500 ( .A(n_24), .Y(n_500) );
INVx1_ASAP7_75t_L g512 ( .A(n_25), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_26), .A2(n_142), .B(n_210), .C(n_224), .Y(n_223) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_27), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_28), .Y(n_468) );
INVx1_ASAP7_75t_L g529 ( .A(n_29), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_30), .A2(n_162), .B(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g144 ( .A(n_31), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g188 ( .A1(n_32), .A2(n_157), .B(n_189), .C(n_190), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_33), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_34), .A2(n_177), .B(n_494), .C(n_496), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g122 ( .A1(n_35), .A2(n_123), .B1(n_418), .B2(n_419), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_35), .Y(n_418) );
INVxp67_ASAP7_75t_L g530 ( .A(n_36), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_37), .B(n_226), .Y(n_225) );
CKINVDCx14_ASAP7_75t_R g492 ( .A(n_38), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_39), .A2(n_142), .B(n_210), .C(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g115 ( .A(n_40), .Y(n_115) );
AOI222xp33_ASAP7_75t_L g432 ( .A1(n_41), .A2(n_433), .B1(n_702), .B2(n_703), .C1(n_709), .C2(n_713), .Y(n_432) );
A2O1A1Ixp33_ASAP7_75t_L g459 ( .A1(n_42), .A2(n_179), .B(n_460), .C(n_461), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_43), .B(n_203), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_44), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_45), .B(n_153), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_46), .B(n_162), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_47), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_48), .Y(n_526) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_49), .A2(n_157), .B(n_189), .C(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g176 ( .A(n_50), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_51), .A2(n_704), .B1(n_705), .B2(n_706), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_51), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_52), .A2(n_84), .B1(n_707), .B2(n_708), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_52), .Y(n_708) );
INVx1_ASAP7_75t_L g251 ( .A(n_53), .Y(n_251) );
INVx1_ASAP7_75t_L g450 ( .A(n_54), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_55), .B(n_162), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g214 ( .A(n_56), .Y(n_214) );
CKINVDCx14_ASAP7_75t_R g458 ( .A(n_57), .Y(n_458) );
INVx1_ASAP7_75t_L g160 ( .A(n_58), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_59), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_60), .B(n_168), .Y(n_269) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_61), .A2(n_149), .B(n_209), .C(n_267), .Y(n_266) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_62), .A2(n_104), .B1(n_116), .B2(n_718), .Y(n_103) );
INVx1_ASAP7_75t_L g138 ( .A(n_63), .Y(n_138) );
INVx1_ASAP7_75t_SL g495 ( .A(n_64), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_65), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_66), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_67), .B(n_153), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_68), .B(n_168), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_69), .B(n_154), .Y(n_240) );
INVx1_ASAP7_75t_L g503 ( .A(n_70), .Y(n_503) );
CKINVDCx16_ASAP7_75t_R g171 ( .A(n_71), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_72), .B(n_193), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g141 ( .A1(n_73), .A2(n_142), .B(n_147), .C(n_157), .Y(n_141) );
CKINVDCx16_ASAP7_75t_R g265 ( .A(n_74), .Y(n_265) );
INVx1_ASAP7_75t_L g112 ( .A(n_75), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_76), .A2(n_162), .B(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_77), .B(n_428), .Y(n_427) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_78), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_79), .A2(n_162), .B(n_478), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_80), .A2(n_203), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g479 ( .A(n_81), .Y(n_479) );
CKINVDCx16_ASAP7_75t_R g509 ( .A(n_82), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_83), .B(n_192), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_84), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_85), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_86), .A2(n_162), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g482 ( .A(n_87), .Y(n_482) );
INVx2_ASAP7_75t_L g136 ( .A(n_88), .Y(n_136) );
INVx1_ASAP7_75t_L g471 ( .A(n_89), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_90), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_91), .B(n_178), .Y(n_241) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_92), .B(n_109), .C(n_110), .Y(n_108) );
OR2x2_ASAP7_75t_L g423 ( .A(n_92), .B(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g436 ( .A(n_92), .B(n_425), .Y(n_436) );
INVx2_ASAP7_75t_L g440 ( .A(n_92), .Y(n_440) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_93), .A2(n_142), .B(n_157), .C(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_94), .B(n_162), .Y(n_187) );
INVx1_ASAP7_75t_L g191 ( .A(n_95), .Y(n_191) );
INVxp67_ASAP7_75t_L g268 ( .A(n_96), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_97), .B(n_134), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_98), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g148 ( .A(n_99), .Y(n_148) );
INVx1_ASAP7_75t_L g236 ( .A(n_100), .Y(n_236) );
INVx2_ASAP7_75t_L g453 ( .A(n_101), .Y(n_453) );
AND2x2_ASAP7_75t_L g253 ( .A(n_102), .B(n_196), .Y(n_253) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
BUFx4f_ASAP7_75t_SL g718 ( .A(n_105), .Y(n_718) );
INVx2_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_SL g106 ( .A(n_107), .B(n_113), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g425 ( .A(n_109), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVxp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AO21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_121), .B(n_431), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g717 ( .A(n_119), .Y(n_717) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_420), .B(n_427), .Y(n_121) );
INVx1_ASAP7_75t_L g419 ( .A(n_123), .Y(n_419) );
XNOR2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_127), .Y(n_123) );
INVx2_ASAP7_75t_L g437 ( .A(n_127), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_127), .A2(n_435), .B1(n_711), .B2(n_712), .Y(n_710) );
NAND2x1p5_ASAP7_75t_L g127 ( .A(n_128), .B(n_361), .Y(n_127) );
AND4x1_ASAP7_75t_L g128 ( .A(n_129), .B(n_301), .C(n_316), .D(n_341), .Y(n_128) );
NOR2xp33_ASAP7_75t_SL g129 ( .A(n_130), .B(n_274), .Y(n_129) );
OAI21xp33_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_182), .B(n_254), .Y(n_130) );
AND2x2_ASAP7_75t_L g304 ( .A(n_131), .B(n_200), .Y(n_304) );
AND2x2_ASAP7_75t_L g317 ( .A(n_131), .B(n_199), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_131), .B(n_183), .Y(n_367) );
INVx1_ASAP7_75t_L g371 ( .A(n_131), .Y(n_371) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_167), .Y(n_131) );
INVx2_ASAP7_75t_L g288 ( .A(n_132), .Y(n_288) );
BUFx2_ASAP7_75t_L g315 ( .A(n_132), .Y(n_315) );
AO21x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_140), .B(n_165), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_133), .B(n_166), .Y(n_165) );
INVx3_ASAP7_75t_L g168 ( .A(n_133), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_133), .B(n_198), .Y(n_197) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_133), .A2(n_235), .B(n_242), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_133), .B(n_475), .Y(n_474) );
AO21x2_ASAP7_75t_L g498 ( .A1(n_133), .A2(n_499), .B(n_505), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_133), .B(n_515), .Y(n_514) );
INVx4_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_134), .A2(n_222), .B(n_223), .Y(n_221) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_134), .Y(n_262) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g244 ( .A(n_135), .Y(n_244) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x2_ASAP7_75t_SL g196 ( .A(n_136), .B(n_137), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_161), .Y(n_140) );
INVx5_ASAP7_75t_L g172 ( .A(n_142), .Y(n_172) );
AND2x6_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_143), .Y(n_156) );
BUFx3_ASAP7_75t_L g180 ( .A(n_143), .Y(n_180) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g164 ( .A(n_144), .Y(n_164) );
INVx1_ASAP7_75t_L g230 ( .A(n_144), .Y(n_230) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_146), .Y(n_151) );
INVx3_ASAP7_75t_L g154 ( .A(n_146), .Y(n_154) );
AND2x2_ASAP7_75t_L g163 ( .A(n_146), .B(n_164), .Y(n_163) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_146), .Y(n_178) );
INVx1_ASAP7_75t_L g226 ( .A(n_146), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B(n_152), .C(n_155), .Y(n_147) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_150), .B(n_453), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_150), .B(n_482), .Y(n_481) );
OAI22xp33_ASAP7_75t_L g528 ( .A1(n_150), .A2(n_153), .B1(n_529), .B2(n_530), .Y(n_528) );
INVx4_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g193 ( .A(n_151), .Y(n_193) );
INVx2_ASAP7_75t_L g174 ( .A(n_153), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_153), .B(n_268), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_153), .A2(n_208), .B(n_512), .C(n_513), .Y(n_511) );
INVx5_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_154), .B(n_462), .Y(n_461) );
HB1xp67_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx3_ASAP7_75t_L g496 ( .A(n_156), .Y(n_496) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
O2A1O1Ixp33_ASAP7_75t_SL g170 ( .A1(n_158), .A2(n_171), .B(n_172), .C(n_173), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_L g264 ( .A1(n_158), .A2(n_172), .B(n_265), .C(n_266), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_SL g449 ( .A1(n_158), .A2(n_172), .B(n_450), .C(n_451), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_SL g457 ( .A1(n_158), .A2(n_172), .B(n_458), .C(n_459), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_SL g478 ( .A1(n_158), .A2(n_172), .B(n_479), .C(n_480), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_158), .A2(n_172), .B(n_492), .C(n_493), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_SL g525 ( .A1(n_158), .A2(n_172), .B(n_526), .C(n_527), .Y(n_525) );
INVx4_ASAP7_75t_SL g158 ( .A(n_159), .Y(n_158) );
AND2x4_ASAP7_75t_L g162 ( .A(n_159), .B(n_163), .Y(n_162) );
BUFx3_ASAP7_75t_L g210 ( .A(n_159), .Y(n_210) );
NAND2x1p5_ASAP7_75t_L g237 ( .A(n_159), .B(n_163), .Y(n_237) );
BUFx2_ASAP7_75t_L g203 ( .A(n_162), .Y(n_203) );
INVx1_ASAP7_75t_L g209 ( .A(n_164), .Y(n_209) );
AND2x2_ASAP7_75t_L g255 ( .A(n_167), .B(n_200), .Y(n_255) );
INVx2_ASAP7_75t_L g271 ( .A(n_167), .Y(n_271) );
AND2x2_ASAP7_75t_L g280 ( .A(n_167), .B(n_199), .Y(n_280) );
AND2x2_ASAP7_75t_L g359 ( .A(n_167), .B(n_288), .Y(n_359) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_181), .Y(n_167) );
INVx2_ASAP7_75t_L g189 ( .A(n_172), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_177), .B(n_495), .Y(n_494) );
INVx4_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g460 ( .A(n_178), .Y(n_460) );
INVx2_ASAP7_75t_L g473 ( .A(n_179), .Y(n_473) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_180), .Y(n_195) );
INVx1_ASAP7_75t_L g483 ( .A(n_180), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_216), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_183), .B(n_286), .Y(n_324) );
INVx1_ASAP7_75t_L g412 ( .A(n_183), .Y(n_412) );
AND2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_199), .Y(n_183) );
AND2x2_ASAP7_75t_L g270 ( .A(n_184), .B(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g284 ( .A(n_184), .B(n_285), .Y(n_284) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_184), .Y(n_313) );
OR2x2_ASAP7_75t_L g345 ( .A(n_184), .B(n_287), .Y(n_345) );
AND2x2_ASAP7_75t_L g353 ( .A(n_184), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g386 ( .A(n_184), .B(n_355), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_184), .B(n_255), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_184), .B(n_315), .Y(n_411) );
AND2x2_ASAP7_75t_L g417 ( .A(n_184), .B(n_304), .Y(n_417) );
INVx5_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
BUFx2_ASAP7_75t_L g277 ( .A(n_185), .Y(n_277) );
AND2x2_ASAP7_75t_L g307 ( .A(n_185), .B(n_287), .Y(n_307) );
AND2x2_ASAP7_75t_L g340 ( .A(n_185), .B(n_300), .Y(n_340) );
AND2x2_ASAP7_75t_L g360 ( .A(n_185), .B(n_200), .Y(n_360) );
AND2x2_ASAP7_75t_L g394 ( .A(n_185), .B(n_260), .Y(n_394) );
OR2x6_ASAP7_75t_L g185 ( .A(n_186), .B(n_197), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_196), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_194), .C(n_195), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g250 ( .A1(n_192), .A2(n_195), .B(n_251), .C(n_252), .Y(n_250) );
O2A1O1Ixp5_ASAP7_75t_L g470 ( .A1(n_192), .A2(n_471), .B(n_472), .C(n_473), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g502 ( .A1(n_192), .A2(n_473), .B(n_503), .C(n_504), .Y(n_502) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g212 ( .A(n_196), .Y(n_212) );
INVx1_ASAP7_75t_L g215 ( .A(n_196), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_196), .A2(n_248), .B(n_249), .Y(n_247) );
OA21x2_ASAP7_75t_L g455 ( .A1(n_196), .A2(n_456), .B(n_463), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_196), .A2(n_237), .B(n_509), .C(n_510), .Y(n_508) );
AND2x4_ASAP7_75t_L g300 ( .A(n_199), .B(n_271), .Y(n_300) );
AND2x2_ASAP7_75t_L g311 ( .A(n_199), .B(n_307), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_199), .B(n_287), .Y(n_350) );
INVx2_ASAP7_75t_L g365 ( .A(n_199), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_199), .B(n_299), .Y(n_388) );
AND2x2_ASAP7_75t_L g407 ( .A(n_199), .B(n_359), .Y(n_407) );
INVx5_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_200), .Y(n_306) );
AND2x2_ASAP7_75t_L g314 ( .A(n_200), .B(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g355 ( .A(n_200), .B(n_271), .Y(n_355) );
OR2x6_ASAP7_75t_L g200 ( .A(n_201), .B(n_213), .Y(n_200) );
AOI21xp5_ASAP7_75t_SL g201 ( .A1(n_202), .A2(n_204), .B(n_211), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_208), .Y(n_205) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_209), .B(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_212), .B(n_506), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
AO21x2_ASAP7_75t_L g466 ( .A1(n_215), .A2(n_467), .B(n_474), .Y(n_466) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_218), .B(n_231), .Y(n_217) );
AND2x2_ASAP7_75t_L g278 ( .A(n_218), .B(n_261), .Y(n_278) );
INVx1_ASAP7_75t_SL g218 ( .A(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_219), .B(n_234), .Y(n_258) );
OR2x2_ASAP7_75t_L g291 ( .A(n_219), .B(n_261), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_219), .B(n_261), .Y(n_296) );
AND2x2_ASAP7_75t_L g323 ( .A(n_219), .B(n_260), .Y(n_323) );
AND2x2_ASAP7_75t_L g375 ( .A(n_219), .B(n_233), .Y(n_375) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_220), .B(n_245), .Y(n_283) );
AND2x2_ASAP7_75t_L g319 ( .A(n_220), .B(n_234), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_227), .B(n_228), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_228), .A2(n_240), .B(n_241), .Y(n_239) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx3_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_231), .B(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g309 ( .A(n_232), .B(n_291), .Y(n_309) );
OR2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_245), .Y(n_232) );
OAI322xp33_ASAP7_75t_L g274 ( .A1(n_233), .A2(n_275), .A3(n_279), .B1(n_281), .B2(n_284), .C1(n_289), .C2(n_297), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_233), .B(n_260), .Y(n_282) );
OR2x2_ASAP7_75t_L g292 ( .A(n_233), .B(n_246), .Y(n_292) );
AND2x2_ASAP7_75t_L g294 ( .A(n_233), .B(n_246), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_233), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_233), .B(n_261), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_233), .B(n_390), .Y(n_389) );
INVx5_ASAP7_75t_SL g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_234), .B(n_278), .Y(n_404) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_238), .Y(n_235) );
OAI21xp5_ASAP7_75t_L g467 ( .A1(n_237), .A2(n_468), .B(n_469), .Y(n_467) );
OAI21xp5_ASAP7_75t_L g499 ( .A1(n_237), .A2(n_500), .B(n_501), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
INVx2_ASAP7_75t_L g523 ( .A(n_244), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_245), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g272 ( .A(n_245), .B(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_245), .B(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g334 ( .A(n_245), .B(n_261), .Y(n_334) );
AOI211xp5_ASAP7_75t_SL g362 ( .A1(n_245), .A2(n_363), .B(n_366), .C(n_378), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_245), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g400 ( .A(n_245), .B(n_375), .Y(n_400) );
INVx5_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g328 ( .A(n_246), .B(n_261), .Y(n_328) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_246), .Y(n_337) );
AND2x2_ASAP7_75t_L g377 ( .A(n_246), .B(n_375), .Y(n_377) );
AND2x2_ASAP7_75t_SL g408 ( .A(n_246), .B(n_278), .Y(n_408) );
AND2x2_ASAP7_75t_L g415 ( .A(n_246), .B(n_374), .Y(n_415) );
OR2x6_ASAP7_75t_L g246 ( .A(n_247), .B(n_253), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_256), .B1(n_270), .B2(n_272), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_255), .B(n_277), .Y(n_325) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx1_ASAP7_75t_L g273 ( .A(n_258), .Y(n_273) );
OR2x2_ASAP7_75t_L g333 ( .A(n_258), .B(n_334), .Y(n_333) );
OAI221xp5_ASAP7_75t_SL g381 ( .A1(n_258), .A2(n_382), .B1(n_384), .B2(n_385), .C(n_387), .Y(n_381) );
INVx2_ASAP7_75t_L g320 ( .A(n_259), .Y(n_320) );
AND2x2_ASAP7_75t_L g293 ( .A(n_260), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g383 ( .A(n_260), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_260), .B(n_375), .Y(n_396) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVxp67_ASAP7_75t_L g338 ( .A(n_261), .Y(n_338) );
AND2x2_ASAP7_75t_L g374 ( .A(n_261), .B(n_375), .Y(n_374) );
OA21x2_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_263), .B(n_269), .Y(n_261) );
OA21x2_ASAP7_75t_L g447 ( .A1(n_262), .A2(n_448), .B(n_454), .Y(n_447) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_262), .A2(n_477), .B(n_484), .Y(n_476) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_262), .A2(n_490), .B(n_497), .Y(n_489) );
AND2x2_ASAP7_75t_L g376 ( .A(n_270), .B(n_315), .Y(n_376) );
AND2x2_ASAP7_75t_L g286 ( .A(n_271), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_271), .B(n_344), .Y(n_343) );
NOR2xp33_ASAP7_75t_SL g357 ( .A(n_273), .B(n_320), .Y(n_357) );
INVx1_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g363 ( .A(n_276), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
OR2x2_ASAP7_75t_L g349 ( .A(n_277), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g414 ( .A(n_277), .B(n_359), .Y(n_414) );
INVx2_ASAP7_75t_L g347 ( .A(n_278), .Y(n_347) );
NAND4xp25_ASAP7_75t_SL g410 ( .A(n_279), .B(n_411), .C(n_412), .D(n_413), .Y(n_410) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_280), .B(n_344), .Y(n_379) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_SL g416 ( .A(n_283), .Y(n_416) );
O2A1O1Ixp33_ASAP7_75t_SL g378 ( .A1(n_284), .A2(n_347), .B(n_351), .C(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g373 ( .A(n_286), .B(n_365), .Y(n_373) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_287), .Y(n_299) );
INVx1_ASAP7_75t_L g354 ( .A(n_287), .Y(n_354) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_288), .Y(n_331) );
AOI211xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_292), .B(n_293), .C(n_295), .Y(n_289) );
AND2x2_ASAP7_75t_L g310 ( .A(n_290), .B(n_294), .Y(n_310) );
OAI322xp33_ASAP7_75t_SL g348 ( .A1(n_290), .A2(n_349), .A3(n_351), .B1(n_352), .B2(n_356), .C1(n_357), .C2(n_358), .Y(n_348) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g370 ( .A(n_292), .B(n_296), .Y(n_370) );
INVx1_ASAP7_75t_L g351 ( .A(n_294), .Y(n_351) );
INVx1_ASAP7_75t_SL g369 ( .A(n_296), .Y(n_369) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
AOI222xp33_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_308), .B1(n_310), .B2(n_311), .C1(n_312), .C2(n_720), .Y(n_301) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_303), .B(n_305), .Y(n_302) );
OAI322xp33_ASAP7_75t_L g391 ( .A1(n_303), .A2(n_365), .A3(n_370), .B1(n_392), .B2(n_393), .C1(n_395), .C2(n_396), .Y(n_391) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_304), .A2(n_318), .B1(n_342), .B2(n_346), .C(n_348), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
OAI222xp33_ASAP7_75t_L g321 ( .A1(n_309), .A2(n_322), .B1(n_324), .B2(n_325), .C1(n_326), .C2(n_329), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g387 ( .A1(n_311), .A2(n_318), .B1(n_388), .B2(n_389), .Y(n_387) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
AOI211xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_318), .B(n_321), .C(n_332), .Y(n_316) );
O2A1O1Ixp33_ASAP7_75t_L g397 ( .A1(n_318), .A2(n_355), .B(n_398), .C(n_401), .Y(n_397) );
AND2x4_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AND2x2_ASAP7_75t_L g327 ( .A(n_319), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_SL g390 ( .A(n_323), .Y(n_390) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_330), .B(n_355), .Y(n_384) );
BUFx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AOI21xp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .B(n_339), .Y(n_332) );
OAI221xp5_ASAP7_75t_SL g401 ( .A1(n_333), .A2(n_402), .B1(n_403), .B2(n_404), .C(n_405), .Y(n_401) );
INVxp33_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_337), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_344), .B(n_355), .Y(n_395) );
INVx2_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
AND2x2_ASAP7_75t_L g406 ( .A(n_359), .B(n_365), .Y(n_406) );
AND4x1_ASAP7_75t_L g361 ( .A(n_362), .B(n_380), .C(n_397), .D(n_409), .Y(n_361) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OAI221xp5_ASAP7_75t_SL g366 ( .A1(n_367), .A2(n_368), .B1(n_370), .B2(n_371), .C(n_372), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_374), .B1(n_376), .B2(n_377), .Y(n_372) );
INVx1_ASAP7_75t_L g402 ( .A(n_373), .Y(n_402) );
INVx1_ASAP7_75t_SL g392 ( .A(n_377), .Y(n_392) );
NOR2xp33_ASAP7_75t_SL g380 ( .A(n_381), .B(n_391), .Y(n_380) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_393), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_400), .A2(n_406), .B1(n_407), .B2(n_408), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_415), .B1(n_416), .B2(n_417), .Y(n_409) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx2_ASAP7_75t_L g430 ( .A(n_423), .Y(n_430) );
NOR2x2_ASAP7_75t_L g715 ( .A(n_424), .B(n_440), .Y(n_715) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g439 ( .A(n_425), .B(n_440), .Y(n_439) );
AOI21xp33_ASAP7_75t_L g431 ( .A1(n_427), .A2(n_432), .B(n_716), .Y(n_431) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_437), .B1(n_438), .B2(n_441), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx6_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g711 ( .A(n_439), .Y(n_711) );
BUFx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g712 ( .A(n_442), .Y(n_712) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_628), .Y(n_442) );
NOR4xp25_ASAP7_75t_L g443 ( .A(n_444), .B(n_570), .C(n_600), .D(n_610), .Y(n_443) );
OAI211xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_485), .B(n_533), .C(n_560), .Y(n_444) );
OAI222xp33_ASAP7_75t_L g655 ( .A1(n_445), .A2(n_575), .B1(n_656), .B2(n_657), .C1(n_658), .C2(n_659), .Y(n_655) );
OR2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_464), .Y(n_445) );
AOI33xp33_ASAP7_75t_L g581 ( .A1(n_446), .A2(n_568), .A3(n_569), .B1(n_582), .B2(n_587), .B3(n_589), .Y(n_581) );
OAI211xp5_ASAP7_75t_SL g638 ( .A1(n_446), .A2(n_639), .B(n_641), .C(n_643), .Y(n_638) );
OR2x2_ASAP7_75t_L g654 ( .A(n_446), .B(n_640), .Y(n_654) );
INVx1_ASAP7_75t_L g687 ( .A(n_446), .Y(n_687) );
OR2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_455), .Y(n_446) );
INVx2_ASAP7_75t_L g564 ( .A(n_447), .Y(n_564) );
AND2x2_ASAP7_75t_L g580 ( .A(n_447), .B(n_476), .Y(n_580) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_447), .Y(n_615) );
AND2x2_ASAP7_75t_L g644 ( .A(n_447), .B(n_455), .Y(n_644) );
INVx2_ASAP7_75t_L g544 ( .A(n_455), .Y(n_544) );
BUFx3_ASAP7_75t_L g552 ( .A(n_455), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_455), .B(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g563 ( .A(n_455), .B(n_564), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_455), .B(n_465), .Y(n_592) );
AND2x2_ASAP7_75t_L g661 ( .A(n_455), .B(n_595), .Y(n_661) );
INVx2_ASAP7_75t_SL g555 ( .A(n_464), .Y(n_555) );
OR2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_476), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_465), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g597 ( .A(n_465), .Y(n_597) );
AND2x2_ASAP7_75t_L g608 ( .A(n_465), .B(n_564), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_465), .B(n_593), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_465), .B(n_595), .Y(n_640) );
AND2x2_ASAP7_75t_L g699 ( .A(n_465), .B(n_644), .Y(n_699) );
INVx4_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g569 ( .A(n_466), .B(n_476), .Y(n_569) );
AND2x2_ASAP7_75t_L g579 ( .A(n_466), .B(n_580), .Y(n_579) );
BUFx3_ASAP7_75t_L g601 ( .A(n_466), .Y(n_601) );
AND3x2_ASAP7_75t_L g660 ( .A(n_466), .B(n_661), .C(n_662), .Y(n_660) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_476), .Y(n_551) );
INVx1_ASAP7_75t_SL g595 ( .A(n_476), .Y(n_595) );
NAND3xp33_ASAP7_75t_L g607 ( .A(n_476), .B(n_544), .C(n_608), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_486), .B(n_516), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g630 ( .A1(n_486), .A2(n_579), .B(n_631), .C(n_633), .Y(n_630) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_488), .B(n_507), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_488), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_SL g647 ( .A(n_488), .Y(n_647) );
AND2x2_ASAP7_75t_L g668 ( .A(n_488), .B(n_518), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_488), .B(n_577), .Y(n_696) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_498), .Y(n_488) );
AND2x2_ASAP7_75t_L g541 ( .A(n_489), .B(n_532), .Y(n_541) );
INVx2_ASAP7_75t_L g548 ( .A(n_489), .Y(n_548) );
AND2x2_ASAP7_75t_L g568 ( .A(n_489), .B(n_518), .Y(n_568) );
AND2x2_ASAP7_75t_L g618 ( .A(n_489), .B(n_507), .Y(n_618) );
INVx1_ASAP7_75t_L g622 ( .A(n_489), .Y(n_622) );
INVx2_ASAP7_75t_SL g532 ( .A(n_498), .Y(n_532) );
BUFx2_ASAP7_75t_L g558 ( .A(n_498), .Y(n_558) );
AND2x2_ASAP7_75t_L g685 ( .A(n_498), .B(n_507), .Y(n_685) );
INVx3_ASAP7_75t_SL g518 ( .A(n_507), .Y(n_518) );
AND2x2_ASAP7_75t_L g540 ( .A(n_507), .B(n_541), .Y(n_540) );
AND2x4_ASAP7_75t_L g547 ( .A(n_507), .B(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g577 ( .A(n_507), .B(n_537), .Y(n_577) );
OR2x2_ASAP7_75t_L g586 ( .A(n_507), .B(n_532), .Y(n_586) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_507), .Y(n_604) );
AND2x2_ASAP7_75t_L g609 ( .A(n_507), .B(n_562), .Y(n_609) );
AND2x2_ASAP7_75t_L g637 ( .A(n_507), .B(n_520), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_507), .B(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g675 ( .A(n_507), .B(n_519), .Y(n_675) );
OR2x6_ASAP7_75t_L g507 ( .A(n_508), .B(n_514), .Y(n_507) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
AND2x2_ASAP7_75t_L g599 ( .A(n_518), .B(n_548), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_518), .B(n_541), .Y(n_627) );
AND2x2_ASAP7_75t_L g645 ( .A(n_518), .B(n_562), .Y(n_645) );
OR2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_532), .Y(n_519) );
AND2x2_ASAP7_75t_L g546 ( .A(n_520), .B(n_532), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_520), .B(n_575), .Y(n_574) );
BUFx3_ASAP7_75t_L g584 ( .A(n_520), .Y(n_584) );
OR2x2_ASAP7_75t_L g632 ( .A(n_520), .B(n_552), .Y(n_632) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_524), .B(n_531), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AO21x2_ASAP7_75t_L g537 ( .A1(n_522), .A2(n_538), .B(n_539), .Y(n_537) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g538 ( .A(n_524), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_531), .Y(n_539) );
AND2x2_ASAP7_75t_L g567 ( .A(n_532), .B(n_537), .Y(n_567) );
INVx1_ASAP7_75t_L g575 ( .A(n_532), .Y(n_575) );
AND2x2_ASAP7_75t_L g670 ( .A(n_532), .B(n_548), .Y(n_670) );
AOI222xp33_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_542), .B1(n_545), .B2(n_549), .C1(n_553), .C2(n_556), .Y(n_533) );
INVx1_ASAP7_75t_L g665 ( .A(n_534), .Y(n_665) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_540), .Y(n_534) );
AND2x2_ASAP7_75t_L g561 ( .A(n_535), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g572 ( .A(n_535), .B(n_541), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_535), .B(n_563), .Y(n_588) );
OAI222xp33_ASAP7_75t_L g610 ( .A1(n_535), .A2(n_611), .B1(n_616), .B2(n_617), .C1(n_625), .C2(n_627), .Y(n_610) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g598 ( .A(n_537), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_537), .B(n_618), .Y(n_658) );
AND2x2_ASAP7_75t_L g669 ( .A(n_537), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g677 ( .A(n_540), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_542), .B(n_593), .Y(n_656) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_544), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g614 ( .A(n_544), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
INVx3_ASAP7_75t_L g559 ( .A(n_547), .Y(n_559) );
O2A1O1Ixp33_ASAP7_75t_L g649 ( .A1(n_547), .A2(n_650), .B(n_653), .C(n_655), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_547), .B(n_584), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_547), .B(n_567), .Y(n_689) );
AND2x2_ASAP7_75t_L g562 ( .A(n_548), .B(n_558), .Y(n_562) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
INVx1_ASAP7_75t_L g589 ( .A(n_551), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_552), .B(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g641 ( .A(n_552), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g680 ( .A(n_552), .B(n_580), .Y(n_680) );
INVx1_ASAP7_75t_L g692 ( .A(n_552), .Y(n_692) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_555), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
INVx1_ASAP7_75t_L g673 ( .A(n_558), .Y(n_673) );
A2O1A1Ixp33_ASAP7_75t_SL g560 ( .A1(n_561), .A2(n_563), .B(n_565), .C(n_569), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_561), .A2(n_591), .B1(n_606), .B2(n_609), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_562), .B(n_576), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_562), .B(n_584), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_563), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_SL g626 ( .A(n_563), .Y(n_626) );
AND2x2_ASAP7_75t_L g633 ( .A(n_563), .B(n_613), .Y(n_633) );
INVx2_ASAP7_75t_L g594 ( .A(n_564), .Y(n_594) );
INVxp67_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NOR4xp25_ASAP7_75t_L g571 ( .A(n_568), .B(n_572), .C(n_573), .D(n_576), .Y(n_571) );
INVx1_ASAP7_75t_SL g642 ( .A(n_569), .Y(n_642) );
AND2x2_ASAP7_75t_L g686 ( .A(n_569), .B(n_687), .Y(n_686) );
OAI211xp5_ASAP7_75t_SL g570 ( .A1(n_571), .A2(n_578), .B(n_581), .C(n_590), .Y(n_570) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_577), .B(n_647), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_579), .A2(n_698), .B1(n_699), .B2(n_700), .Y(n_697) );
INVx1_ASAP7_75t_SL g652 ( .A(n_580), .Y(n_652) );
AND2x2_ASAP7_75t_L g691 ( .A(n_580), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_584), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_588), .B(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_589), .B(n_614), .Y(n_674) );
OAI21xp5_ASAP7_75t_SL g590 ( .A1(n_591), .A2(n_596), .B(n_598), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx1_ASAP7_75t_L g666 ( .A(n_593), .Y(n_666) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
INVx2_ASAP7_75t_L g694 ( .A(n_594), .Y(n_694) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_595), .Y(n_621) );
OAI21xp33_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B(n_605), .Y(n_600) );
CKINVDCx16_ASAP7_75t_R g613 ( .A(n_601), .Y(n_613) );
OR2x2_ASAP7_75t_L g651 ( .A(n_601), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AOI21xp33_ASAP7_75t_SL g646 ( .A1(n_604), .A2(n_647), .B(n_648), .Y(n_646) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_608), .A2(n_635), .B1(n_638), .B2(n_645), .C(n_646), .Y(n_634) );
INVx1_ASAP7_75t_SL g678 ( .A(n_609), .Y(n_678) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
OR2x2_ASAP7_75t_L g625 ( .A(n_613), .B(n_626), .Y(n_625) );
INVxp67_ASAP7_75t_L g662 ( .A(n_615), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_619), .B1(n_622), .B2(n_623), .Y(n_617) );
INVx1_ASAP7_75t_L g657 ( .A(n_618), .Y(n_657) );
INVxp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_621), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NOR4xp25_ASAP7_75t_L g628 ( .A(n_629), .B(n_663), .C(n_676), .D(n_688), .Y(n_628) );
NAND3xp33_ASAP7_75t_SL g629 ( .A(n_630), .B(n_634), .C(n_649), .Y(n_629) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_632), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_639), .B(n_644), .Y(n_648) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI221xp5_ASAP7_75t_SL g676 ( .A1(n_651), .A2(n_677), .B1(n_678), .B2(n_679), .C(n_681), .Y(n_676) );
O2A1O1Ixp33_ASAP7_75t_L g667 ( .A1(n_653), .A2(n_668), .B(n_669), .C(n_671), .Y(n_667) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_654), .A2(n_672), .B1(n_674), .B2(n_675), .Y(n_671) );
INVx2_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
A2O1A1Ixp33_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B(n_666), .C(n_667), .Y(n_663) );
INVx1_ASAP7_75t_L g682 ( .A(n_675), .Y(n_682) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OAI21xp5_ASAP7_75t_SL g681 ( .A1(n_682), .A2(n_683), .B(n_686), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
OAI221xp5_ASAP7_75t_SL g688 ( .A1(n_689), .A2(n_690), .B1(n_693), .B2(n_695), .C(n_697), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVxp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVx3_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
endmodule