module fake_jpeg_12391_n_549 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_549);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_549;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_17),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_52),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_55),
.Y(n_126)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_64),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_10),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_65),
.B(n_75),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g156 ( 
.A(n_69),
.Y(n_156)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_73),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_38),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_34),
.B(n_10),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_76),
.B(n_96),
.Y(n_130)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_79),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_85),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_42),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_86),
.A2(n_42),
.B1(n_44),
.B2(n_20),
.Y(n_136)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_87),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_22),
.A2(n_10),
.B(n_2),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_88),
.A2(n_29),
.B(n_30),
.C(n_26),
.Y(n_145)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_32),
.Y(n_139)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_103),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_22),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_105),
.B(n_139),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_53),
.B1(n_100),
.B2(n_91),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_109),
.A2(n_143),
.B1(n_50),
.B2(n_40),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_28),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_110),
.B(n_113),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_82),
.A2(n_42),
.B1(n_35),
.B2(n_33),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_112),
.A2(n_145),
.B(n_155),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_70),
.B(n_43),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_46),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_122),
.B(n_28),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_136),
.A2(n_99),
.B1(n_30),
.B2(n_29),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_54),
.A2(n_50),
.B1(n_40),
.B2(n_44),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_97),
.A2(n_35),
.B1(n_40),
.B2(n_50),
.Y(n_155)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_73),
.Y(n_157)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

AOI21xp33_ASAP7_75t_SL g160 ( 
.A1(n_89),
.A2(n_32),
.B(n_35),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_52),
.Y(n_188)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_95),
.Y(n_164)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_164),
.Y(n_226)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_55),
.Y(n_165)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_156),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_166),
.B(n_194),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_159),
.A2(n_103),
.B1(n_81),
.B2(n_80),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_167),
.A2(n_169),
.B1(n_147),
.B2(n_141),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_115),
.A2(n_81),
.B1(n_80),
.B2(n_59),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_170),
.A2(n_184),
.B1(n_158),
.B2(n_149),
.Y(n_231)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_107),
.Y(n_172)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_173),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_132),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_174),
.Y(n_247)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_175),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_176),
.Y(n_242)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_178),
.Y(n_249)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_179),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_124),
.A2(n_58),
.B1(n_90),
.B2(n_78),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_180),
.A2(n_182),
.B1(n_192),
.B2(n_204),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_128),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_181),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_155),
.A2(n_67),
.B1(n_74),
.B2(n_72),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_154),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_183),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_143),
.A2(n_62),
.B1(n_71),
.B2(n_66),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

AO22x1_ASAP7_75t_SL g186 ( 
.A1(n_150),
.A2(n_96),
.B1(n_69),
.B2(n_26),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_186),
.B(n_59),
.Y(n_228)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_123),
.Y(n_187)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

OAI21xp33_ASAP7_75t_L g261 ( 
.A1(n_188),
.A2(n_199),
.B(n_200),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_112),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_190),
.Y(n_227)
);

BUFx16f_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_130),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_191),
.B(n_210),
.Y(n_239)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_193),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_130),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_111),
.Y(n_195)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_195),
.Y(n_238)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_134),
.Y(n_196)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_196),
.Y(n_241)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_127),
.Y(n_197)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_197),
.Y(n_260)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_117),
.Y(n_198)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_198),
.Y(n_272)
);

AND2x4_ASAP7_75t_SL g199 ( 
.A(n_139),
.B(n_39),
.Y(n_199)
);

NAND2x1_ASAP7_75t_L g200 ( 
.A(n_105),
.B(n_50),
.Y(n_200)
);

OA22x2_ASAP7_75t_L g202 ( 
.A1(n_106),
.A2(n_40),
.B1(n_20),
.B2(n_30),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_202),
.A2(n_20),
.B1(n_149),
.B2(n_147),
.Y(n_229)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_140),
.Y(n_203)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_203),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_124),
.A2(n_41),
.B1(n_48),
.B2(n_47),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_144),
.Y(n_205)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_205),
.Y(n_253)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_148),
.Y(n_207)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_207),
.Y(n_254)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_114),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_153),
.Y(n_209)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_209),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_121),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_108),
.Y(n_211)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_211),
.Y(n_275)
);

BUFx24_ASAP7_75t_L g212 ( 
.A(n_146),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_212),
.Y(n_267)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_142),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_213),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_104),
.A2(n_41),
.B1(n_48),
.B2(n_47),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_214),
.A2(n_222),
.B1(n_225),
.B2(n_182),
.Y(n_248)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_119),
.Y(n_215)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_215),
.Y(n_276)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_120),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_216),
.B(n_218),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_217),
.B(n_224),
.Y(n_269)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_125),
.Y(n_218)
);

BUFx4f_ASAP7_75t_L g219 ( 
.A(n_129),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_219),
.Y(n_262)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_152),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_220),
.B(n_221),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_158),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_116),
.A2(n_21),
.B1(n_46),
.B2(n_43),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_116),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_223),
.B(n_18),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_118),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_118),
.A2(n_21),
.B1(n_29),
.B2(n_26),
.Y(n_225)
);

AOI21x1_ASAP7_75t_L g297 ( 
.A1(n_228),
.A2(n_263),
.B(n_266),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_229),
.A2(n_243),
.B1(n_244),
.B2(n_252),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_231),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_234),
.A2(n_245),
.B1(n_18),
.B2(n_14),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_171),
.B(n_141),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_236),
.B(n_263),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_189),
.A2(n_138),
.B1(n_137),
.B2(n_135),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_204),
.A2(n_138),
.B1(n_137),
.B2(n_135),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_201),
.A2(n_133),
.B1(n_126),
.B2(n_45),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_248),
.B(n_187),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_188),
.A2(n_133),
.B1(n_126),
.B2(n_45),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_171),
.B(n_45),
.C(n_2),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_186),
.C(n_169),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_206),
.A2(n_45),
.B1(n_3),
.B2(n_5),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_258),
.A2(n_13),
.B(n_15),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_199),
.B(n_0),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_199),
.A2(n_45),
.B1(n_3),
.B2(n_5),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_265),
.A2(n_167),
.B1(n_198),
.B2(n_195),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_200),
.B(n_0),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_266),
.B(n_273),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_184),
.A2(n_12),
.B1(n_5),
.B2(n_6),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_268),
.A2(n_262),
.B1(n_255),
.B2(n_276),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_186),
.B(n_0),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_274),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_168),
.B(n_6),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_279),
.B(n_175),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_170),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_280),
.B(n_288),
.C(n_292),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_227),
.B(n_202),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_282),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_284),
.B(n_299),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_237),
.A2(n_248),
.B1(n_228),
.B2(n_273),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_285),
.A2(n_306),
.B1(n_321),
.B2(n_262),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_286),
.B(n_301),
.Y(n_348)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_251),
.Y(n_287)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_287),
.Y(n_329)
);

MAJx2_ASAP7_75t_L g288 ( 
.A(n_239),
.B(n_183),
.C(n_181),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_251),
.Y(n_290)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_290),
.Y(n_332)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_275),
.Y(n_291)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_291),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_236),
.B(n_176),
.C(n_226),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_231),
.A2(n_202),
.B1(n_177),
.B2(n_196),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_293),
.A2(n_302),
.B1(n_305),
.B2(n_307),
.Y(n_339)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_294),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_295),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_296),
.A2(n_312),
.B1(n_328),
.B2(n_257),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_297),
.A2(n_304),
.B(n_317),
.Y(n_347)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_271),
.Y(n_298)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_298),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_269),
.B(n_213),
.Y(n_299)
);

A2O1A1Ixp33_ASAP7_75t_L g300 ( 
.A1(n_256),
.A2(n_212),
.B(n_210),
.C(n_190),
.Y(n_300)
);

NOR3xp33_ASAP7_75t_L g335 ( 
.A(n_300),
.B(n_240),
.C(n_271),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_264),
.B(n_249),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_237),
.A2(n_193),
.B1(n_185),
.B2(n_208),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_230),
.Y(n_303)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_303),
.Y(n_344)
);

AO22x1_ASAP7_75t_L g304 ( 
.A1(n_229),
.A2(n_212),
.B1(n_190),
.B2(n_219),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_252),
.A2(n_219),
.B1(n_7),
.B2(n_9),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_268),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_306)
);

OAI22x1_ASAP7_75t_L g368 ( 
.A1(n_309),
.A2(n_305),
.B1(n_312),
.B2(n_296),
.Y(n_368)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_230),
.Y(n_310)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_310),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_246),
.B(n_13),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_311),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_246),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_249),
.Y(n_313)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_313),
.Y(n_357)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_247),
.Y(n_314)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_314),
.Y(n_363)
);

BUFx2_ASAP7_75t_SL g315 ( 
.A(n_242),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_315),
.Y(n_338)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_270),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_316),
.B(n_319),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_259),
.B(n_258),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_324),
.Y(n_330)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_253),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_253),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_320),
.B(n_322),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_254),
.B(n_13),
.Y(n_322)
);

BUFx12_ASAP7_75t_L g323 ( 
.A(n_257),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_323),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_254),
.B(n_15),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_255),
.B(n_16),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_325),
.B(n_326),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_260),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_276),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_327),
.B(n_277),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_278),
.A2(n_16),
.B1(n_240),
.B2(n_235),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_335),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_297),
.A2(n_233),
.B(n_235),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_336),
.A2(n_350),
.B(n_370),
.Y(n_397)
);

AO22x1_ASAP7_75t_L g342 ( 
.A1(n_285),
.A2(n_241),
.B1(n_233),
.B2(n_232),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_342),
.A2(n_362),
.B(n_364),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_283),
.B(n_260),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_343),
.B(n_346),
.C(n_367),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_345),
.A2(n_314),
.B1(n_316),
.B2(n_290),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_292),
.B(n_267),
.C(n_277),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_282),
.A2(n_241),
.B(n_232),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_282),
.A2(n_238),
.B(n_272),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_351),
.A2(n_352),
.B(n_360),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_286),
.A2(n_238),
.B(n_272),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_328),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_353),
.B(n_303),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_356),
.B(n_351),
.Y(n_401)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_359),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_280),
.A2(n_271),
.B(n_250),
.Y(n_360)
);

OA21x2_ASAP7_75t_L g362 ( 
.A1(n_293),
.A2(n_302),
.B(n_304),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_295),
.A2(n_250),
.B(n_16),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_283),
.B(n_250),
.C(n_16),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_368),
.Y(n_403)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_298),
.Y(n_369)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_369),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_300),
.A2(n_304),
.B(n_317),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_308),
.A2(n_318),
.B1(n_289),
.B2(n_281),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_371),
.A2(n_362),
.B1(n_339),
.B2(n_342),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_349),
.B(n_308),
.Y(n_372)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_372),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_373),
.A2(n_375),
.B1(n_401),
.B2(n_332),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_359),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_374),
.B(n_377),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_345),
.A2(n_325),
.B1(n_324),
.B2(n_287),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_349),
.B(n_291),
.Y(n_376)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_376),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_361),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_313),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_378),
.B(n_380),
.C(n_389),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_350),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_379),
.B(n_385),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_337),
.B(n_288),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_381),
.Y(n_438)
);

AOI322xp5_ASAP7_75t_L g383 ( 
.A1(n_371),
.A2(n_306),
.A3(n_326),
.B1(n_310),
.B2(n_323),
.C1(n_294),
.C2(n_320),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_383),
.B(n_390),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_354),
.Y(n_385)
);

OA22x2_ASAP7_75t_L g387 ( 
.A1(n_362),
.A2(n_319),
.B1(n_327),
.B2(n_323),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_387),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_358),
.A2(n_323),
.B1(n_331),
.B2(n_356),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_388),
.A2(n_393),
.B(n_394),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_348),
.B(n_343),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_354),
.B(n_361),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_365),
.B(n_367),
.Y(n_391)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_391),
.Y(n_426)
);

AOI32xp33_ASAP7_75t_L g393 ( 
.A1(n_336),
.A2(n_330),
.A3(n_352),
.B1(n_360),
.B2(n_370),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_364),
.A2(n_366),
.B1(n_353),
.B2(n_339),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_346),
.B(n_330),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_395),
.B(n_408),
.C(n_340),
.Y(n_428)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_329),
.Y(n_396)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_396),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_398),
.A2(n_368),
.B1(n_341),
.B2(n_357),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_365),
.B(n_363),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_399),
.B(n_400),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_333),
.Y(n_400)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_329),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_402),
.Y(n_437)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_332),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_404),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_368),
.A2(n_342),
.B1(n_362),
.B2(n_344),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_407),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_347),
.B(n_363),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_409),
.A2(n_416),
.B1(n_440),
.B2(n_387),
.Y(n_452)
);

OAI21xp33_ASAP7_75t_L g412 ( 
.A1(n_377),
.A2(n_347),
.B(n_333),
.Y(n_412)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_412),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_403),
.A2(n_401),
.B1(n_375),
.B2(n_397),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_399),
.Y(n_418)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_418),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_378),
.B(n_344),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_419),
.B(n_425),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_376),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_420),
.B(n_422),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_400),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_389),
.B(n_355),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_395),
.B(n_355),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_427),
.B(n_405),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_428),
.B(n_429),
.C(n_406),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_380),
.B(n_392),
.C(n_408),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_384),
.Y(n_430)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_430),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_397),
.A2(n_340),
.B(n_341),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_433),
.B(n_386),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_391),
.B(n_338),
.Y(n_435)
);

CKINVDCx14_ASAP7_75t_R g465 ( 
.A(n_435),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_436),
.A2(n_404),
.B1(n_396),
.B2(n_402),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_392),
.B(n_338),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g455 ( 
.A(n_439),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_403),
.A2(n_401),
.B1(n_382),
.B2(n_374),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_441),
.B(n_443),
.C(n_444),
.Y(n_473)
);

XNOR2x1_ASAP7_75t_SL g442 ( 
.A(n_416),
.B(n_393),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_SL g481 ( 
.A(n_442),
.B(n_453),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_406),
.C(n_372),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_413),
.B(n_382),
.C(n_398),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_413),
.B(n_388),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_446),
.B(n_448),
.Y(n_468)
);

AOI21x1_ASAP7_75t_L g483 ( 
.A1(n_447),
.A2(n_432),
.B(n_431),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_419),
.B(n_394),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_421),
.B(n_426),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_449),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_452),
.A2(n_456),
.B1(n_462),
.B2(n_414),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_423),
.A2(n_386),
.B1(n_405),
.B2(n_387),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_421),
.B(n_387),
.Y(n_457)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_457),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_458),
.A2(n_464),
.B1(n_431),
.B2(n_433),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_428),
.B(n_357),
.C(n_384),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_459),
.B(n_466),
.C(n_438),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_415),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_460),
.B(n_410),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_423),
.A2(n_334),
.B1(n_369),
.B2(n_409),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_417),
.B(n_334),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_463),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_436),
.A2(n_431),
.B1(n_417),
.B2(n_410),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_427),
.B(n_425),
.C(n_426),
.Y(n_466)
);

XNOR2x1_ASAP7_75t_L g467 ( 
.A(n_440),
.B(n_415),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_467),
.B(n_452),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_SL g469 ( 
.A(n_442),
.B(n_432),
.C(n_434),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_469),
.A2(n_468),
.B(n_487),
.Y(n_507)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_471),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_465),
.B(n_424),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_472),
.B(n_474),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_445),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_475),
.B(n_482),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_461),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_476),
.B(n_461),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_477),
.B(n_483),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_454),
.B(n_437),
.Y(n_478)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_478),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_480),
.A2(n_488),
.B1(n_456),
.B2(n_453),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_443),
.B(n_414),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_459),
.B(n_437),
.C(n_430),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_484),
.B(n_489),
.C(n_455),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_485),
.A2(n_450),
.B1(n_463),
.B2(n_467),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_441),
.B(n_411),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_486),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_464),
.A2(n_458),
.B1(n_457),
.B2(n_444),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_466),
.B(n_451),
.C(n_446),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_490),
.A2(n_507),
.B1(n_487),
.B2(n_479),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_SL g517 ( 
.A1(n_491),
.A2(n_494),
.B1(n_499),
.B2(n_492),
.Y(n_517)
);

MAJx2_ASAP7_75t_L g493 ( 
.A(n_473),
.B(n_448),
.C(n_451),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_493),
.B(n_496),
.Y(n_516)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_495),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_489),
.B(n_462),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_498),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_477),
.B(n_485),
.Y(n_499)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_499),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_470),
.B(n_478),
.Y(n_500)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_500),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_474),
.B(n_473),
.C(n_484),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_502),
.B(n_498),
.C(n_496),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_470),
.B(n_479),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_504),
.B(n_481),
.Y(n_514)
);

XNOR2x1_ASAP7_75t_SL g506 ( 
.A(n_481),
.B(n_488),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_SL g521 ( 
.A(n_506),
.B(n_492),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_511),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_490),
.A2(n_480),
.B1(n_483),
.B2(n_469),
.Y(n_512)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_512),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_505),
.B(n_468),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_513),
.B(n_520),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g528 ( 
.A1(n_514),
.A2(n_503),
.B(n_491),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_504),
.A2(n_476),
.B1(n_494),
.B2(n_500),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_515),
.B(n_517),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_518),
.B(n_499),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_502),
.B(n_497),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_521),
.B(n_506),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_521),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_525),
.B(n_528),
.Y(n_533)
);

OAI21xp33_ASAP7_75t_L g527 ( 
.A1(n_514),
.A2(n_507),
.B(n_501),
.Y(n_527)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_527),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_518),
.A2(n_495),
.B(n_493),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_529),
.A2(n_530),
.B(n_512),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_508),
.A2(n_516),
.B(n_519),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_523),
.B(n_515),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_532),
.B(n_535),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_522),
.B(n_516),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_534),
.B(n_510),
.Y(n_538)
);

MAJx2_ASAP7_75t_L g540 ( 
.A(n_536),
.B(n_527),
.C(n_511),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_538),
.B(n_539),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_533),
.B(n_537),
.C(n_526),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_540),
.B(n_532),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_542),
.B(n_541),
.C(n_531),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_544),
.B(n_545),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_542),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_546),
.B(n_543),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_547),
.B(n_531),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_548),
.B(n_509),
.Y(n_549)
);


endmodule