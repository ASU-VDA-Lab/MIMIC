module fake_jpeg_823_n_440 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_440);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_440;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_67),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_20),
.B(n_8),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_46),
.B(n_47),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_31),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_17),
.A2(n_8),
.B1(n_15),
.B2(n_2),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_49),
.A2(n_23),
.B1(n_38),
.B2(n_39),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_50),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_51),
.Y(n_124)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_52),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_34),
.Y(n_54)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_62),
.B(n_70),
.Y(n_121)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_63),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_23),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_20),
.B(n_8),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_77),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_27),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_73),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_27),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_28),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_82),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_28),
.B(n_10),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_32),
.Y(n_82)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_86),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_32),
.B(n_10),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_87),
.B(n_23),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_88),
.B(n_134),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_21),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_94),
.B(n_110),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_49),
.A2(n_37),
.B1(n_40),
.B2(n_36),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_95),
.A2(n_98),
.B1(n_107),
.B2(n_128),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_L g96 ( 
.A1(n_46),
.A2(n_33),
.B(n_29),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_96),
.B(n_129),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_58),
.A2(n_37),
.B1(n_40),
.B2(n_36),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_100),
.A2(n_137),
.B1(n_70),
.B2(n_26),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_60),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_54),
.A2(n_25),
.B1(n_39),
.B2(n_33),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_108),
.A2(n_127),
.B1(n_83),
.B2(n_57),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_33),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_80),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_122),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_54),
.A2(n_25),
.B1(n_30),
.B2(n_29),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_72),
.A2(n_30),
.B1(n_29),
.B2(n_26),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_73),
.B(n_24),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_75),
.B(n_24),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_82),
.A2(n_30),
.B1(n_26),
.B2(n_24),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_92),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_138),
.B(n_149),
.Y(n_216)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_140),
.Y(n_205)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_141),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_142),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_90),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_143),
.B(n_148),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_147),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_99),
.B(n_44),
.Y(n_149)
);

NAND2xp33_ASAP7_75t_SL g203 ( 
.A(n_150),
.B(n_175),
.Y(n_203)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_117),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_153),
.B(n_155),
.Y(n_210)
);

NOR2xp67_ASAP7_75t_L g155 ( 
.A(n_89),
.B(n_79),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_51),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_156),
.Y(n_214)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_159),
.Y(n_198)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_160),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_110),
.B(n_47),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_173),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_94),
.A2(n_62),
.B(n_79),
.C(n_41),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_162),
.A2(n_172),
.B(n_59),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_104),
.B(n_56),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_163),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_122),
.A2(n_63),
.B1(n_48),
.B2(n_50),
.Y(n_164)
);

AOI22x1_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_174),
.B1(n_133),
.B2(n_125),
.Y(n_186)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_91),
.Y(n_165)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_115),
.Y(n_166)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_102),
.Y(n_167)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_118),
.Y(n_169)
);

INVx4_ASAP7_75t_SL g200 ( 
.A(n_169),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_170),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_101),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_180),
.Y(n_196)
);

NAND2x1_ASAP7_75t_SL g172 ( 
.A(n_118),
.B(n_52),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_102),
.B(n_86),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_97),
.A2(n_45),
.B1(n_69),
.B2(n_53),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_111),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g176 ( 
.A(n_114),
.B(n_64),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_126),
.C(n_112),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_115),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_177),
.A2(n_178),
.B1(n_181),
.B2(n_124),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_111),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_SL g209 ( 
.A(n_179),
.B(n_135),
.C(n_133),
.Y(n_209)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_103),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_132),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_157),
.A2(n_114),
.B1(n_104),
.B2(n_119),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_183),
.A2(n_177),
.B1(n_166),
.B2(n_144),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_158),
.A2(n_136),
.B1(n_113),
.B2(n_53),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_185),
.A2(n_194),
.B1(n_211),
.B2(n_164),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_186),
.A2(n_106),
.B1(n_119),
.B2(n_120),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_187),
.B(n_202),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_135),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_176),
.C(n_172),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_161),
.A2(n_136),
.B1(n_69),
.B2(n_50),
.Y(n_194)
);

NOR3xp33_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_169),
.C(n_112),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_151),
.A2(n_45),
.B1(n_86),
.B2(n_85),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_150),
.A2(n_126),
.B1(n_124),
.B2(n_123),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

AOI32xp33_ASAP7_75t_L g215 ( 
.A1(n_138),
.A2(n_125),
.A3(n_120),
.B1(n_68),
.B2(n_66),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_152),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_202),
.A2(n_162),
.B(n_172),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_218),
.A2(n_209),
.B(n_206),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_210),
.A2(n_141),
.B(n_146),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_219),
.A2(n_227),
.B(n_233),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_176),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_220),
.B(n_231),
.C(n_196),
.Y(n_259)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_221),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_216),
.B(n_153),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_222),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_223),
.B(n_237),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_196),
.Y(n_224)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_224),
.Y(n_269)
);

XNOR2x1_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_199),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_203),
.A2(n_195),
.B(n_216),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_195),
.A2(n_154),
.B1(n_174),
.B2(n_165),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_228),
.A2(n_249),
.B1(n_198),
.B2(n_193),
.Y(n_256)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_189),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_229),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_214),
.A2(n_145),
.B1(n_167),
.B2(n_123),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_230),
.A2(n_245),
.B1(n_76),
.B2(n_78),
.Y(n_277)
);

MAJx2_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_181),
.C(n_159),
.Y(n_231)
);

NAND3xp33_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_170),
.C(n_148),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_190),
.B(n_160),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_234),
.B(n_239),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_192),
.A2(n_169),
.B(n_180),
.Y(n_235)
);

NAND2xp33_ASAP7_75t_SL g279 ( 
.A(n_235),
.B(n_240),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_236),
.Y(n_273)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_238),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_187),
.B(n_168),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_247),
.B1(n_200),
.B2(n_197),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_139),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_243),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_184),
.Y(n_245)
);

NOR2x1_ASAP7_75t_L g246 ( 
.A(n_186),
.B(n_147),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_248),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_194),
.B(n_140),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_185),
.A2(n_142),
.B1(n_85),
.B2(n_84),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_251),
.A2(n_41),
.B(n_171),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_228),
.A2(n_186),
.B1(n_211),
.B2(n_182),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_252),
.A2(n_253),
.B1(n_258),
.B2(n_268),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_223),
.A2(n_182),
.B1(n_193),
.B2(n_201),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_255),
.A2(n_256),
.B1(n_261),
.B2(n_267),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_257),
.B(n_224),
.C(n_234),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_244),
.A2(n_201),
.B1(n_199),
.B2(n_184),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_259),
.B(n_231),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_218),
.A2(n_197),
.B1(n_188),
.B2(n_196),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_244),
.A2(n_188),
.B(n_198),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_266),
.A2(n_275),
.B(n_226),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_244),
.A2(n_248),
.B1(n_247),
.B2(n_239),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_227),
.A2(n_106),
.B1(n_217),
.B2(n_207),
.Y(n_268)
);

A2O1A1Ixp33_ASAP7_75t_L g270 ( 
.A1(n_225),
.A2(n_208),
.B(n_205),
.C(n_217),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_229),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_220),
.A2(n_208),
.B1(n_205),
.B2(n_61),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_272),
.A2(n_276),
.B1(n_238),
.B2(n_93),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_242),
.A2(n_226),
.B(n_235),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_242),
.A2(n_103),
.B1(n_76),
.B2(n_78),
.Y(n_276)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_277),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_280),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_265),
.B(n_222),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_281),
.B(n_282),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_266),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_258),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_283),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_260),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_284),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_271),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_291),
.C(n_292),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_250),
.B(n_219),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_287),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_268),
.Y(n_288)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_288),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_261),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_290),
.B(n_301),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_221),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_262),
.A2(n_249),
.B1(n_246),
.B2(n_240),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_293),
.A2(n_302),
.B1(n_255),
.B2(n_276),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_298),
.C(n_300),
.Y(n_317)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_296),
.Y(n_316)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_297),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_259),
.B(n_245),
.C(n_236),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_260),
.Y(n_299)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_299),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_245),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_250),
.B(n_236),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_262),
.A2(n_81),
.B1(n_41),
.B2(n_171),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_270),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_278),
.B(n_274),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_306),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_278),
.B(n_171),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_305),
.B(n_303),
.C(n_291),
.Y(n_329)
);

OAI21x1_ASAP7_75t_R g306 ( 
.A1(n_279),
.A2(n_0),
.B(n_1),
.Y(n_306)
);

OA22x2_ASAP7_75t_L g307 ( 
.A1(n_267),
.A2(n_93),
.B1(n_64),
.B2(n_22),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_277),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_294),
.A2(n_262),
.B1(n_264),
.B2(n_252),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_312),
.A2(n_313),
.B1(n_319),
.B2(n_332),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_290),
.A2(n_262),
.B1(n_264),
.B2(n_253),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_315),
.B(n_321),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_286),
.B(n_251),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_318),
.B(n_300),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_297),
.A2(n_256),
.B1(n_270),
.B2(n_275),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_285),
.A2(n_272),
.B1(n_269),
.B2(n_274),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_SL g351 ( 
.A(n_322),
.B(n_328),
.C(n_306),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_285),
.A2(n_269),
.B1(n_279),
.B2(n_273),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_307),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_305),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_301),
.B(n_273),
.Y(n_330)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_330),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_292),
.B(n_254),
.C(n_263),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_307),
.C(n_306),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_293),
.A2(n_254),
.B1(n_263),
.B2(n_64),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_334),
.B(n_337),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_295),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_338),
.B(n_351),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_339),
.B(n_355),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_309),
.B(n_298),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_340),
.B(n_341),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_317),
.B(n_280),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_308),
.Y(n_342)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_342),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_333),
.B(n_299),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_343),
.B(n_352),
.Y(n_358)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_324),
.Y(n_344)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_344),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_302),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_345),
.B(n_349),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_346),
.B(n_356),
.C(n_323),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_314),
.B(n_333),
.Y(n_347)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_347),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_311),
.B(n_326),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_325),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_350),
.B(n_353),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_310),
.B(n_254),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_323),
.A2(n_296),
.B(n_289),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_326),
.B(n_331),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_354),
.B(n_337),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_329),
.B(n_307),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_318),
.B(n_289),
.C(n_93),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_348),
.A2(n_325),
.B1(n_320),
.B2(n_312),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_357),
.A2(n_370),
.B1(n_374),
.B2(n_22),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_SL g388 ( 
.A(n_362),
.B(n_11),
.Y(n_388)
);

BUFx12_ASAP7_75t_L g363 ( 
.A(n_339),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_363),
.B(n_367),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_336),
.A2(n_320),
.B1(n_319),
.B2(n_313),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_366),
.A2(n_335),
.B1(n_353),
.B2(n_351),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_345),
.B(n_310),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_348),
.A2(n_316),
.B1(n_327),
.B2(n_315),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_340),
.B(n_321),
.C(n_330),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_371),
.B(n_372),
.Y(n_386)
);

OAI321xp33_ASAP7_75t_L g374 ( 
.A1(n_336),
.A2(n_316),
.A3(n_328),
.B1(n_324),
.B2(n_322),
.C(n_332),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_373),
.B(n_341),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_376),
.B(n_12),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_375),
.B(n_334),
.C(n_356),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_377),
.B(n_378),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_375),
.B(n_355),
.C(n_346),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_358),
.Y(n_379)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_379),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_380),
.A2(n_364),
.B1(n_363),
.B2(n_3),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_359),
.A2(n_19),
.B(n_22),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_381),
.A2(n_388),
.B(n_389),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_373),
.B(n_0),
.C(n_1),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_383),
.C(n_387),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_371),
.B(n_0),
.C(n_1),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_385),
.A2(n_370),
.B1(n_357),
.B2(n_360),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_362),
.B(n_0),
.C(n_1),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_369),
.A2(n_11),
.B(n_2),
.Y(n_389)
);

AOI21x1_ASAP7_75t_SL g390 ( 
.A1(n_369),
.A2(n_11),
.B(n_2),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_390),
.A2(n_365),
.B1(n_368),
.B2(n_366),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_361),
.B(n_6),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_391),
.B(n_13),
.Y(n_396)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_392),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_395),
.A2(n_4),
.B1(n_5),
.B2(n_13),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_396),
.B(n_4),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_364),
.C(n_363),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_397),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_398),
.B(n_402),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_376),
.B(n_377),
.C(n_386),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_399),
.B(n_405),
.C(n_382),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_400),
.B(n_381),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_380),
.A2(n_5),
.B1(n_2),
.B2(n_3),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_384),
.B(n_13),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_404),
.A2(n_393),
.B(n_405),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_383),
.B(n_1),
.C(n_3),
.Y(n_405)
);

A2O1A1Ixp33_ASAP7_75t_SL g407 ( 
.A1(n_398),
.A2(n_390),
.B(n_389),
.C(n_387),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_410),
.Y(n_422)
);

OAI211xp5_ASAP7_75t_L g408 ( 
.A1(n_401),
.A2(n_395),
.B(n_394),
.C(n_399),
.Y(n_408)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_408),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g424 ( 
.A(n_411),
.B(n_413),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_412),
.B(n_414),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_403),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_415),
.B(n_416),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_397),
.A2(n_4),
.B(n_5),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_409),
.B(n_406),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_418),
.A2(n_419),
.B(n_421),
.Y(n_431)
);

NOR2x1_ASAP7_75t_L g419 ( 
.A(n_417),
.B(n_400),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_406),
.B(n_393),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_420),
.B(n_407),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_407),
.B(n_402),
.Y(n_421)
);

NOR3xp33_ASAP7_75t_L g435 ( 
.A(n_427),
.B(n_428),
.C(n_429),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_424),
.B(n_14),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_423),
.B(n_14),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_418),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_430),
.A2(n_432),
.B(n_14),
.Y(n_434)
);

A2O1A1Ixp33_ASAP7_75t_SL g432 ( 
.A1(n_422),
.A2(n_421),
.B(n_425),
.C(n_426),
.Y(n_432)
);

NAND4xp25_ASAP7_75t_SL g433 ( 
.A(n_431),
.B(n_14),
.C(n_15),
.D(n_16),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_433),
.B(n_434),
.Y(n_436)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_435),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_437),
.B(n_16),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_438),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_439),
.B(n_436),
.Y(n_440)
);


endmodule