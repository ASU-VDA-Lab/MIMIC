module fake_ibex_738_n_963 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_168, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_963);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_963;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_418;
wire n_256;
wire n_510;
wire n_193;
wire n_845;
wire n_947;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_909;
wire n_545;
wire n_862;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_375;
wire n_280;
wire n_340;
wire n_317;
wire n_698;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_832;
wire n_798;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_604;
wire n_441;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_490;
wire n_407;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_953;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_960;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_262;
wire n_433;
wire n_299;
wire n_439;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_456;
wire n_368;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_581;
wire n_416;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_200;
wire n_506;
wire n_444;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_520;
wire n_411;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_397;
wire n_366;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_285;
wire n_247;
wire n_379;
wire n_320;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_440;
wire n_268;
wire n_858;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_683;
wire n_631;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_912;
wire n_921;
wire n_677;
wire n_489;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_16),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_62),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_68),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_85),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_44),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_72),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_61),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_79),
.Y(n_181)
);

BUFx2_ASAP7_75t_SL g182 ( 
.A(n_73),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_3),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_161),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_51),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_167),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_137),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_49),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_57),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_1),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_127),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_86),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_132),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_105),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_75),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_50),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_3),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_81),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_143),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_42),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_114),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_4),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_22),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_63),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_7),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_25),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_88),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_24),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_34),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_30),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_152),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_106),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_151),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_46),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_150),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_109),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_123),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_43),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_126),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_145),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_141),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_96),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_53),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_138),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_30),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_31),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_154),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_140),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_70),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_56),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_93),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_18),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_18),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_158),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_25),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_120),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_135),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_131),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_100),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_92),
.B(n_80),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_15),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_8),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_117),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_84),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_32),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_172),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_89),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_107),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_134),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_50),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_44),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_5),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_168),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_64),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_112),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_41),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_99),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_48),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_11),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_22),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_9),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_21),
.Y(n_266)
);

INVxp67_ASAP7_75t_SL g267 ( 
.A(n_1),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_113),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_34),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_43),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_10),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_163),
.Y(n_272)
);

INVxp67_ASAP7_75t_SL g273 ( 
.A(n_6),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_5),
.Y(n_274)
);

INVxp33_ASAP7_75t_L g275 ( 
.A(n_148),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_139),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_67),
.Y(n_277)
);

INVxp67_ASAP7_75t_SL g278 ( 
.A(n_121),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_58),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_24),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_116),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_115),
.Y(n_282)
);

BUFx8_ASAP7_75t_SL g283 ( 
.A(n_103),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_153),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_149),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_60),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_32),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_104),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_101),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_27),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_66),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_111),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_170),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_74),
.Y(n_294)
);

NOR2xp67_ASAP7_75t_L g295 ( 
.A(n_125),
.B(n_155),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_39),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_7),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_133),
.Y(n_298)
);

NOR2xp67_ASAP7_75t_L g299 ( 
.A(n_71),
.B(n_130),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_147),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_97),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_90),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_102),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_136),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_203),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_208),
.B(n_0),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_208),
.B(n_0),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_203),
.Y(n_308)
);

OAI21x1_ASAP7_75t_L g309 ( 
.A1(n_194),
.A2(n_76),
.B(n_164),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_215),
.B(n_2),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_173),
.Y(n_311)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_241),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_283),
.Y(n_313)
);

AND2x4_ASAP7_75t_L g314 ( 
.A(n_215),
.B(n_2),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_202),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_207),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_202),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_204),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_211),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_204),
.Y(n_320)
);

AND2x4_ASAP7_75t_L g321 ( 
.A(n_198),
.B(n_12),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_226),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_231),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_207),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_210),
.Y(n_325)
);

AND2x6_ASAP7_75t_L g326 ( 
.A(n_231),
.B(n_52),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_276),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_227),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_227),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_198),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_173),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_206),
.B(n_14),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_302),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_275),
.B(n_15),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_229),
.B(n_17),
.Y(n_335)
);

AND2x6_ASAP7_75t_L g336 ( 
.A(n_210),
.B(n_54),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_302),
.Y(n_337)
);

AND2x4_ASAP7_75t_L g338 ( 
.A(n_245),
.B(n_19),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_283),
.B(n_55),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_245),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_298),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_298),
.Y(n_342)
);

OAI21x1_ASAP7_75t_L g343 ( 
.A1(n_300),
.A2(n_91),
.B(n_162),
.Y(n_343)
);

NOR2x1_ASAP7_75t_L g344 ( 
.A(n_174),
.B(n_19),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_263),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_236),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_230),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_189),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_247),
.B(n_20),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_241),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_205),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_230),
.B(n_26),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_189),
.B(n_28),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_184),
.B(n_28),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_300),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_249),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_279),
.B(n_29),
.Y(n_357)
);

INVx5_ASAP7_75t_L g358 ( 
.A(n_301),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_303),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_303),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_249),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_304),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_218),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_304),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_218),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_222),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_255),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_249),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_222),
.Y(n_369)
);

OA21x2_ASAP7_75t_L g370 ( 
.A1(n_175),
.A2(n_98),
.B(n_159),
.Y(n_370)
);

INVx6_ASAP7_75t_L g371 ( 
.A(n_301),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_290),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_176),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_179),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_270),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_375)
);

AND2x2_ASAP7_75t_SL g376 ( 
.A(n_180),
.B(n_165),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_186),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_188),
.Y(n_378)
);

NAND2x1p5_ASAP7_75t_L g379 ( 
.A(n_205),
.B(n_59),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_288),
.B(n_33),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_301),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_209),
.B(n_35),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_249),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_287),
.B(n_36),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_190),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_192),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_195),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_196),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_199),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_209),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_287),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_297),
.B(n_37),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_296),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_289),
.B(n_37),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_217),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_297),
.A2(n_185),
.B1(n_181),
.B2(n_292),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_177),
.B(n_38),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_219),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_220),
.Y(n_399)
);

OR2x6_ASAP7_75t_L g400 ( 
.A(n_391),
.B(n_182),
.Y(n_400)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_358),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_353),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_353),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_381),
.B(n_178),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_330),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_381),
.B(n_178),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_353),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_382),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_382),
.Y(n_409)
);

OR2x6_ASAP7_75t_L g410 ( 
.A(n_391),
.B(n_182),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_382),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_330),
.Y(n_412)
);

BUFx10_ASAP7_75t_L g413 ( 
.A(n_371),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_314),
.B(n_212),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_358),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_371),
.B(n_221),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_371),
.B(n_224),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_358),
.B(n_187),
.Y(n_418)
);

NOR2x1p5_ASAP7_75t_L g419 ( 
.A(n_313),
.B(n_267),
.Y(n_419)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_358),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_382),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_371),
.B(n_225),
.Y(n_422)
);

AND2x4_ASAP7_75t_SL g423 ( 
.A(n_367),
.B(n_296),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_340),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_305),
.A2(n_237),
.B1(n_212),
.B2(n_197),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_321),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_350),
.B(n_228),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_314),
.B(n_237),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_314),
.B(n_183),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_340),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_321),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_347),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_390),
.Y(n_433)
);

NAND2xp33_ASAP7_75t_L g434 ( 
.A(n_326),
.B(n_244),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_321),
.Y(n_435)
);

AND3x2_ASAP7_75t_L g436 ( 
.A(n_339),
.B(n_273),
.C(n_278),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_323),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_345),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_313),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_345),
.B(n_296),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_305),
.B(n_232),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_389),
.B(n_373),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_373),
.B(n_233),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_380),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_338),
.Y(n_445)
);

AND3x1_ASAP7_75t_L g446 ( 
.A(n_375),
.B(n_201),
.C(n_191),
.Y(n_446)
);

INVx4_ASAP7_75t_L g447 ( 
.A(n_326),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_323),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_309),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_374),
.B(n_193),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_314),
.B(n_213),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_323),
.Y(n_452)
);

BUFx10_ASAP7_75t_L g453 ( 
.A(n_338),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_327),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_308),
.B(n_238),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_319),
.B(n_193),
.Y(n_456)
);

AND2x6_ASAP7_75t_L g457 ( 
.A(n_338),
.B(n_240),
.Y(n_457)
);

BUFx4f_ASAP7_75t_L g458 ( 
.A(n_376),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_374),
.B(n_200),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_377),
.B(n_388),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_309),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_398),
.B(n_243),
.Y(n_462)
);

AND2x6_ASAP7_75t_L g463 ( 
.A(n_306),
.B(n_248),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_393),
.B(n_239),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_380),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_355),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_306),
.B(n_246),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_394),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_327),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_316),
.B(n_250),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_327),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_327),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_398),
.B(n_251),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_316),
.B(n_252),
.Y(n_474)
);

AND2x6_ASAP7_75t_L g475 ( 
.A(n_394),
.B(n_253),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_324),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_327),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_324),
.B(n_257),
.Y(n_478)
);

INVx6_ASAP7_75t_L g479 ( 
.A(n_312),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_325),
.Y(n_480)
);

BUFx4f_ASAP7_75t_L g481 ( 
.A(n_376),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_335),
.B(n_254),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_325),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_341),
.A2(n_265),
.B1(n_266),
.B2(n_264),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_341),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_312),
.B(n_258),
.Y(n_486)
);

NAND3xp33_ASAP7_75t_L g487 ( 
.A(n_310),
.B(n_274),
.C(n_256),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_342),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_376),
.A2(n_181),
.B1(n_185),
.B2(n_292),
.Y(n_489)
);

OAI22xp33_ASAP7_75t_L g490 ( 
.A1(n_375),
.A2(n_260),
.B1(n_262),
.B2(n_269),
.Y(n_490)
);

BUFx8_ASAP7_75t_SL g491 ( 
.A(n_311),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_342),
.B(n_214),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_312),
.B(n_261),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_332),
.B(n_216),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_332),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_334),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_359),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_359),
.A2(n_280),
.B1(n_271),
.B2(n_294),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_354),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_335),
.B(n_307),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_360),
.B(n_216),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_360),
.B(n_223),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_362),
.B(n_277),
.Y(n_503)
);

AND2x6_ASAP7_75t_L g504 ( 
.A(n_334),
.B(n_281),
.Y(n_504)
);

BUFx4f_ASAP7_75t_L g505 ( 
.A(n_379),
.Y(n_505)
);

AND2x2_ASAP7_75t_SL g506 ( 
.A(n_354),
.B(n_282),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_364),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_364),
.B(n_234),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_357),
.A2(n_272),
.B1(n_234),
.B2(n_235),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_312),
.B(n_284),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_378),
.B(n_235),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_315),
.Y(n_512)
);

INVx4_ASAP7_75t_L g513 ( 
.A(n_326),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_336),
.A2(n_285),
.B1(n_291),
.B2(n_293),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_386),
.B(n_242),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_385),
.B(n_242),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_379),
.B(n_386),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_317),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_318),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_357),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_379),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_387),
.B(n_259),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_432),
.Y(n_523)
);

NOR2xp67_ASAP7_75t_L g524 ( 
.A(n_439),
.B(n_352),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_438),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_485),
.B(n_336),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_485),
.B(n_336),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_447),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_476),
.B(n_336),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_500),
.B(n_349),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_412),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_480),
.B(n_336),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_483),
.B(n_336),
.Y(n_533)
);

OR2x6_ASAP7_75t_L g534 ( 
.A(n_400),
.B(n_331),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_458),
.A2(n_346),
.B1(n_392),
.B2(n_384),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_481),
.A2(n_399),
.B1(n_395),
.B2(n_387),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_413),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_447),
.B(n_259),
.Y(n_538)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_499),
.B(n_397),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_413),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_492),
.B(n_395),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_491),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_488),
.B(n_399),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g544 ( 
.A(n_440),
.B(n_351),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_400),
.Y(n_545)
);

NOR2x2_ASAP7_75t_L g546 ( 
.A(n_400),
.B(n_320),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_497),
.B(n_344),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_513),
.B(n_268),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_404),
.B(n_268),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_513),
.Y(n_550)
);

NOR2x1_ASAP7_75t_L g551 ( 
.A(n_419),
.B(n_410),
.Y(n_551)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_456),
.B(n_348),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_430),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_410),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_501),
.B(n_272),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_481),
.A2(n_333),
.B1(n_337),
.B2(n_322),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_410),
.B(n_348),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_505),
.B(n_286),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_505),
.B(n_286),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_406),
.B(n_363),
.Y(n_560)
);

NAND2x1p5_ASAP7_75t_L g561 ( 
.A(n_521),
.B(n_363),
.Y(n_561)
);

INVx5_ASAP7_75t_L g562 ( 
.A(n_401),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_496),
.B(n_363),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_507),
.B(n_328),
.Y(n_564)
);

O2A1O1Ixp33_ASAP7_75t_L g565 ( 
.A1(n_490),
.A2(n_495),
.B(n_403),
.C(n_407),
.Y(n_565)
);

OR2x2_ASAP7_75t_L g566 ( 
.A(n_520),
.B(n_495),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_433),
.Y(n_567)
);

INVx5_ASAP7_75t_L g568 ( 
.A(n_401),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_434),
.A2(n_370),
.B(n_343),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_442),
.B(n_460),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_446),
.A2(n_506),
.B1(n_425),
.B2(n_484),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_502),
.B(n_365),
.Y(n_572)
);

A2O1A1Ixp33_ASAP7_75t_L g573 ( 
.A1(n_408),
.A2(n_337),
.B(n_329),
.C(n_343),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_453),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_405),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_453),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_402),
.Y(n_577)
);

OR2x6_ASAP7_75t_L g578 ( 
.A(n_444),
.B(n_365),
.Y(n_578)
);

NOR2x2_ASAP7_75t_L g579 ( 
.A(n_423),
.B(n_329),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_509),
.A2(n_370),
.B1(n_366),
.B2(n_369),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_475),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_508),
.B(n_369),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_468),
.B(n_494),
.Y(n_583)
);

AND2x6_ASAP7_75t_SL g584 ( 
.A(n_464),
.B(n_372),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_424),
.Y(n_585)
);

AND2x2_ASAP7_75t_SL g586 ( 
.A(n_514),
.B(n_370),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_425),
.A2(n_299),
.B1(n_295),
.B2(n_361),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_450),
.B(n_356),
.Y(n_588)
);

OAI22xp33_ASAP7_75t_L g589 ( 
.A1(n_490),
.A2(n_368),
.B1(n_361),
.B2(n_356),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_459),
.B(n_356),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_409),
.B(n_361),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_519),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_414),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_426),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_463),
.A2(n_457),
.B1(n_475),
.B2(n_504),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_512),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_518),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_411),
.B(n_368),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_421),
.B(n_368),
.Y(n_599)
);

NOR2xp67_ASAP7_75t_L g600 ( 
.A(n_487),
.B(n_40),
.Y(n_600)
);

OAI22xp33_ASAP7_75t_L g601 ( 
.A1(n_465),
.A2(n_383),
.B1(n_42),
.B2(n_45),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_467),
.Y(n_602)
);

NOR3xp33_ASAP7_75t_L g603 ( 
.A(n_522),
.B(n_41),
.C(n_47),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_428),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_515),
.B(n_110),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_463),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_466),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_467),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_449),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_482),
.B(n_65),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_515),
.B(n_457),
.Y(n_611)
);

OAI221xp5_ASAP7_75t_L g612 ( 
.A1(n_498),
.A2(n_69),
.B1(n_77),
.B2(n_78),
.C(n_82),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_577),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_523),
.B(n_429),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_545),
.B(n_554),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_528),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_525),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_529),
.A2(n_533),
.B(n_532),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_529),
.A2(n_445),
.B(n_435),
.Y(n_619)
);

OR2x6_ASAP7_75t_L g620 ( 
.A(n_534),
.B(n_429),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_594),
.Y(n_621)
);

NAND2x1p5_ASAP7_75t_L g622 ( 
.A(n_557),
.B(n_537),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_557),
.B(n_593),
.Y(n_623)
);

BUFx2_ASAP7_75t_L g624 ( 
.A(n_584),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_L g625 ( 
.A1(n_569),
.A2(n_517),
.B(n_431),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_578),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_533),
.A2(n_527),
.B(n_526),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_570),
.A2(n_451),
.B1(n_498),
.B2(n_484),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_570),
.B(n_504),
.Y(n_629)
);

INVxp33_ASAP7_75t_L g630 ( 
.A(n_551),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_577),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_571),
.A2(n_504),
.B1(n_473),
.B2(n_443),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_604),
.A2(n_511),
.B1(n_422),
.B2(n_417),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_578),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_581),
.A2(n_417),
.B1(n_422),
.B2(n_416),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_574),
.B(n_418),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_526),
.A2(n_461),
.B(n_449),
.Y(n_637)
);

INVx5_ASAP7_75t_L g638 ( 
.A(n_562),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_566),
.Y(n_639)
);

OR2x6_ASAP7_75t_L g640 ( 
.A(n_534),
.B(n_571),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_550),
.Y(n_641)
);

A2O1A1Ixp33_ASAP7_75t_L g642 ( 
.A1(n_565),
.A2(n_462),
.B(n_473),
.C(n_443),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_583),
.B(n_539),
.Y(n_643)
);

HB1xp67_ASAP7_75t_L g644 ( 
.A(n_578),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_602),
.B(n_462),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_596),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_524),
.B(n_436),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_536),
.B(n_427),
.Y(n_648)
);

OR2x6_ASAP7_75t_L g649 ( 
.A(n_534),
.B(n_420),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_611),
.A2(n_461),
.B(n_449),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_544),
.B(n_415),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_L g652 ( 
.A1(n_573),
.A2(n_493),
.B(n_486),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_562),
.Y(n_653)
);

CKINVDCx8_ASAP7_75t_R g654 ( 
.A(n_542),
.Y(n_654)
);

OR2x6_ASAP7_75t_SL g655 ( 
.A(n_579),
.B(n_441),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_574),
.B(n_427),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_608),
.B(n_441),
.Y(n_657)
);

NAND3xp33_ASAP7_75t_SL g658 ( 
.A(n_606),
.B(n_474),
.C(n_455),
.Y(n_658)
);

BUFx6f_ASAP7_75t_SL g659 ( 
.A(n_540),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_585),
.Y(n_660)
);

O2A1O1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_535),
.A2(n_470),
.B(n_478),
.C(n_503),
.Y(n_661)
);

A2O1A1Ixp33_ASAP7_75t_L g662 ( 
.A1(n_560),
.A2(n_510),
.B(n_478),
.C(n_503),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_576),
.B(n_516),
.Y(n_663)
);

BUFx4f_ASAP7_75t_L g664 ( 
.A(n_561),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_585),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_543),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_561),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_541),
.B(n_479),
.Y(n_668)
);

INVx5_ASAP7_75t_L g669 ( 
.A(n_562),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_607),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_549),
.B(n_479),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_552),
.B(n_477),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_555),
.Y(n_673)
);

BUFx8_ASAP7_75t_L g674 ( 
.A(n_546),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_586),
.A2(n_556),
.B1(n_582),
.B2(n_572),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_543),
.Y(n_676)
);

O2A1O1Ixp33_ASAP7_75t_L g677 ( 
.A1(n_601),
.A2(n_472),
.B(n_471),
.C(n_469),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_567),
.Y(n_678)
);

INVxp33_ASAP7_75t_SL g679 ( 
.A(n_610),
.Y(n_679)
);

NOR3xp33_ASAP7_75t_SL g680 ( 
.A(n_558),
.B(n_83),
.C(n_87),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_547),
.B(n_454),
.Y(n_681)
);

O2A1O1Ixp33_ASAP7_75t_L g682 ( 
.A1(n_589),
.A2(n_452),
.B(n_448),
.C(n_437),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_592),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_591),
.A2(n_94),
.B(n_95),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_575),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_564),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_564),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_559),
.B(n_553),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_580),
.A2(n_118),
.B1(n_119),
.B2(n_122),
.Y(n_689)
);

O2A1O1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_587),
.A2(n_124),
.B(n_128),
.C(n_129),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_609),
.Y(n_691)
);

BUFx8_ASAP7_75t_SL g692 ( 
.A(n_588),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_568),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_597),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_643),
.B(n_563),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_617),
.Y(n_696)
);

A2O1A1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_661),
.A2(n_600),
.B(n_603),
.C(n_605),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_639),
.B(n_538),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_654),
.Y(n_699)
);

O2A1O1Ixp33_ASAP7_75t_L g700 ( 
.A1(n_642),
.A2(n_587),
.B(n_590),
.C(n_612),
.Y(n_700)
);

INVx5_ASAP7_75t_L g701 ( 
.A(n_638),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_620),
.B(n_548),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_653),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_620),
.B(n_531),
.Y(n_704)
);

OA21x2_ASAP7_75t_L g705 ( 
.A1(n_625),
.A2(n_598),
.B(n_599),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_674),
.Y(n_706)
);

OAI22x1_ASAP7_75t_L g707 ( 
.A1(n_626),
.A2(n_142),
.B1(n_144),
.B2(n_146),
.Y(n_707)
);

A2O1A1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_687),
.A2(n_676),
.B(n_666),
.C(n_629),
.Y(n_708)
);

BUFx2_ASAP7_75t_R g709 ( 
.A(n_655),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_694),
.Y(n_710)
);

A2O1A1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_662),
.A2(n_156),
.B(n_157),
.C(n_619),
.Y(n_711)
);

OR2x2_ASAP7_75t_L g712 ( 
.A(n_640),
.B(n_620),
.Y(n_712)
);

O2A1O1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_633),
.A2(n_640),
.B(n_658),
.C(n_614),
.Y(n_713)
);

AOI221xp5_ASAP7_75t_L g714 ( 
.A1(n_645),
.A2(n_651),
.B1(n_644),
.B2(n_634),
.C(n_624),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_640),
.A2(n_649),
.B1(n_623),
.B2(n_679),
.Y(n_715)
);

BUFx4f_ASAP7_75t_SL g716 ( 
.A(n_674),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_657),
.B(n_646),
.Y(n_717)
);

A2O1A1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_677),
.A2(n_689),
.B(n_682),
.C(n_656),
.Y(n_718)
);

O2A1O1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_635),
.A2(n_670),
.B(n_663),
.C(n_681),
.Y(n_719)
);

INVx8_ASAP7_75t_L g720 ( 
.A(n_659),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_630),
.B(n_623),
.Y(n_721)
);

OAI22x1_ASAP7_75t_L g722 ( 
.A1(n_689),
.A2(n_647),
.B1(n_622),
.B2(n_667),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_616),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_649),
.A2(n_615),
.B1(n_647),
.B2(n_659),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_649),
.B(n_646),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_616),
.Y(n_726)
);

INVx4_ASAP7_75t_L g727 ( 
.A(n_638),
.Y(n_727)
);

A2O1A1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_690),
.A2(n_683),
.B(n_680),
.C(n_685),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_615),
.A2(n_688),
.B1(n_692),
.B2(n_664),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_671),
.A2(n_668),
.B(n_636),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_638),
.Y(n_731)
);

AOI211x1_ASAP7_75t_L g732 ( 
.A1(n_672),
.A2(n_613),
.B(n_631),
.C(n_684),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_669),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_660),
.A2(n_665),
.B(n_621),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_669),
.B(n_693),
.Y(n_735)
);

NAND2x1p5_ASAP7_75t_L g736 ( 
.A(n_641),
.B(n_664),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_639),
.A2(n_489),
.B1(n_523),
.B2(n_571),
.Y(n_737)
);

A2O1A1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_661),
.A2(n_632),
.B(n_481),
.C(n_458),
.Y(n_738)
);

OAI21xp33_ASAP7_75t_L g739 ( 
.A1(n_614),
.A2(n_523),
.B(n_432),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_691),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_640),
.B(n_649),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_643),
.B(n_523),
.Y(n_742)
);

OAI22xp33_ASAP7_75t_L g743 ( 
.A1(n_640),
.A2(n_489),
.B1(n_396),
.B2(n_523),
.Y(n_743)
);

BUFx8_ASAP7_75t_L g744 ( 
.A(n_659),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_SL g745 ( 
.A(n_617),
.B(n_523),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_617),
.B(n_523),
.Y(n_746)
);

AO31x2_ASAP7_75t_L g747 ( 
.A1(n_675),
.A2(n_573),
.A3(n_569),
.B(n_650),
.Y(n_747)
);

A2O1A1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_661),
.A2(n_632),
.B(n_481),
.C(n_458),
.Y(n_748)
);

OAI21xp5_ASAP7_75t_L g749 ( 
.A1(n_627),
.A2(n_618),
.B(n_637),
.Y(n_749)
);

OAI21xp5_ASAP7_75t_L g750 ( 
.A1(n_627),
.A2(n_618),
.B(n_637),
.Y(n_750)
);

OAI21xp5_ASAP7_75t_L g751 ( 
.A1(n_627),
.A2(n_618),
.B(n_637),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_678),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_SL g753 ( 
.A(n_617),
.B(n_523),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_691),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_678),
.Y(n_755)
);

OAI221xp5_ASAP7_75t_L g756 ( 
.A1(n_673),
.A2(n_571),
.B1(n_523),
.B2(n_535),
.C(n_639),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_686),
.Y(n_757)
);

AOI21xp33_ASAP7_75t_L g758 ( 
.A1(n_614),
.A2(n_432),
.B(n_523),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_643),
.B(n_530),
.Y(n_759)
);

A2O1A1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_661),
.A2(n_632),
.B(n_481),
.C(n_458),
.Y(n_760)
);

O2A1O1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_642),
.A2(n_648),
.B(n_571),
.C(n_628),
.Y(n_761)
);

OA21x2_ASAP7_75t_L g762 ( 
.A1(n_652),
.A2(n_569),
.B(n_573),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_678),
.Y(n_763)
);

INVxp67_ASAP7_75t_SL g764 ( 
.A(n_639),
.Y(n_764)
);

AO31x2_ASAP7_75t_L g765 ( 
.A1(n_675),
.A2(n_573),
.A3(n_569),
.B(n_650),
.Y(n_765)
);

A2O1A1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_661),
.A2(n_632),
.B(n_481),
.C(n_458),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_654),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_640),
.B(n_649),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_643),
.B(n_530),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_640),
.A2(n_458),
.B1(n_481),
.B2(n_571),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_654),
.Y(n_771)
);

OAI21x1_ASAP7_75t_SL g772 ( 
.A1(n_666),
.A2(n_595),
.B(n_676),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_678),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_L g774 ( 
.A1(n_686),
.A2(n_481),
.B1(n_458),
.B2(n_687),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_654),
.Y(n_775)
);

NAND2x1p5_ASAP7_75t_L g776 ( 
.A(n_664),
.B(n_617),
.Y(n_776)
);

A2O1A1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_661),
.A2(n_632),
.B(n_481),
.C(n_458),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_643),
.B(n_523),
.Y(n_778)
);

AO31x2_ASAP7_75t_L g779 ( 
.A1(n_675),
.A2(n_573),
.A3(n_569),
.B(n_650),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_686),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_678),
.Y(n_781)
);

NAND2x1_ASAP7_75t_L g782 ( 
.A(n_653),
.B(n_686),
.Y(n_782)
);

A2O1A1Ixp33_ASAP7_75t_L g783 ( 
.A1(n_661),
.A2(n_632),
.B(n_481),
.C(n_458),
.Y(n_783)
);

NAND2x1_ASAP7_75t_L g784 ( 
.A(n_653),
.B(n_686),
.Y(n_784)
);

A2O1A1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_661),
.A2(n_632),
.B(n_481),
.C(n_458),
.Y(n_785)
);

AO31x2_ASAP7_75t_L g786 ( 
.A1(n_675),
.A2(n_573),
.A3(n_569),
.B(n_650),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_617),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_643),
.B(n_530),
.Y(n_788)
);

AO31x2_ASAP7_75t_L g789 ( 
.A1(n_718),
.A2(n_711),
.A3(n_738),
.B(n_760),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_743),
.B(n_739),
.Y(n_790)
);

OAI221xp5_ASAP7_75t_L g791 ( 
.A1(n_756),
.A2(n_737),
.B1(n_770),
.B2(n_714),
.C(n_715),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_SL g792 ( 
.A1(n_745),
.A2(n_753),
.B1(n_768),
.B2(n_741),
.Y(n_792)
);

OAI221xp5_ASAP7_75t_L g793 ( 
.A1(n_713),
.A2(n_695),
.B1(n_758),
.B2(n_788),
.C(n_759),
.Y(n_793)
);

OR2x6_ASAP7_75t_L g794 ( 
.A(n_720),
.B(n_741),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_768),
.A2(n_778),
.B1(n_742),
.B2(n_746),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_769),
.B(n_764),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_748),
.A2(n_783),
.B1(n_785),
.B2(n_777),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_696),
.B(n_712),
.Y(n_798)
);

INVx4_ASAP7_75t_L g799 ( 
.A(n_701),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_710),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_757),
.B(n_780),
.Y(n_801)
);

AO31x2_ASAP7_75t_L g802 ( 
.A1(n_766),
.A2(n_697),
.A3(n_708),
.B(n_722),
.Y(n_802)
);

A2O1A1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_700),
.A2(n_719),
.B(n_730),
.C(n_728),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_787),
.A2(n_774),
.B1(n_698),
.B2(n_702),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_776),
.B(n_729),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_721),
.B(n_724),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_752),
.B(n_755),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_SL g808 ( 
.A1(n_744),
.A2(n_720),
.B1(n_716),
.B2(n_701),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_701),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_744),
.Y(n_810)
);

AOI211xp5_ASAP7_75t_L g811 ( 
.A1(n_704),
.A2(n_725),
.B(n_717),
.C(n_773),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_763),
.B(n_781),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_732),
.B(n_734),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_703),
.A2(n_727),
.B1(n_733),
.B2(n_731),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_762),
.B(n_703),
.Y(n_815)
);

INVx6_ASAP7_75t_L g816 ( 
.A(n_727),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_735),
.B(n_731),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_699),
.Y(n_818)
);

INVx4_ASAP7_75t_L g819 ( 
.A(n_771),
.Y(n_819)
);

OAI22xp33_ASAP7_75t_L g820 ( 
.A1(n_706),
.A2(n_775),
.B1(n_767),
.B2(n_736),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_705),
.A2(n_784),
.B(n_782),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_709),
.B(n_723),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_707),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_723),
.A2(n_726),
.B1(n_740),
.B2(n_754),
.Y(n_824)
);

AO31x2_ASAP7_75t_L g825 ( 
.A1(n_747),
.A2(n_786),
.A3(n_779),
.B(n_765),
.Y(n_825)
);

OAI21x1_ASAP7_75t_L g826 ( 
.A1(n_747),
.A2(n_765),
.B(n_779),
.Y(n_826)
);

AO21x2_ASAP7_75t_L g827 ( 
.A1(n_749),
.A2(n_751),
.B(n_750),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_743),
.B(n_620),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_787),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_743),
.B(n_620),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_742),
.B(n_778),
.Y(n_831)
);

OR2x6_ASAP7_75t_L g832 ( 
.A(n_720),
.B(n_489),
.Y(n_832)
);

BUFx12f_ASAP7_75t_L g833 ( 
.A(n_744),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_743),
.A2(n_640),
.B1(n_534),
.B2(n_481),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_761),
.B(n_666),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_761),
.B(n_666),
.Y(n_836)
);

AO31x2_ASAP7_75t_L g837 ( 
.A1(n_718),
.A2(n_573),
.A3(n_711),
.B(n_738),
.Y(n_837)
);

BUFx8_ASAP7_75t_L g838 ( 
.A(n_699),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_743),
.A2(n_640),
.B1(n_534),
.B2(n_481),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_744),
.Y(n_840)
);

OAI21x1_ASAP7_75t_SL g841 ( 
.A1(n_770),
.A2(n_772),
.B(n_713),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_743),
.A2(n_640),
.B1(n_534),
.B2(n_481),
.Y(n_842)
);

O2A1O1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_756),
.A2(n_743),
.B(n_642),
.C(n_571),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_815),
.Y(n_844)
);

OR2x6_ASAP7_75t_L g845 ( 
.A(n_841),
.B(n_821),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_825),
.B(n_826),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_825),
.B(n_827),
.Y(n_847)
);

INVxp67_ASAP7_75t_L g848 ( 
.A(n_829),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_815),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_813),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_790),
.A2(n_828),
.B1(n_830),
.B2(n_791),
.Y(n_851)
);

OR2x6_ASAP7_75t_L g852 ( 
.A(n_821),
.B(n_797),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_843),
.A2(n_803),
.B(n_793),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_SL g854 ( 
.A1(n_824),
.A2(n_799),
.B(n_823),
.Y(n_854)
);

OAI222xp33_ASAP7_75t_L g855 ( 
.A1(n_791),
.A2(n_842),
.B1(n_839),
.B2(n_834),
.C1(n_792),
.C2(n_832),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_793),
.A2(n_835),
.B(n_836),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_802),
.Y(n_857)
);

AOI222xp33_ASAP7_75t_L g858 ( 
.A1(n_831),
.A2(n_795),
.B1(n_806),
.B2(n_807),
.C1(n_812),
.C2(n_796),
.Y(n_858)
);

INVxp67_ASAP7_75t_L g859 ( 
.A(n_801),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_802),
.Y(n_860)
);

OAI221xp5_ASAP7_75t_L g861 ( 
.A1(n_804),
.A2(n_811),
.B1(n_832),
.B2(n_808),
.C(n_807),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_809),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_800),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_847),
.B(n_789),
.Y(n_864)
);

BUFx2_ASAP7_75t_L g865 ( 
.A(n_844),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_847),
.B(n_837),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_847),
.B(n_837),
.Y(n_867)
);

OR2x2_ASAP7_75t_L g868 ( 
.A(n_844),
.B(n_805),
.Y(n_868)
);

OAI21xp33_ASAP7_75t_L g869 ( 
.A1(n_861),
.A2(n_832),
.B(n_798),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_850),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_861),
.A2(n_851),
.B1(n_858),
.B2(n_853),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_845),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_849),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_846),
.B(n_817),
.Y(n_874)
);

AOI211xp5_ASAP7_75t_L g875 ( 
.A1(n_855),
.A2(n_820),
.B(n_822),
.C(n_810),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_852),
.B(n_794),
.Y(n_876)
);

INVxp67_ASAP7_75t_SL g877 ( 
.A(n_859),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_859),
.A2(n_794),
.B1(n_816),
.B2(n_814),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_864),
.B(n_866),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_870),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_872),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_872),
.B(n_852),
.Y(n_882)
);

AND2x4_ASAP7_75t_SL g883 ( 
.A(n_876),
.B(n_845),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_864),
.B(n_857),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_864),
.B(n_857),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_866),
.B(n_857),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_873),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_866),
.B(n_860),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_867),
.B(n_860),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_865),
.Y(n_890)
);

NAND2x1_ASAP7_75t_L g891 ( 
.A(n_881),
.B(n_876),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_880),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_879),
.B(n_867),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_879),
.B(n_868),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_879),
.B(n_877),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_880),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_884),
.B(n_867),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_884),
.B(n_874),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_884),
.B(n_874),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_885),
.B(n_886),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_885),
.B(n_886),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_885),
.B(n_818),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_890),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_886),
.B(n_874),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_901),
.B(n_888),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_902),
.A2(n_869),
.B1(n_871),
.B2(n_875),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_892),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_901),
.B(n_888),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_903),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_893),
.B(n_888),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_892),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_900),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_896),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_896),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_898),
.B(n_889),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_891),
.B(n_883),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_894),
.Y(n_917)
);

OR2x2_ASAP7_75t_L g918 ( 
.A(n_900),
.B(n_890),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_893),
.B(n_898),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_912),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_907),
.Y(n_921)
);

NAND3xp33_ASAP7_75t_L g922 ( 
.A(n_906),
.B(n_875),
.C(n_869),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_919),
.B(n_899),
.Y(n_923)
);

AOI332xp33_ASAP7_75t_L g924 ( 
.A1(n_917),
.A2(n_851),
.A3(n_904),
.B1(n_899),
.B2(n_895),
.B3(n_897),
.C1(n_863),
.C2(n_889),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_919),
.B(n_904),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_912),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_911),
.Y(n_927)
);

OAI21xp33_ASAP7_75t_L g928 ( 
.A1(n_918),
.A2(n_894),
.B(n_897),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_913),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_914),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_918),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_910),
.B(n_889),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_910),
.B(n_887),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_921),
.Y(n_934)
);

AOI221xp5_ASAP7_75t_SL g935 ( 
.A1(n_928),
.A2(n_915),
.B1(n_905),
.B2(n_908),
.C(n_855),
.Y(n_935)
);

O2A1O1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_922),
.A2(n_909),
.B(n_878),
.C(n_848),
.Y(n_936)
);

OAI31xp33_ASAP7_75t_L g937 ( 
.A1(n_920),
.A2(n_916),
.A3(n_909),
.B(n_876),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_921),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_926),
.A2(n_876),
.B1(n_882),
.B2(n_916),
.Y(n_939)
);

NAND2x1_ASAP7_75t_L g940 ( 
.A(n_923),
.B(n_916),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_SL g941 ( 
.A1(n_937),
.A2(n_936),
.B(n_939),
.Y(n_941)
);

AOI221xp5_ASAP7_75t_L g942 ( 
.A1(n_935),
.A2(n_940),
.B1(n_938),
.B2(n_934),
.C(n_931),
.Y(n_942)
);

NOR2x1_ASAP7_75t_L g943 ( 
.A(n_940),
.B(n_840),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_934),
.B(n_923),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_940),
.Y(n_945)
);

AOI221xp5_ASAP7_75t_L g946 ( 
.A1(n_935),
.A2(n_929),
.B1(n_930),
.B2(n_927),
.C(n_933),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_944),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_946),
.B(n_925),
.Y(n_948)
);

AND4x1_ASAP7_75t_L g949 ( 
.A(n_943),
.B(n_833),
.C(n_838),
.D(n_858),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_945),
.Y(n_950)
);

NAND5xp2_ASAP7_75t_L g951 ( 
.A(n_948),
.B(n_941),
.C(n_942),
.D(n_924),
.E(n_853),
.Y(n_951)
);

NAND4xp25_ASAP7_75t_SL g952 ( 
.A(n_947),
.B(n_932),
.C(n_925),
.D(n_854),
.Y(n_952)
);

AOI211xp5_ASAP7_75t_L g953 ( 
.A1(n_950),
.A2(n_947),
.B(n_949),
.C(n_876),
.Y(n_953)
);

NAND4xp75_ASAP7_75t_L g954 ( 
.A(n_948),
.B(n_838),
.C(n_856),
.D(n_927),
.Y(n_954)
);

XOR2xp5_ASAP7_75t_L g955 ( 
.A(n_954),
.B(n_862),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_952),
.Y(n_956)
);

XNOR2xp5_ASAP7_75t_L g957 ( 
.A(n_955),
.B(n_956),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_955),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_958),
.B(n_953),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_959),
.Y(n_960)
);

NAND3xp33_ASAP7_75t_L g961 ( 
.A(n_960),
.B(n_957),
.C(n_819),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_961),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_962),
.A2(n_951),
.B1(n_819),
.B2(n_848),
.Y(n_963)
);


endmodule