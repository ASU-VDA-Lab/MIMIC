module fake_jpeg_25766_n_194 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_194);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_194;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_9),
.B(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_1),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_17),
.B(n_19),
.C(n_34),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_47),
.Y(n_59)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_23),
.Y(n_57)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx5_ASAP7_75t_SL g65 ( 
.A(n_44),
.Y(n_65)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_26),
.B(n_33),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_27),
.Y(n_58)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_22),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_50),
.B(n_29),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_27),
.C(n_19),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_30),
.Y(n_78)
);

NOR3xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_33),
.C(n_23),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_52),
.A2(n_74),
.B(n_16),
.Y(n_93)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_46),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_58),
.B(n_68),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_60),
.A2(n_61),
.B(n_17),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_31),
.B(n_29),
.C(n_28),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_73),
.Y(n_83)
);

BUFx16f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_20),
.B1(n_26),
.B2(n_21),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_42),
.B1(n_45),
.B2(n_40),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_31),
.Y(n_68)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

NAND2x1_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_26),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_28),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_15),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_32),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_78),
.B(n_92),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_85),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_55),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_75),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_58),
.A2(n_35),
.B1(n_20),
.B2(n_34),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_86),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_38),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_90),
.Y(n_105)
);

AND2x6_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_14),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_37),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_95),
.Y(n_106)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_32),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_98),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_53),
.A2(n_20),
.B1(n_16),
.B2(n_25),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_65),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

OAI22x1_ASAP7_75t_SL g100 ( 
.A1(n_67),
.A2(n_21),
.B1(n_2),
.B2(n_3),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_56),
.B(n_55),
.C(n_71),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_72),
.A2(n_30),
.B1(n_25),
.B2(n_21),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_72),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_70),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_103),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_99),
.B1(n_88),
.B2(n_101),
.Y(n_127)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_113),
.Y(n_129)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_66),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_115),
.B(n_119),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_83),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_116),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_117),
.A2(n_121),
.B(n_75),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_66),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_80),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_98),
.B(n_86),
.Y(n_136)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_135),
.B1(n_110),
.B2(n_121),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_91),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_1),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_104),
.B(n_91),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_131),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_79),
.Y(n_131)
);

AND2x4_ASAP7_75t_SL g133 ( 
.A(n_115),
.B(n_100),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_133),
.A2(n_138),
.B(n_140),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_92),
.B1(n_82),
.B2(n_94),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_136),
.B(n_139),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_78),
.C(n_84),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_107),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_111),
.A2(n_93),
.B1(n_90),
.B2(n_89),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_87),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_89),
.B(n_2),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_142),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_133),
.A2(n_108),
.B1(n_105),
.B2(n_135),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_149),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_133),
.A2(n_105),
.B1(n_108),
.B2(n_121),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_145),
.A2(n_146),
.B(n_142),
.Y(n_164)
);

AOI221xp5_ASAP7_75t_L g146 ( 
.A1(n_137),
.A2(n_110),
.B1(n_104),
.B2(n_107),
.C(n_112),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_147),
.B(n_155),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_106),
.C(n_112),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_150),
.C(n_138),
.Y(n_160)
);

MAJx2_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_116),
.C(n_123),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_152),
.B(n_153),
.Y(n_158)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

INVxp67_ASAP7_75t_SL g167 ( 
.A(n_154),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_161),
.C(n_125),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_141),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_143),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_162),
.B(n_157),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_150),
.B(n_140),
.Y(n_163)
);

AOI321xp33_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_164),
.A3(n_11),
.B1(n_15),
.B2(n_10),
.C(n_6),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_151),
.A2(n_134),
.B(n_132),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_166),
.A2(n_145),
.B1(n_144),
.B2(n_127),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_134),
.C(n_132),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_156),
.C(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_169),
.B(n_173),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_172),
.Y(n_180)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_155),
.C(n_125),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_175),
.Y(n_181)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_167),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_114),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_182),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_170),
.B(n_168),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_177),
.A2(n_165),
.B(n_163),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_184),
.A2(n_186),
.B(n_3),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_179),
.A2(n_113),
.B1(n_160),
.B2(n_81),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_SL g189 ( 
.A1(n_185),
.A2(n_187),
.B(n_64),
.C(n_118),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_159),
.C(n_173),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_180),
.A2(n_181),
.B1(n_159),
.B2(n_81),
.Y(n_187)
);

AOI322xp5_ASAP7_75t_L g188 ( 
.A1(n_183),
.A2(n_180),
.A3(n_118),
.B1(n_5),
.B2(n_6),
.C1(n_3),
.C2(n_4),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_188),
.A2(n_189),
.B1(n_186),
.B2(n_5),
.Y(n_192)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_190),
.Y(n_191)
);

OAI321xp33_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_4),
.A3(n_5),
.B1(n_8),
.B2(n_118),
.C(n_191),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_8),
.Y(n_194)
);


endmodule