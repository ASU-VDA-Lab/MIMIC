module fake_ariane_2533_n_1702 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1702);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1702;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_73),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_150),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_23),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_72),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_105),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_103),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_155),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_95),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_126),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_67),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_84),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_108),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_146),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_129),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_33),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_65),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_35),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_68),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_66),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_115),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_81),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_97),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_100),
.Y(n_182)
);

BUFx10_ASAP7_75t_L g183 ( 
.A(n_137),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_83),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_122),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_152),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_133),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_8),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_130),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_33),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_41),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_111),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_53),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_96),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_82),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_46),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_12),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_19),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_86),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_18),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_144),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_99),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_52),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_12),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_87),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_91),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_26),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_139),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_15),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_147),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g212 ( 
.A(n_61),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_70),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_124),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_10),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_75),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_3),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_116),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_123),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_142),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_101),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_119),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_19),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_132),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_114),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_26),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_106),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_4),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_120),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_8),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_113),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_127),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_31),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_31),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_34),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_74),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_6),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_107),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_71),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_16),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_13),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_24),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_56),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_136),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_145),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_37),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_125),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_77),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_34),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_141),
.Y(n_250)
);

BUFx10_ASAP7_75t_L g251 ( 
.A(n_14),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_10),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_92),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_20),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_157),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_15),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_53),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_60),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_156),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_57),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_36),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_69),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_1),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_93),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_44),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_0),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_55),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_79),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_9),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_118),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_52),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_58),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_21),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_21),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_85),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_151),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_143),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_89),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_90),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_138),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_28),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_5),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_37),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_45),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_20),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_80),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_121),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_35),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_41),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_88),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_27),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_76),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_24),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_59),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_102),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_63),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_49),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_62),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_1),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_3),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_64),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_16),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_14),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_42),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_38),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_9),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_11),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_32),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_154),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_2),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_11),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_55),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_117),
.Y(n_313)
);

BUFx2_ASAP7_75t_SL g314 ( 
.A(n_7),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_28),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_4),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_44),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_27),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_289),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_230),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_166),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_230),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_230),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_230),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_230),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_190),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_306),
.Y(n_327)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_160),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_306),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_225),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_225),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_262),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_262),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_173),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_280),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_280),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_189),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_193),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_209),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_191),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_197),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_227),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_204),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_238),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_176),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_245),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_188),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_234),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_205),
.Y(n_349)
);

INVxp33_ASAP7_75t_L g350 ( 
.A(n_215),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_173),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_217),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_223),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_192),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_226),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_237),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_261),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_314),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_274),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_188),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_194),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_257),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_281),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_282),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_176),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_293),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_303),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_312),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_167),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_168),
.Y(n_370)
);

CKINVDCx14_ASAP7_75t_R g371 ( 
.A(n_183),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_174),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_249),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_249),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_175),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_198),
.Y(n_376)
);

INVxp33_ASAP7_75t_SL g377 ( 
.A(n_297),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_178),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_218),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_172),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_216),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_224),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_229),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_244),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_214),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_259),
.Y(n_386)
);

INVxp33_ASAP7_75t_SL g387 ( 
.A(n_297),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_260),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_264),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_251),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_288),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_270),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_278),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_279),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_236),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_251),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_320),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_319),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_320),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_321),
.Y(n_400)
);

NAND2xp33_ASAP7_75t_SL g401 ( 
.A(n_328),
.B(n_300),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_380),
.B(n_219),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_325),
.Y(n_403)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_347),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_322),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_348),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_322),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_325),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_323),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_347),
.B(n_255),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_323),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_324),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_326),
.Y(n_413)
);

OAI21x1_ASAP7_75t_L g414 ( 
.A1(n_330),
.A2(n_298),
.B(n_295),
.Y(n_414)
);

NOR2x1_ASAP7_75t_L g415 ( 
.A(n_330),
.B(n_216),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_360),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_369),
.B(n_250),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_338),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_360),
.B(n_301),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_324),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_331),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_331),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_332),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_332),
.Y(n_424)
);

OAI21x1_ASAP7_75t_L g425 ( 
.A1(n_333),
.A2(n_212),
.B(n_186),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_333),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_369),
.B(n_370),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_335),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_370),
.B(n_183),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_335),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_336),
.Y(n_431)
);

OA21x2_ASAP7_75t_L g432 ( 
.A1(n_336),
.A2(n_231),
.B(n_171),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_327),
.Y(n_433)
);

NOR2xp67_ASAP7_75t_L g434 ( 
.A(n_372),
.B(n_171),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_372),
.Y(n_435)
);

CKINVDCx14_ASAP7_75t_R g436 ( 
.A(n_371),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_375),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_327),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_339),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_375),
.B(n_250),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_378),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_381),
.B(n_378),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_381),
.B(n_158),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_329),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_R g445 ( 
.A(n_354),
.B(n_187),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_379),
.B(n_382),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_385),
.B(n_183),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_379),
.B(n_158),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_344),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_329),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_382),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_383),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_357),
.Y(n_453)
);

AND2x6_ASAP7_75t_L g454 ( 
.A(n_383),
.B(n_211),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_384),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_365),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_384),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_386),
.B(n_251),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_386),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_388),
.B(n_159),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_388),
.B(n_159),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_389),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_359),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_389),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_346),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_392),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_392),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_393),
.B(n_256),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_361),
.B(n_376),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_393),
.B(n_231),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_409),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_404),
.B(n_377),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_400),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_409),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_R g475 ( 
.A(n_413),
.B(n_342),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_450),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_408),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_429),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_409),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_404),
.B(n_387),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_L g481 ( 
.A1(n_470),
.A2(n_395),
.B1(n_365),
.B2(n_350),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_445),
.B(n_390),
.Y(n_482)
);

NAND2xp33_ASAP7_75t_L g483 ( 
.A(n_448),
.B(n_161),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_429),
.B(n_394),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_408),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_408),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_429),
.B(n_334),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_398),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_397),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_412),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_412),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_458),
.B(n_351),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_412),
.Y(n_493)
);

AND2x6_ASAP7_75t_L g494 ( 
.A(n_458),
.B(n_211),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_404),
.B(n_394),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_450),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_458),
.B(n_396),
.Y(n_497)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_457),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_423),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_408),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_423),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_404),
.B(n_358),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_423),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_408),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_397),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_469),
.B(n_345),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_423),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_423),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_399),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_423),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_399),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_468),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_405),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_405),
.Y(n_514)
);

INVx8_ASAP7_75t_L g515 ( 
.A(n_454),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_407),
.Y(n_516)
);

NAND2xp33_ASAP7_75t_SL g517 ( 
.A(n_398),
.B(n_300),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_468),
.B(n_161),
.Y(n_518)
);

CKINVDCx11_ASAP7_75t_R g519 ( 
.A(n_406),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_470),
.A2(n_373),
.B1(n_374),
.B2(n_302),
.Y(n_520)
);

NAND3xp33_ASAP7_75t_L g521 ( 
.A(n_457),
.B(n_363),
.C(n_362),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_468),
.B(n_162),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_407),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_411),
.Y(n_524)
);

BUFx10_ASAP7_75t_L g525 ( 
.A(n_410),
.Y(n_525)
);

OR2x6_ASAP7_75t_L g526 ( 
.A(n_470),
.B(n_442),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_411),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_420),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_420),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_403),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_408),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_446),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_456),
.B(n_364),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_450),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_418),
.B(n_299),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_446),
.B(n_337),
.Y(n_536)
);

NAND3xp33_ASAP7_75t_L g537 ( 
.A(n_457),
.B(n_163),
.C(n_162),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_446),
.B(n_163),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_446),
.B(n_337),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_427),
.B(n_340),
.Y(n_540)
);

OAI22xp33_ASAP7_75t_L g541 ( 
.A1(n_456),
.A2(n_316),
.B1(n_305),
.B2(n_307),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_447),
.B(n_340),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_457),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_422),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_457),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_422),
.Y(n_546)
);

INVx5_ASAP7_75t_L g547 ( 
.A(n_454),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_470),
.A2(n_256),
.B1(n_265),
.B2(n_367),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_457),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_453),
.B(n_391),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_431),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_431),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_417),
.A2(n_256),
.B1(n_265),
.B2(n_366),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_431),
.Y(n_554)
);

OAI21xp33_ASAP7_75t_SL g555 ( 
.A1(n_427),
.A2(n_343),
.B(n_341),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_SL g556 ( 
.A1(n_439),
.A2(n_265),
.B1(n_304),
.B2(n_317),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_448),
.B(n_341),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_401),
.B(n_164),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_462),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_427),
.B(n_343),
.Y(n_560)
);

OR2x6_ASAP7_75t_L g561 ( 
.A(n_442),
.B(n_349),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_449),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_450),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_462),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_450),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_462),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_417),
.B(n_349),
.Y(n_567)
);

INVx5_ASAP7_75t_L g568 ( 
.A(n_454),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_450),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_403),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_403),
.Y(n_571)
);

INVxp67_ASAP7_75t_SL g572 ( 
.A(n_416),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_430),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_417),
.A2(n_368),
.B1(n_367),
.B2(n_366),
.Y(n_574)
);

BUFx6f_ASAP7_75t_SL g575 ( 
.A(n_417),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_440),
.B(n_352),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_403),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_430),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_433),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_433),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_460),
.B(n_164),
.Y(n_581)
);

AO21x2_ASAP7_75t_L g582 ( 
.A1(n_414),
.A2(n_368),
.B(n_356),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_432),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_433),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_440),
.B(n_352),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_438),
.Y(n_586)
);

AO21x2_ASAP7_75t_L g587 ( 
.A1(n_414),
.A2(n_356),
.B(n_355),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_416),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_435),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_416),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_465),
.Y(n_591)
);

OR2x6_ASAP7_75t_L g592 ( 
.A(n_440),
.B(n_353),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_460),
.B(n_353),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_440),
.B(n_355),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_438),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_435),
.B(n_304),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_437),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_437),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_438),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_441),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_461),
.B(n_443),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_432),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_461),
.B(n_165),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_444),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_441),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_451),
.B(n_305),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_432),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_451),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_452),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_444),
.Y(n_610)
);

AND3x2_ASAP7_75t_L g611 ( 
.A(n_410),
.B(n_307),
.C(n_317),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_454),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_444),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_443),
.B(n_195),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_434),
.B(n_308),
.Y(n_615)
);

OAI22xp33_ASAP7_75t_L g616 ( 
.A1(n_402),
.A2(n_308),
.B1(n_315),
.B2(n_310),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_452),
.B(n_165),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_414),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_532),
.B(n_455),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_528),
.Y(n_620)
);

NAND2xp33_ASAP7_75t_SL g621 ( 
.A(n_562),
.B(n_455),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_528),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_600),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_600),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_600),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_601),
.B(n_459),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_489),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_492),
.B(n_436),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_505),
.Y(n_629)
);

AND2x6_ASAP7_75t_L g630 ( 
.A(n_618),
.B(n_464),
.Y(n_630)
);

INVxp67_ASAP7_75t_SL g631 ( 
.A(n_532),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_528),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_505),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_478),
.B(n_512),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_557),
.B(n_593),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_492),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_509),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_492),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_478),
.B(n_512),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_492),
.B(n_464),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_487),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_614),
.B(n_466),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_525),
.B(n_466),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_509),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_511),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_550),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_484),
.B(n_467),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_550),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_487),
.B(n_467),
.Y(n_649)
);

INVxp67_ASAP7_75t_SL g650 ( 
.A(n_590),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_539),
.B(n_434),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_488),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_511),
.Y(n_653)
);

OAI22xp33_ASAP7_75t_L g654 ( 
.A1(n_561),
.A2(n_424),
.B1(n_421),
.B2(n_428),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_535),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_561),
.A2(n_432),
.B1(n_421),
.B2(n_426),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_539),
.B(n_419),
.Y(n_657)
);

NAND2xp33_ASAP7_75t_L g658 ( 
.A(n_573),
.B(n_454),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_525),
.B(n_169),
.Y(n_659)
);

OAI22xp33_ASAP7_75t_L g660 ( 
.A1(n_561),
.A2(n_428),
.B1(n_426),
.B2(n_424),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_533),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_588),
.Y(n_662)
);

INVx4_ASAP7_75t_L g663 ( 
.A(n_515),
.Y(n_663)
);

OR2x6_ASAP7_75t_L g664 ( 
.A(n_592),
.B(n_419),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_588),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_591),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_539),
.B(n_415),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_588),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_513),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_513),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_526),
.A2(n_561),
.B1(n_592),
.B2(n_539),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_514),
.Y(n_672)
);

AND2x6_ASAP7_75t_SL g673 ( 
.A(n_506),
.B(n_463),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_494),
.A2(n_415),
.B1(n_287),
.B2(n_290),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_494),
.B(n_432),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_590),
.Y(n_676)
);

INVxp67_ASAP7_75t_L g677 ( 
.A(n_473),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_516),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_516),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_544),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_592),
.B(n_310),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_525),
.B(n_169),
.Y(n_682)
);

INVxp67_ASAP7_75t_L g683 ( 
.A(n_542),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_525),
.B(n_170),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_494),
.B(n_207),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_523),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_494),
.B(n_248),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_494),
.B(n_268),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_555),
.B(n_170),
.Y(n_689)
);

AOI221xp5_ASAP7_75t_L g690 ( 
.A1(n_541),
.A2(n_311),
.B1(n_315),
.B2(n_318),
.C(n_235),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_494),
.B(n_275),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_523),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_524),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_561),
.A2(n_454),
.B1(n_287),
.B2(n_290),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_555),
.B(n_177),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_494),
.B(n_177),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_578),
.B(n_179),
.Y(n_697)
);

NOR3xp33_ASAP7_75t_L g698 ( 
.A(n_591),
.B(n_556),
.C(n_517),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_540),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_472),
.B(n_179),
.Y(n_700)
);

OR2x2_ASAP7_75t_L g701 ( 
.A(n_481),
.B(n_311),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_578),
.B(n_180),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_527),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_480),
.B(n_180),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_527),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_540),
.B(n_181),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_544),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_560),
.B(n_181),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_560),
.B(n_182),
.Y(n_709)
);

A2O1A1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_589),
.A2(n_425),
.B(n_199),
.C(n_228),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_578),
.B(n_536),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_578),
.B(n_182),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_589),
.B(n_597),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_529),
.Y(n_714)
);

AND2x6_ASAP7_75t_SL g715 ( 
.A(n_519),
.B(n_201),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_597),
.B(n_184),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_592),
.B(n_425),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_598),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_598),
.B(n_605),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_SL g720 ( 
.A1(n_548),
.A2(n_283),
.B1(n_254),
.B2(n_252),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_605),
.A2(n_454),
.B1(n_425),
.B2(n_291),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_608),
.B(n_184),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_608),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_596),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_590),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_609),
.A2(n_454),
.B1(n_240),
.B2(n_208),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_609),
.B(n_185),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_502),
.B(n_567),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_526),
.A2(n_454),
.B1(n_246),
.B2(n_241),
.Y(n_729)
);

NAND3xp33_ASAP7_75t_L g730 ( 
.A(n_497),
.B(n_210),
.C(n_233),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_546),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_596),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_546),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_576),
.B(n_185),
.Y(n_734)
);

BUFx2_ASAP7_75t_L g735 ( 
.A(n_475),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_606),
.B(n_242),
.Y(n_736)
);

OR2x6_ASAP7_75t_L g737 ( 
.A(n_592),
.B(n_211),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_554),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_606),
.B(n_263),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_573),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_590),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_583),
.B(n_309),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_585),
.B(n_313),
.Y(n_743)
);

BUFx4f_ASAP7_75t_L g744 ( 
.A(n_526),
.Y(n_744)
);

BUFx6f_ASAP7_75t_SL g745 ( 
.A(n_615),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_583),
.B(n_186),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_583),
.B(n_186),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_594),
.B(n_266),
.Y(n_748)
);

NOR3xp33_ASAP7_75t_L g749 ( 
.A(n_518),
.B(n_267),
.C(n_269),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_559),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_564),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_588),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_583),
.B(n_186),
.Y(n_753)
);

O2A1O1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_564),
.A2(n_271),
.B(n_273),
.C(n_284),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_602),
.B(n_186),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_615),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_574),
.B(n_495),
.Y(n_757)
);

O2A1O1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_566),
.A2(n_285),
.B(n_2),
.C(n_5),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_554),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_602),
.B(n_186),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_522),
.B(n_0),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_581),
.B(n_6),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_603),
.B(n_7),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_526),
.B(n_196),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_526),
.B(n_200),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_590),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_615),
.B(n_296),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_483),
.A2(n_294),
.B1(n_292),
.B2(n_286),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_566),
.A2(n_211),
.B1(n_186),
.B2(n_212),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_615),
.B(n_277),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_602),
.B(n_186),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_579),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_572),
.B(n_276),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_611),
.Y(n_774)
);

A2O1A1Ixp33_ASAP7_75t_L g775 ( 
.A1(n_551),
.A2(n_272),
.B(n_258),
.C(n_253),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_551),
.A2(n_211),
.B1(n_212),
.B2(n_239),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_579),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_580),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_R g779 ( 
.A(n_666),
.B(n_575),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_646),
.B(n_482),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_676),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_635),
.A2(n_610),
.B1(n_599),
.B2(n_586),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_627),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_654),
.B(n_476),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_620),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_620),
.Y(n_786)
);

BUFx8_ASAP7_75t_L g787 ( 
.A(n_735),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_663),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_676),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_622),
.Y(n_790)
);

A2O1A1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_762),
.A2(n_552),
.B(n_618),
.C(n_521),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_622),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_628),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_652),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_632),
.Y(n_795)
);

INVx4_ASAP7_75t_L g796 ( 
.A(n_737),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_661),
.B(n_553),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_683),
.B(n_626),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_673),
.Y(n_799)
);

INVx5_ASAP7_75t_L g800 ( 
.A(n_630),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_636),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_671),
.A2(n_575),
.B1(n_538),
.B2(n_616),
.Y(n_802)
);

OAI22xp5_ASAP7_75t_SL g803 ( 
.A1(n_648),
.A2(n_520),
.B1(n_537),
.B2(n_521),
.Y(n_803)
);

A2O1A1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_762),
.A2(n_552),
.B(n_618),
.C(n_610),
.Y(n_804)
);

INVx4_ASAP7_75t_L g805 ( 
.A(n_737),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_SL g806 ( 
.A1(n_736),
.A2(n_575),
.B1(n_537),
.B2(n_582),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_640),
.B(n_580),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_654),
.B(n_476),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_732),
.B(n_641),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_699),
.B(n_558),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_642),
.B(n_584),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_629),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_632),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_724),
.B(n_739),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_633),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_643),
.B(n_586),
.Y(n_816)
);

AOI221xp5_ASAP7_75t_SL g817 ( 
.A1(n_689),
.A2(n_617),
.B1(n_549),
.B2(n_545),
.C(n_543),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_681),
.Y(n_818)
);

BUFx8_ASAP7_75t_L g819 ( 
.A(n_745),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_638),
.A2(n_613),
.B1(n_595),
.B2(n_599),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_655),
.B(n_498),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_681),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_SL g823 ( 
.A1(n_720),
.A2(n_222),
.B1(n_202),
.B2(n_203),
.Y(n_823)
);

BUFx4f_ASAP7_75t_L g824 ( 
.A(n_737),
.Y(n_824)
);

NAND2x1p5_ASAP7_75t_L g825 ( 
.A(n_744),
.B(n_498),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_657),
.B(n_595),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_634),
.A2(n_498),
.B1(n_602),
.B2(n_545),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_774),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_744),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_637),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_634),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_639),
.B(n_604),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_725),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_644),
.Y(n_834)
);

NOR2x1p5_ASAP7_75t_L g835 ( 
.A(n_701),
.B(n_612),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_639),
.B(n_471),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_645),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_649),
.B(n_471),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_706),
.Y(n_839)
);

NAND2x1p5_ASAP7_75t_L g840 ( 
.A(n_663),
.B(n_498),
.Y(n_840)
);

OR2x4_ASAP7_75t_L g841 ( 
.A(n_761),
.B(n_543),
.Y(n_841)
);

OR2x6_ASAP7_75t_L g842 ( 
.A(n_664),
.B(n_515),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_653),
.Y(n_843)
);

INVx4_ASAP7_75t_L g844 ( 
.A(n_745),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_728),
.B(n_474),
.Y(n_845)
);

BUFx4f_ASAP7_75t_L g846 ( 
.A(n_664),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_647),
.B(n_479),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_756),
.B(n_549),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_700),
.B(n_479),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_660),
.B(n_476),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_664),
.B(n_612),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_704),
.B(n_708),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_680),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_761),
.A2(n_607),
.B1(n_508),
.B2(n_499),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_669),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_709),
.B(n_631),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_670),
.B(n_490),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_672),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_677),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_707),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_731),
.Y(n_861)
);

INVx4_ASAP7_75t_L g862 ( 
.A(n_725),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_678),
.B(n_491),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_698),
.B(n_612),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_679),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_686),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_692),
.B(n_693),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_660),
.B(n_476),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_667),
.Y(n_869)
);

OR2x2_ASAP7_75t_SL g870 ( 
.A(n_730),
.B(n_715),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_725),
.Y(n_871)
);

INVx1_ASAP7_75t_SL g872 ( 
.A(n_621),
.Y(n_872)
);

OR2x2_ASAP7_75t_L g873 ( 
.A(n_748),
.B(n_570),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_703),
.B(n_705),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_695),
.A2(n_493),
.B1(n_607),
.B2(n_501),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_749),
.B(n_612),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_651),
.B(n_499),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_717),
.B(n_713),
.Y(n_878)
);

AND2x6_ASAP7_75t_L g879 ( 
.A(n_717),
.B(n_476),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_725),
.Y(n_880)
);

AND2x2_ASAP7_75t_SL g881 ( 
.A(n_729),
.B(n_496),
.Y(n_881)
);

OR2x4_ASAP7_75t_L g882 ( 
.A(n_763),
.B(n_496),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_767),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_714),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_718),
.B(n_570),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_741),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_719),
.B(n_496),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_723),
.B(n_571),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_741),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_741),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_763),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_690),
.B(n_571),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_695),
.A2(n_757),
.B1(n_729),
.B2(n_694),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_659),
.B(n_501),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_740),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_758),
.A2(n_530),
.B(n_577),
.C(n_503),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_733),
.Y(n_897)
);

BUFx2_ASAP7_75t_SL g898 ( 
.A(n_630),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_682),
.B(n_503),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_741),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_682),
.B(n_507),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_684),
.A2(n_507),
.B1(n_508),
.B2(n_510),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_623),
.B(n_496),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_684),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_624),
.B(n_496),
.Y(n_905)
);

NOR2xp67_ASAP7_75t_L g906 ( 
.A(n_770),
.B(n_577),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_766),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_716),
.B(n_722),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_766),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_711),
.B(n_530),
.Y(n_910)
);

OAI22xp33_ASAP7_75t_L g911 ( 
.A1(n_727),
.A2(n_563),
.B1(n_510),
.B2(n_569),
.Y(n_911)
);

BUFx4f_ASAP7_75t_L g912 ( 
.A(n_630),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_625),
.Y(n_913)
);

INVx5_ASAP7_75t_L g914 ( 
.A(n_630),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_630),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_734),
.B(n_563),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_619),
.A2(n_569),
.B1(n_486),
.B2(n_500),
.Y(n_917)
);

INVx1_ASAP7_75t_SL g918 ( 
.A(n_764),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_750),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_743),
.B(n_534),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_662),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_SL g922 ( 
.A(n_765),
.B(n_515),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_751),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_665),
.B(n_534),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_694),
.A2(n_587),
.B1(n_582),
.B2(n_515),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_650),
.B(n_531),
.Y(n_926)
);

INVx1_ASAP7_75t_SL g927 ( 
.A(n_773),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_R g928 ( 
.A(n_658),
.B(n_515),
.Y(n_928)
);

NOR2x2_ASAP7_75t_L g929 ( 
.A(n_668),
.B(n_13),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_752),
.B(n_534),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_778),
.B(n_534),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_697),
.B(n_531),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_738),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_685),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_702),
.B(n_504),
.Y(n_935)
);

INVx5_ASAP7_75t_L g936 ( 
.A(n_759),
.Y(n_936)
);

INVx1_ASAP7_75t_SL g937 ( 
.A(n_687),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_772),
.B(n_565),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_702),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_772),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_777),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_777),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_778),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_712),
.B(n_587),
.Y(n_944)
);

NAND3xp33_ASAP7_75t_SL g945 ( 
.A(n_754),
.B(n_206),
.C(n_213),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_798),
.B(n_768),
.Y(n_946)
);

A2O1A1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_891),
.A2(n_710),
.B(n_742),
.C(n_775),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_787),
.Y(n_948)
);

OAI21x1_ASAP7_75t_L g949 ( 
.A1(n_887),
.A2(n_746),
.B(n_747),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_831),
.B(n_918),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_783),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_852),
.A2(n_710),
.B(n_742),
.C(n_775),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_816),
.A2(n_753),
.B(n_771),
.Y(n_953)
);

OR2x2_ASAP7_75t_L g954 ( 
.A(n_794),
.B(n_696),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_831),
.B(n_656),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_829),
.B(n_844),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_845),
.A2(n_746),
.B(n_753),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_908),
.B(n_656),
.Y(n_958)
);

AOI221xp5_ASAP7_75t_L g959 ( 
.A1(n_797),
.A2(n_726),
.B1(n_776),
.B2(n_721),
.C(n_769),
.Y(n_959)
);

INVxp67_ASAP7_75t_L g960 ( 
.A(n_859),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_839),
.A2(n_760),
.B(n_755),
.C(n_726),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_787),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_824),
.B(n_565),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_927),
.B(n_688),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_869),
.B(n_755),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_819),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_869),
.B(n_809),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_881),
.A2(n_691),
.B1(n_776),
.B2(n_760),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_812),
.Y(n_969)
);

INVx6_ASAP7_75t_L g970 ( 
.A(n_819),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_818),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_809),
.B(n_674),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_904),
.A2(n_675),
.B1(n_721),
.B2(n_565),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_793),
.B(n_486),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_815),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_779),
.Y(n_976)
);

INVx6_ASAP7_75t_L g977 ( 
.A(n_844),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_872),
.B(n_485),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_779),
.B(n_565),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_838),
.B(n_531),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_847),
.A2(n_587),
.B(n_582),
.Y(n_981)
);

OAI21x1_ASAP7_75t_SL g982 ( 
.A1(n_867),
.A2(n_769),
.B(n_18),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_814),
.B(n_477),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_802),
.B(n_500),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_822),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_883),
.B(n_531),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_821),
.B(n_856),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_780),
.B(n_485),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_896),
.A2(n_504),
.B(n_22),
.C(n_23),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_801),
.B(n_504),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_894),
.A2(n_901),
.B(n_899),
.C(n_893),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_801),
.B(n_220),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_811),
.B(n_568),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_781),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_830),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_896),
.A2(n_17),
.B(n_22),
.C(n_25),
.Y(n_996)
);

OR2x6_ASAP7_75t_SL g997 ( 
.A(n_799),
.B(n_221),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_826),
.B(n_568),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_915),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_874),
.A2(n_17),
.B(n_25),
.C(n_29),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_834),
.B(n_568),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_893),
.A2(n_232),
.B1(n_243),
.B2(n_247),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_939),
.A2(n_29),
.B(n_30),
.C(n_32),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_910),
.A2(n_878),
.B(n_920),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_892),
.B(n_30),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_841),
.B(n_36),
.Y(n_1006)
);

CKINVDCx16_ASAP7_75t_R g1007 ( 
.A(n_823),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_915),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_SL g1009 ( 
.A(n_881),
.B(n_796),
.Y(n_1009)
);

AO21x1_ASAP7_75t_L g1010 ( 
.A1(n_901),
.A2(n_911),
.B(n_808),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_837),
.B(n_547),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_843),
.B(n_547),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_935),
.A2(n_547),
.B(n_212),
.C(n_40),
.Y(n_1013)
);

INVx4_ASAP7_75t_L g1014 ( 
.A(n_879),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_855),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_882),
.Y(n_1016)
);

INVx2_ASAP7_75t_SL g1017 ( 
.A(n_828),
.Y(n_1017)
);

O2A1O1Ixp5_ASAP7_75t_L g1018 ( 
.A1(n_804),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_1018)
);

NOR3xp33_ASAP7_75t_L g1019 ( 
.A(n_945),
.B(n_39),
.C(n_42),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_781),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_796),
.B(n_547),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_935),
.A2(n_212),
.B(n_45),
.C(n_46),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_805),
.B(n_212),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_945),
.A2(n_43),
.B(n_47),
.C(n_48),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_870),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_858),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_865),
.A2(n_43),
.B1(n_47),
.B2(n_48),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_805),
.B(n_49),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_842),
.B(n_50),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_919),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_841),
.B(n_50),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_866),
.B(n_51),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_853),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_781),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_887),
.A2(n_112),
.B(n_78),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_912),
.B(n_54),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_884),
.B(n_94),
.Y(n_1037)
);

AND2x6_ASAP7_75t_L g1038 ( 
.A(n_851),
.B(n_864),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_849),
.A2(n_832),
.B(n_836),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_916),
.A2(n_924),
.B(n_930),
.Y(n_1040)
);

AO22x1_ASAP7_75t_L g1041 ( 
.A1(n_864),
.A2(n_98),
.B1(n_104),
.B2(n_109),
.Y(n_1041)
);

NOR2xp67_ASAP7_75t_L g1042 ( 
.A(n_895),
.B(n_110),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_810),
.B(n_128),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_R g1044 ( 
.A(n_846),
.B(n_134),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_923),
.A2(n_135),
.B1(n_148),
.B2(n_153),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_781),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_800),
.A2(n_914),
.B1(n_807),
.B2(n_784),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_882),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_R g1049 ( 
.A(n_846),
.B(n_880),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_930),
.A2(n_857),
.B(n_863),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_842),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_913),
.B(n_803),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_860),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_842),
.B(n_851),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_804),
.A2(n_903),
.B(n_905),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_835),
.B(n_934),
.Y(n_1056)
);

BUFx8_ASAP7_75t_L g1057 ( 
.A(n_879),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_940),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_848),
.A2(n_791),
.B(n_868),
.C(n_784),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_861),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_785),
.B(n_786),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_850),
.A2(n_868),
.B(n_873),
.C(n_906),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_800),
.A2(n_914),
.B1(n_850),
.B2(n_782),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_825),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_932),
.Y(n_1065)
);

NAND2x1p5_ASAP7_75t_L g1066 ( 
.A(n_800),
.B(n_914),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_937),
.B(n_941),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_943),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_909),
.B(n_921),
.Y(n_1069)
);

AND2x6_ASAP7_75t_L g1070 ( 
.A(n_788),
.B(n_833),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_903),
.A2(n_905),
.B(n_944),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_800),
.A2(n_914),
.B1(n_782),
.B2(n_898),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_825),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_SL g1074 ( 
.A1(n_827),
.A2(n_880),
.B(n_917),
.C(n_888),
.Y(n_1074)
);

AOI21x1_ASAP7_75t_L g1075 ( 
.A1(n_931),
.A2(n_938),
.B(n_885),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_926),
.A2(n_788),
.B(n_922),
.Y(n_1076)
);

INVx5_ASAP7_75t_L g1077 ( 
.A(n_1014),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_946),
.A2(n_854),
.B(n_875),
.Y(n_1078)
);

O2A1O1Ixp5_ASAP7_75t_SL g1079 ( 
.A1(n_984),
.A2(n_1028),
.B(n_1027),
.C(n_987),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_SL g1080 ( 
.A1(n_1072),
.A2(n_833),
.B(n_932),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_950),
.B(n_813),
.Y(n_1081)
);

OAI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1002),
.A2(n_875),
.B(n_902),
.Y(n_1082)
);

BUFx12f_ASAP7_75t_L g1083 ( 
.A(n_970),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1002),
.A2(n_817),
.B(n_806),
.Y(n_1084)
);

AO31x2_ASAP7_75t_L g1085 ( 
.A1(n_1010),
.A2(n_795),
.A3(n_792),
.B(n_790),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_951),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_967),
.B(n_942),
.Y(n_1087)
);

INVxp67_ASAP7_75t_L g1088 ( 
.A(n_971),
.Y(n_1088)
);

AOI221x1_ASAP7_75t_L g1089 ( 
.A1(n_1019),
.A2(n_921),
.B1(n_933),
.B2(n_877),
.C(n_897),
.Y(n_1089)
);

AO22x1_ASAP7_75t_L g1090 ( 
.A1(n_1057),
.A2(n_876),
.B1(n_929),
.B2(n_879),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_1059),
.A2(n_925),
.B(n_820),
.C(n_907),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_960),
.A2(n_820),
.B1(n_925),
.B2(n_936),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_1063),
.B(n_789),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1005),
.B(n_929),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_1067),
.B(n_921),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_1063),
.B(n_789),
.Y(n_1096)
);

NOR2xp67_ASAP7_75t_L g1097 ( 
.A(n_976),
.B(n_862),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_SL g1098 ( 
.A1(n_1027),
.A2(n_840),
.B(n_789),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_964),
.B(n_921),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_991),
.A2(n_936),
.B(n_789),
.C(n_889),
.Y(n_1100)
);

AO21x1_ASAP7_75t_L g1101 ( 
.A1(n_1047),
.A2(n_862),
.B(n_840),
.Y(n_1101)
);

INVx4_ASAP7_75t_L g1102 ( 
.A(n_1014),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1052),
.B(n_879),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_972),
.B(n_958),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_983),
.B(n_879),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_SL g1106 ( 
.A1(n_1062),
.A2(n_871),
.B(n_886),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_988),
.B(n_936),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_953),
.A2(n_957),
.B(n_952),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_958),
.B(n_936),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1025),
.B(n_871),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_996),
.A2(n_871),
.B(n_886),
.C(n_889),
.Y(n_1111)
);

AO21x2_ASAP7_75t_L g1112 ( 
.A1(n_1071),
.A2(n_928),
.B(n_889),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_969),
.B(n_886),
.Y(n_1113)
);

NOR2x1_ASAP7_75t_SL g1114 ( 
.A(n_994),
.B(n_889),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1074),
.A2(n_1076),
.B(n_1004),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_975),
.B(n_890),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_985),
.Y(n_1117)
);

NAND3xp33_ASAP7_75t_SL g1118 ( 
.A(n_1024),
.B(n_928),
.C(n_890),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_1065),
.Y(n_1119)
);

NAND2x1p5_ASAP7_75t_L g1120 ( 
.A(n_1054),
.B(n_890),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_995),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1015),
.B(n_1026),
.Y(n_1122)
);

OA21x2_ASAP7_75t_L g1123 ( 
.A1(n_1055),
.A2(n_900),
.B(n_981),
.Y(n_1123)
);

NOR2xp67_ASAP7_75t_SL g1124 ( 
.A(n_948),
.B(n_900),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1075),
.A2(n_900),
.B(n_949),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_955),
.A2(n_947),
.B(n_978),
.Y(n_1126)
);

NAND3xp33_ASAP7_75t_L g1127 ( 
.A(n_1022),
.B(n_1000),
.C(n_1031),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_980),
.A2(n_1050),
.B(n_1047),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_954),
.B(n_1043),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1035),
.A2(n_980),
.B(n_1066),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1029),
.B(n_1030),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1006),
.A2(n_989),
.B(n_959),
.C(n_1018),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_992),
.A2(n_990),
.B1(n_1032),
.B2(n_1029),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_965),
.A2(n_961),
.B(n_974),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1056),
.B(n_1038),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1038),
.B(n_1054),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1058),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_1051),
.A2(n_993),
.B(n_998),
.Y(n_1138)
);

AOI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1023),
.A2(n_1041),
.B(n_979),
.Y(n_1139)
);

AOI21x1_ASAP7_75t_L g1140 ( 
.A1(n_963),
.A2(n_1048),
.B(n_1016),
.Y(n_1140)
);

AOI221xp5_ASAP7_75t_SL g1141 ( 
.A1(n_1003),
.A2(n_1013),
.B1(n_1036),
.B2(n_1045),
.C(n_986),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_997),
.B(n_1017),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1068),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_962),
.B(n_956),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_1045),
.A2(n_1042),
.B(n_1037),
.C(n_968),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1064),
.A2(n_1073),
.B(n_999),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1038),
.B(n_956),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1038),
.B(n_1049),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_973),
.A2(n_1069),
.B(n_1009),
.C(n_1008),
.Y(n_1149)
);

NOR2xp67_ASAP7_75t_SL g1150 ( 
.A(n_966),
.B(n_970),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1001),
.A2(n_1011),
.B(n_1012),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1070),
.A2(n_1061),
.B(n_1021),
.Y(n_1152)
);

OAI21xp33_ASAP7_75t_SL g1153 ( 
.A1(n_1061),
.A2(n_1057),
.B(n_1060),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1070),
.A2(n_1053),
.B(n_1033),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_994),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_994),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_977),
.B(n_1070),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1020),
.A2(n_1034),
.B(n_1046),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_1020),
.A2(n_1034),
.B(n_1046),
.C(n_1044),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_977),
.B(n_1034),
.Y(n_1160)
);

NOR3xp33_ASAP7_75t_L g1161 ( 
.A(n_1046),
.B(n_635),
.C(n_946),
.Y(n_1161)
);

BUFx4_ASAP7_75t_SL g1162 ( 
.A(n_948),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1040),
.A2(n_1075),
.B(n_1055),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_1030),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_SL g1165 ( 
.A1(n_1072),
.A2(n_1014),
.B(n_1063),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_950),
.B(n_798),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1039),
.A2(n_635),
.B(n_912),
.Y(n_1167)
);

A2O1A1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_946),
.A2(n_635),
.B(n_1059),
.C(n_991),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_946),
.A2(n_635),
.B1(n_661),
.B2(n_831),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1040),
.A2(n_1075),
.B(n_1055),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1040),
.A2(n_1075),
.B(n_1055),
.Y(n_1171)
);

NAND2x1p5_ASAP7_75t_L g1172 ( 
.A(n_1014),
.B(n_824),
.Y(n_1172)
);

INVx2_ASAP7_75t_SL g1173 ( 
.A(n_977),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_948),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_1054),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_SL g1176 ( 
.A1(n_1072),
.A2(n_1014),
.B(n_1063),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1039),
.A2(n_635),
.B(n_912),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_946),
.A2(n_635),
.B(n_661),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_SL g1179 ( 
.A1(n_955),
.A2(n_989),
.B(n_982),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_950),
.B(n_798),
.Y(n_1180)
);

CKINVDCx6p67_ASAP7_75t_R g1181 ( 
.A(n_948),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1039),
.A2(n_635),
.B(n_912),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_950),
.B(n_798),
.Y(n_1183)
);

INVxp67_ASAP7_75t_SL g1184 ( 
.A(n_1072),
.Y(n_1184)
);

AOI221x1_ASAP7_75t_L g1185 ( 
.A1(n_1019),
.A2(n_1022),
.B1(n_991),
.B2(n_1002),
.C(n_947),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_946),
.A2(n_635),
.B1(n_661),
.B2(n_831),
.Y(n_1186)
);

CKINVDCx11_ASAP7_75t_R g1187 ( 
.A(n_997),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_1065),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_1030),
.Y(n_1189)
);

OR2x6_ASAP7_75t_L g1190 ( 
.A(n_1014),
.B(n_844),
.Y(n_1190)
);

NOR2x1_ASAP7_75t_SL g1191 ( 
.A(n_1014),
.B(n_737),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1040),
.A2(n_1075),
.B(n_1055),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_946),
.B(n_661),
.Y(n_1193)
);

XNOR2xp5_ASAP7_75t_L g1194 ( 
.A(n_962),
.B(n_550),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1039),
.A2(n_635),
.B(n_912),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_951),
.Y(n_1196)
);

OAI22x1_ASAP7_75t_L g1197 ( 
.A1(n_1052),
.A2(n_550),
.B1(n_904),
.B2(n_1005),
.Y(n_1197)
);

NOR2xp67_ASAP7_75t_L g1198 ( 
.A(n_976),
.B(n_666),
.Y(n_1198)
);

NOR2x1_ASAP7_75t_SL g1199 ( 
.A(n_1014),
.B(n_737),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_1065),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_948),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1039),
.A2(n_635),
.B(n_912),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_950),
.B(n_798),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_950),
.B(n_798),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1193),
.B(n_1166),
.Y(n_1205)
);

O2A1O1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1168),
.A2(n_1193),
.B(n_1178),
.C(n_1186),
.Y(n_1206)
);

OAI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1169),
.A2(n_1185),
.B1(n_1184),
.B2(n_1203),
.Y(n_1207)
);

CKINVDCx16_ASAP7_75t_R g1208 ( 
.A(n_1083),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1168),
.A2(n_1145),
.B(n_1161),
.Y(n_1209)
);

NOR2x1_ASAP7_75t_L g1210 ( 
.A(n_1198),
.B(n_1097),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1122),
.Y(n_1211)
);

INVx5_ASAP7_75t_L g1212 ( 
.A(n_1190),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1085),
.Y(n_1213)
);

AO21x2_ASAP7_75t_L g1214 ( 
.A1(n_1084),
.A2(n_1145),
.B(n_1151),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1192),
.A2(n_1115),
.B(n_1138),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1180),
.B(n_1204),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1125),
.A2(n_1128),
.B(n_1130),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1183),
.B(n_1104),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1086),
.Y(n_1219)
);

O2A1O1Ixp33_ASAP7_75t_SL g1220 ( 
.A1(n_1132),
.A2(n_1111),
.B(n_1100),
.C(n_1103),
.Y(n_1220)
);

CKINVDCx12_ASAP7_75t_R g1221 ( 
.A(n_1131),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1104),
.B(n_1129),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1121),
.Y(n_1223)
);

CKINVDCx6p67_ASAP7_75t_R g1224 ( 
.A(n_1187),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1119),
.B(n_1188),
.Y(n_1225)
);

O2A1O1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1133),
.A2(n_1132),
.B(n_1127),
.C(n_1078),
.Y(n_1226)
);

O2A1O1Ixp33_ASAP7_75t_SL g1227 ( 
.A1(n_1111),
.A2(n_1159),
.B(n_1091),
.C(n_1126),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1167),
.A2(n_1202),
.B(n_1182),
.Y(n_1228)
);

OAI222xp33_ASAP7_75t_L g1229 ( 
.A1(n_1184),
.A2(n_1092),
.B1(n_1081),
.B2(n_1109),
.C1(n_1099),
.C2(n_1087),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1085),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1177),
.A2(n_1195),
.B(n_1079),
.Y(n_1231)
);

OAI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1197),
.A2(n_1082),
.B1(n_1098),
.B2(n_1088),
.Y(n_1232)
);

INVx4_ASAP7_75t_L g1233 ( 
.A(n_1174),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1088),
.B(n_1119),
.Y(n_1234)
);

BUFx10_ASAP7_75t_L g1235 ( 
.A(n_1201),
.Y(n_1235)
);

NAND2x1p5_ASAP7_75t_L g1236 ( 
.A(n_1077),
.B(n_1102),
.Y(n_1236)
);

OR2x2_ASAP7_75t_L g1237 ( 
.A(n_1188),
.B(n_1200),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_1187),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1090),
.A2(n_1150),
.B1(n_1194),
.B2(n_1142),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1200),
.B(n_1095),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1165),
.A2(n_1176),
.B(n_1106),
.Y(n_1241)
);

CKINVDCx16_ASAP7_75t_R g1242 ( 
.A(n_1110),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1117),
.B(n_1196),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1093),
.A2(n_1096),
.B(n_1080),
.Y(n_1244)
);

AO31x2_ASAP7_75t_L g1245 ( 
.A1(n_1089),
.A2(n_1091),
.A3(n_1149),
.B(n_1101),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1123),
.A2(n_1139),
.B(n_1179),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1175),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1085),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1137),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1093),
.A2(n_1096),
.B(n_1134),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1143),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1085),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1118),
.A2(n_1153),
.B1(n_1135),
.B2(n_1117),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1105),
.A2(n_1107),
.B1(n_1164),
.B2(n_1189),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1190),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1120),
.B(n_1157),
.Y(n_1256)
);

OAI222xp33_ASAP7_75t_L g1257 ( 
.A1(n_1147),
.A2(n_1148),
.B1(n_1136),
.B2(n_1113),
.C1(n_1116),
.C2(n_1190),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1123),
.A2(n_1146),
.B(n_1152),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1118),
.A2(n_1112),
.B(n_1077),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1162),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_1162),
.Y(n_1261)
);

AO21x2_ASAP7_75t_L g1262 ( 
.A1(n_1154),
.A2(n_1140),
.B(n_1159),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1112),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_SL g1264 ( 
.A(n_1181),
.B(n_1124),
.Y(n_1264)
);

O2A1O1Ixp33_ASAP7_75t_SL g1265 ( 
.A1(n_1155),
.A2(n_1156),
.B(n_1158),
.C(n_1141),
.Y(n_1265)
);

A2O1A1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1077),
.A2(n_1144),
.B(n_1160),
.C(n_1173),
.Y(n_1266)
);

AO21x2_ASAP7_75t_L g1267 ( 
.A1(n_1191),
.A2(n_1199),
.B(n_1114),
.Y(n_1267)
);

OAI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1175),
.A2(n_1102),
.B1(n_1172),
.B2(n_1120),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1172),
.A2(n_1193),
.B(n_1168),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1175),
.A2(n_1193),
.B1(n_1178),
.B2(n_1186),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1193),
.A2(n_1168),
.B(n_1178),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1168),
.A2(n_1177),
.B(n_1167),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1193),
.A2(n_1197),
.B1(n_1005),
.B2(n_881),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1163),
.A2(n_1171),
.B(n_1170),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1163),
.A2(n_1171),
.B(n_1170),
.Y(n_1275)
);

AOI221xp5_ASAP7_75t_L g1276 ( 
.A1(n_1178),
.A2(n_541),
.B1(n_1193),
.B2(n_1186),
.C(n_1169),
.Y(n_1276)
);

CKINVDCx8_ASAP7_75t_R g1277 ( 
.A(n_1174),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1163),
.A2(n_1171),
.B(n_1170),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1136),
.B(n_1051),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1163),
.A2(n_1171),
.B(n_1170),
.Y(n_1280)
);

OAI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1193),
.A2(n_1168),
.B(n_1178),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1163),
.A2(n_1171),
.B(n_1170),
.Y(n_1282)
);

NOR2x1_ASAP7_75t_L g1283 ( 
.A(n_1198),
.B(n_1097),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1122),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1163),
.A2(n_1171),
.B(n_1170),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1193),
.A2(n_1168),
.B(n_1178),
.Y(n_1286)
);

AOI222xp33_ASAP7_75t_L g1287 ( 
.A1(n_1193),
.A2(n_720),
.B1(n_261),
.B2(n_274),
.C1(n_288),
.C2(n_234),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1122),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1122),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1193),
.A2(n_1197),
.B1(n_1005),
.B2(n_881),
.Y(n_1290)
);

NAND2x1p5_ASAP7_75t_L g1291 ( 
.A(n_1077),
.B(n_1014),
.Y(n_1291)
);

NOR2x1_ASAP7_75t_L g1292 ( 
.A(n_1198),
.B(n_1097),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1136),
.B(n_1051),
.Y(n_1293)
);

CKINVDCx20_ASAP7_75t_R g1294 ( 
.A(n_1187),
.Y(n_1294)
);

BUFx2_ASAP7_75t_SL g1295 ( 
.A(n_1198),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1193),
.A2(n_1197),
.B1(n_1005),
.B2(n_881),
.Y(n_1296)
);

OAI221xp5_ASAP7_75t_L g1297 ( 
.A1(n_1178),
.A2(n_1193),
.B1(n_698),
.B2(n_556),
.C(n_535),
.Y(n_1297)
);

INVx4_ASAP7_75t_L g1298 ( 
.A(n_1083),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1122),
.Y(n_1299)
);

NAND3xp33_ASAP7_75t_L g1300 ( 
.A(n_1193),
.B(n_1168),
.C(n_1178),
.Y(n_1300)
);

NAND2x1p5_ASAP7_75t_L g1301 ( 
.A(n_1077),
.B(n_1014),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1193),
.B(n_1166),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1085),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1164),
.Y(n_1304)
);

INVx2_ASAP7_75t_SL g1305 ( 
.A(n_1162),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1193),
.A2(n_1178),
.B1(n_1186),
.B2(n_1169),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_SL g1307 ( 
.A1(n_1179),
.A2(n_1133),
.B(n_1103),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1122),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1193),
.B(n_1169),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1164),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_1187),
.Y(n_1311)
);

INVx2_ASAP7_75t_SL g1312 ( 
.A(n_1162),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1193),
.A2(n_1168),
.B(n_1178),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_SL g1314 ( 
.A1(n_1184),
.A2(n_881),
.B1(n_1129),
.B2(n_342),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1193),
.B(n_1094),
.Y(n_1315)
);

OA21x2_ASAP7_75t_L g1316 ( 
.A1(n_1108),
.A2(n_1170),
.B(n_1163),
.Y(n_1316)
);

AO21x1_ASAP7_75t_L g1317 ( 
.A1(n_1133),
.A2(n_1126),
.B(n_1084),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1193),
.B(n_1166),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1193),
.B(n_1094),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1163),
.A2(n_1171),
.B(n_1170),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1163),
.A2(n_1171),
.B(n_1170),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1193),
.A2(n_535),
.B1(n_1052),
.B2(n_1007),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1163),
.A2(n_1171),
.B(n_1170),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1193),
.B(n_1094),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1162),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1085),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1162),
.Y(n_1327)
);

O2A1O1Ixp33_ASAP7_75t_SL g1328 ( 
.A1(n_1168),
.A2(n_1145),
.B(n_1132),
.C(n_1178),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1219),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1222),
.B(n_1309),
.Y(n_1330)
);

O2A1O1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1306),
.A2(n_1206),
.B(n_1281),
.C(n_1286),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1309),
.B(n_1205),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1300),
.A2(n_1322),
.B1(n_1276),
.B2(n_1297),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1271),
.A2(n_1313),
.B1(n_1206),
.B2(n_1270),
.Y(n_1334)
);

O2A1O1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1328),
.A2(n_1226),
.B(n_1207),
.C(n_1209),
.Y(n_1335)
);

AOI21x1_ASAP7_75t_SL g1336 ( 
.A1(n_1234),
.A2(n_1318),
.B(n_1302),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1218),
.B(n_1233),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1328),
.A2(n_1272),
.B(n_1241),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1216),
.B(n_1211),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1223),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1207),
.A2(n_1314),
.B1(n_1226),
.B2(n_1269),
.Y(n_1341)
);

O2A1O1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1317),
.A2(n_1232),
.B(n_1227),
.C(n_1220),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1314),
.A2(n_1232),
.B1(n_1273),
.B2(n_1296),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1319),
.B(n_1324),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1228),
.A2(n_1220),
.B(n_1214),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1237),
.B(n_1240),
.Y(n_1346)
);

A2O1A1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1244),
.A2(n_1250),
.B(n_1296),
.C(n_1273),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1316),
.Y(n_1348)
);

BUFx8_ASAP7_75t_L g1349 ( 
.A(n_1260),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1290),
.A2(n_1253),
.B1(n_1304),
.B2(n_1310),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1290),
.A2(n_1253),
.B1(n_1239),
.B2(n_1295),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1242),
.B(n_1243),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_SL g1353 ( 
.A1(n_1266),
.A2(n_1291),
.B(n_1301),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1254),
.A2(n_1238),
.B1(n_1294),
.B2(n_1311),
.Y(n_1354)
);

A2O1A1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1259),
.A2(n_1266),
.B(n_1210),
.C(n_1283),
.Y(n_1355)
);

O2A1O1Ixp5_ASAP7_75t_L g1356 ( 
.A1(n_1229),
.A2(n_1257),
.B(n_1268),
.C(n_1230),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1284),
.B(n_1288),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1289),
.B(n_1299),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1308),
.B(n_1249),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1251),
.B(n_1279),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1212),
.B(n_1279),
.Y(n_1361)
);

O2A1O1Ixp5_ASAP7_75t_L g1362 ( 
.A1(n_1229),
.A2(n_1257),
.B(n_1268),
.C(n_1326),
.Y(n_1362)
);

CKINVDCx20_ASAP7_75t_R g1363 ( 
.A(n_1238),
.Y(n_1363)
);

O2A1O1Ixp5_ASAP7_75t_L g1364 ( 
.A1(n_1213),
.A2(n_1248),
.B(n_1326),
.C(n_1230),
.Y(n_1364)
);

O2A1O1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1287),
.A2(n_1307),
.B(n_1265),
.C(n_1264),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1294),
.A2(n_1311),
.B1(n_1224),
.B2(n_1305),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1293),
.B(n_1256),
.Y(n_1367)
);

O2A1O1Ixp5_ASAP7_75t_L g1368 ( 
.A1(n_1213),
.A2(n_1252),
.B(n_1248),
.C(n_1303),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1212),
.B(n_1293),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1247),
.B(n_1255),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1292),
.Y(n_1371)
);

O2A1O1Ixp5_ASAP7_75t_L g1372 ( 
.A1(n_1252),
.A2(n_1303),
.B(n_1263),
.C(n_1298),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1312),
.A2(n_1327),
.B1(n_1325),
.B2(n_1261),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1208),
.B(n_1245),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1233),
.B(n_1325),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1261),
.A2(n_1327),
.B1(n_1298),
.B2(n_1236),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1236),
.A2(n_1277),
.B1(n_1263),
.B2(n_1221),
.Y(n_1377)
);

O2A1O1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1262),
.A2(n_1267),
.B(n_1245),
.C(n_1235),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1246),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1245),
.B(n_1235),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1245),
.B(n_1258),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1274),
.B(n_1275),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1278),
.A2(n_1280),
.B1(n_1282),
.B2(n_1285),
.Y(n_1383)
);

AOI21x1_ASAP7_75t_SL g1384 ( 
.A1(n_1320),
.A2(n_1321),
.B(n_1323),
.Y(n_1384)
);

NOR2xp67_ASAP7_75t_L g1385 ( 
.A(n_1241),
.B(n_1239),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_SL g1386 ( 
.A1(n_1226),
.A2(n_1168),
.B(n_1145),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1315),
.B(n_1319),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1237),
.B(n_1240),
.Y(n_1388)
);

NOR2xp67_ASAP7_75t_L g1389 ( 
.A(n_1241),
.B(n_1239),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1237),
.B(n_1240),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1309),
.A2(n_1193),
.B1(n_1300),
.B2(n_1322),
.Y(n_1391)
);

O2A1O1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1306),
.A2(n_1168),
.B(n_1206),
.C(n_1271),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1222),
.B(n_1309),
.Y(n_1393)
);

O2A1O1Ixp33_ASAP7_75t_L g1394 ( 
.A1(n_1306),
.A2(n_1168),
.B(n_1206),
.C(n_1271),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1328),
.A2(n_1168),
.B(n_1272),
.Y(n_1395)
);

O2A1O1Ixp5_ASAP7_75t_L g1396 ( 
.A1(n_1317),
.A2(n_1209),
.B(n_1309),
.C(n_1168),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1222),
.B(n_1309),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1225),
.B(n_1310),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1219),
.Y(n_1399)
);

OR2x6_ASAP7_75t_SL g1400 ( 
.A(n_1261),
.B(n_1325),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1231),
.A2(n_1217),
.B(n_1215),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1309),
.A2(n_1193),
.B1(n_1300),
.B2(n_1322),
.Y(n_1402)
);

O2A1O1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1306),
.A2(n_1168),
.B(n_1206),
.C(n_1271),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1225),
.B(n_1310),
.Y(n_1404)
);

O2A1O1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1306),
.A2(n_1168),
.B(n_1206),
.C(n_1271),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1222),
.B(n_1309),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1222),
.B(n_1309),
.Y(n_1407)
);

O2A1O1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1306),
.A2(n_1168),
.B(n_1206),
.C(n_1271),
.Y(n_1408)
);

OAI31xp33_ASAP7_75t_L g1409 ( 
.A1(n_1297),
.A2(n_1232),
.A3(n_1306),
.B(n_1300),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1225),
.B(n_1310),
.Y(n_1410)
);

BUFx2_ASAP7_75t_L g1411 ( 
.A(n_1379),
.Y(n_1411)
);

NOR3xp33_ASAP7_75t_L g1412 ( 
.A(n_1333),
.B(n_1402),
.C(n_1391),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1329),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1349),
.Y(n_1414)
);

NAND2x1p5_ASAP7_75t_L g1415 ( 
.A(n_1338),
.B(n_1395),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1381),
.B(n_1348),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1330),
.B(n_1393),
.Y(n_1417)
);

AO21x2_ASAP7_75t_L g1418 ( 
.A1(n_1345),
.A2(n_1347),
.B(n_1348),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1340),
.Y(n_1419)
);

NAND3xp33_ASAP7_75t_L g1420 ( 
.A(n_1409),
.B(n_1331),
.C(n_1396),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1380),
.B(n_1345),
.Y(n_1421)
);

OAI321xp33_ASAP7_75t_L g1422 ( 
.A1(n_1341),
.A2(n_1334),
.A3(n_1343),
.B1(n_1331),
.B2(n_1335),
.C(n_1342),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1379),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1344),
.B(n_1387),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1396),
.A2(n_1335),
.B(n_1386),
.Y(n_1425)
);

OA21x2_ASAP7_75t_L g1426 ( 
.A1(n_1356),
.A2(n_1362),
.B(n_1372),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1364),
.Y(n_1427)
);

AOI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1351),
.A2(n_1332),
.B1(n_1385),
.B2(n_1389),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1399),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1382),
.Y(n_1430)
);

AO21x2_ASAP7_75t_L g1431 ( 
.A1(n_1378),
.A2(n_1392),
.B(n_1408),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1346),
.B(n_1388),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1364),
.Y(n_1433)
);

AO21x1_ASAP7_75t_SL g1434 ( 
.A1(n_1374),
.A2(n_1405),
.B(n_1394),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1368),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1359),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1398),
.Y(n_1437)
);

OR2x6_ASAP7_75t_L g1438 ( 
.A(n_1353),
.B(n_1342),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1390),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1397),
.B(n_1406),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1404),
.B(n_1410),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1349),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1407),
.B(n_1394),
.Y(n_1443)
);

AOI21xp33_ASAP7_75t_L g1444 ( 
.A1(n_1392),
.A2(n_1403),
.B(n_1408),
.Y(n_1444)
);

OA21x2_ASAP7_75t_L g1445 ( 
.A1(n_1356),
.A2(n_1372),
.B(n_1383),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1403),
.A2(n_1405),
.B(n_1401),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1401),
.Y(n_1447)
);

OA21x2_ASAP7_75t_L g1448 ( 
.A1(n_1355),
.A2(n_1360),
.B(n_1339),
.Y(n_1448)
);

OA21x2_ASAP7_75t_L g1449 ( 
.A1(n_1357),
.A2(n_1358),
.B(n_1367),
.Y(n_1449)
);

OA21x2_ASAP7_75t_L g1450 ( 
.A1(n_1370),
.A2(n_1350),
.B(n_1361),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1413),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1443),
.B(n_1352),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1431),
.B(n_1337),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1431),
.B(n_1371),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1449),
.B(n_1416),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1449),
.B(n_1369),
.Y(n_1456)
);

INVxp67_ASAP7_75t_L g1457 ( 
.A(n_1434),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1443),
.B(n_1436),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1413),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1419),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1449),
.B(n_1416),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1450),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1449),
.B(n_1354),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1416),
.B(n_1377),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1421),
.B(n_1375),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1429),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1423),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1421),
.B(n_1400),
.Y(n_1468)
);

AO21x2_ASAP7_75t_L g1469 ( 
.A1(n_1446),
.A2(n_1418),
.B(n_1431),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1421),
.B(n_1384),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1418),
.B(n_1365),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1418),
.B(n_1365),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1431),
.B(n_1336),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1411),
.Y(n_1474)
);

AO22x1_ASAP7_75t_L g1475 ( 
.A1(n_1463),
.A2(n_1425),
.B1(n_1412),
.B2(n_1439),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1451),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1451),
.Y(n_1477)
);

NAND3xp33_ASAP7_75t_L g1478 ( 
.A(n_1471),
.B(n_1412),
.C(n_1420),
.Y(n_1478)
);

NOR2x1_ASAP7_75t_R g1479 ( 
.A(n_1468),
.B(n_1414),
.Y(n_1479)
);

OAI221xp5_ASAP7_75t_L g1480 ( 
.A1(n_1453),
.A2(n_1472),
.B1(n_1471),
.B2(n_1428),
.C(n_1420),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1468),
.B(n_1465),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1451),
.Y(n_1482)
);

AOI221xp5_ASAP7_75t_L g1483 ( 
.A1(n_1471),
.A2(n_1422),
.B1(n_1444),
.B2(n_1446),
.C(n_1425),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1455),
.B(n_1439),
.Y(n_1484)
);

BUFx5_ASAP7_75t_L g1485 ( 
.A(n_1462),
.Y(n_1485)
);

OAI33xp33_ASAP7_75t_L g1486 ( 
.A1(n_1453),
.A2(n_1417),
.A3(n_1440),
.B1(n_1436),
.B2(n_1422),
.B3(n_1366),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1455),
.B(n_1432),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1471),
.A2(n_1434),
.B1(n_1444),
.B2(n_1431),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1455),
.B(n_1432),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1468),
.B(n_1437),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1456),
.B(n_1437),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1458),
.B(n_1417),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1472),
.A2(n_1434),
.B1(n_1428),
.B2(n_1426),
.Y(n_1493)
);

OAI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1457),
.A2(n_1438),
.B1(n_1448),
.B2(n_1440),
.Y(n_1494)
);

INVx4_ASAP7_75t_L g1495 ( 
.A(n_1468),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1457),
.A2(n_1438),
.B1(n_1437),
.B2(n_1415),
.Y(n_1496)
);

NAND3xp33_ASAP7_75t_SL g1497 ( 
.A(n_1472),
.B(n_1363),
.C(n_1415),
.Y(n_1497)
);

OAI221xp5_ASAP7_75t_L g1498 ( 
.A1(n_1453),
.A2(n_1426),
.B1(n_1438),
.B2(n_1445),
.C(n_1436),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1465),
.B(n_1441),
.Y(n_1499)
);

A2O1A1Ixp33_ASAP7_75t_L g1500 ( 
.A1(n_1472),
.A2(n_1435),
.B(n_1427),
.C(n_1433),
.Y(n_1500)
);

AO21x2_ASAP7_75t_L g1501 ( 
.A1(n_1469),
.A2(n_1447),
.B(n_1418),
.Y(n_1501)
);

NOR2xp67_ASAP7_75t_L g1502 ( 
.A(n_1455),
.B(n_1456),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_SL g1503 ( 
.A1(n_1462),
.A2(n_1426),
.B1(n_1450),
.B2(n_1438),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1464),
.B(n_1432),
.Y(n_1504)
);

NOR2xp67_ASAP7_75t_L g1505 ( 
.A(n_1456),
.B(n_1430),
.Y(n_1505)
);

NOR2x1_ASAP7_75t_L g1506 ( 
.A(n_1452),
.B(n_1438),
.Y(n_1506)
);

OAI33xp33_ASAP7_75t_L g1507 ( 
.A1(n_1454),
.A2(n_1452),
.A3(n_1473),
.B1(n_1459),
.B2(n_1466),
.B3(n_1460),
.Y(n_1507)
);

AO21x2_ASAP7_75t_L g1508 ( 
.A1(n_1469),
.A2(n_1454),
.B(n_1473),
.Y(n_1508)
);

NAND3xp33_ASAP7_75t_L g1509 ( 
.A(n_1454),
.B(n_1470),
.C(n_1462),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1502),
.B(n_1461),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1501),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1476),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1478),
.B(n_1495),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1477),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1475),
.B(n_1461),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1505),
.B(n_1456),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1482),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1508),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1501),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1491),
.B(n_1461),
.Y(n_1520)
);

NAND3xp33_ASAP7_75t_L g1521 ( 
.A(n_1483),
.B(n_1463),
.C(n_1438),
.Y(n_1521)
);

INVx1_ASAP7_75t_SL g1522 ( 
.A(n_1508),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1491),
.B(n_1461),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1484),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1495),
.Y(n_1525)
);

INVxp67_ASAP7_75t_SL g1526 ( 
.A(n_1493),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1492),
.B(n_1463),
.Y(n_1527)
);

INVxp67_ASAP7_75t_L g1528 ( 
.A(n_1486),
.Y(n_1528)
);

INVx3_ASAP7_75t_L g1529 ( 
.A(n_1485),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1487),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1480),
.B(n_1469),
.Y(n_1531)
);

BUFx2_ASAP7_75t_L g1532 ( 
.A(n_1479),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1489),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1527),
.B(n_1504),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1525),
.B(n_1509),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1532),
.Y(n_1536)
);

AOI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1528),
.A2(n_1488),
.B(n_1486),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1528),
.B(n_1488),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_SL g1539 ( 
.A(n_1532),
.B(n_1498),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1525),
.B(n_1481),
.Y(n_1540)
);

AND2x6_ASAP7_75t_SL g1541 ( 
.A(n_1515),
.B(n_1414),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1532),
.B(n_1507),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1518),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1512),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1512),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1512),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1518),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1514),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1518),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1514),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1525),
.B(n_1491),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_L g1552 ( 
.A(n_1513),
.B(n_1442),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1526),
.B(n_1459),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1520),
.B(n_1523),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1526),
.A2(n_1469),
.B1(n_1503),
.B2(n_1494),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1520),
.B(n_1490),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1517),
.Y(n_1557)
);

NAND4xp25_ASAP7_75t_L g1558 ( 
.A(n_1513),
.B(n_1503),
.C(n_1470),
.D(n_1497),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1520),
.B(n_1499),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1520),
.B(n_1465),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1521),
.B(n_1469),
.Y(n_1561)
);

AOI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1521),
.A2(n_1469),
.B1(n_1494),
.B2(n_1426),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1521),
.B(n_1467),
.Y(n_1563)
);

INVx2_ASAP7_75t_SL g1564 ( 
.A(n_1518),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1511),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1511),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1540),
.B(n_1510),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1540),
.B(n_1510),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1550),
.Y(n_1569)
);

OAI32xp33_ASAP7_75t_L g1570 ( 
.A1(n_1542),
.A2(n_1515),
.A3(n_1531),
.B1(n_1529),
.B2(n_1522),
.Y(n_1570)
);

NAND2x1p5_ASAP7_75t_L g1571 ( 
.A(n_1564),
.B(n_1506),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_SL g1572 ( 
.A(n_1536),
.B(n_1442),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1560),
.B(n_1530),
.Y(n_1573)
);

O2A1O1Ixp33_ASAP7_75t_L g1574 ( 
.A1(n_1538),
.A2(n_1531),
.B(n_1515),
.C(n_1500),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1537),
.B(n_1524),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1537),
.B(n_1524),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1550),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1544),
.Y(n_1578)
);

INVx1_ASAP7_75t_SL g1579 ( 
.A(n_1538),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1560),
.B(n_1530),
.Y(n_1580)
);

O2A1O1Ixp33_ASAP7_75t_SL g1581 ( 
.A1(n_1542),
.A2(n_1531),
.B(n_1496),
.C(n_1474),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1544),
.Y(n_1582)
);

NAND3xp33_ASAP7_75t_L g1583 ( 
.A(n_1539),
.B(n_1500),
.C(n_1511),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1553),
.B(n_1533),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1545),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1553),
.B(n_1533),
.Y(n_1586)
);

INVx1_ASAP7_75t_SL g1587 ( 
.A(n_1541),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1545),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1561),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1546),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1534),
.B(n_1533),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1552),
.B(n_1424),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1564),
.Y(n_1593)
);

BUFx3_ASAP7_75t_L g1594 ( 
.A(n_1543),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1564),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1561),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1561),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1556),
.B(n_1516),
.Y(n_1598)
);

INVxp67_ASAP7_75t_L g1599 ( 
.A(n_1539),
.Y(n_1599)
);

AOI21xp33_ASAP7_75t_L g1600 ( 
.A1(n_1543),
.A2(n_1522),
.B(n_1511),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1556),
.B(n_1516),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1562),
.B(n_1424),
.Y(n_1602)
);

NOR3xp33_ASAP7_75t_L g1603 ( 
.A(n_1575),
.B(n_1558),
.C(n_1547),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1576),
.B(n_1534),
.Y(n_1604)
);

AND3x1_ASAP7_75t_L g1605 ( 
.A(n_1572),
.B(n_1562),
.C(n_1555),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1578),
.Y(n_1606)
);

NOR2xp67_ASAP7_75t_L g1607 ( 
.A(n_1583),
.B(n_1558),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1578),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1573),
.B(n_1559),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1579),
.A2(n_1561),
.B1(n_1555),
.B2(n_1547),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1573),
.B(n_1559),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1580),
.B(n_1551),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1589),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1587),
.Y(n_1614)
);

INVxp67_ASAP7_75t_SL g1615 ( 
.A(n_1572),
.Y(n_1615)
);

OAI221xp5_ASAP7_75t_L g1616 ( 
.A1(n_1599),
.A2(n_1563),
.B1(n_1549),
.B2(n_1547),
.C(n_1543),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1594),
.B(n_1554),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1579),
.B(n_1546),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1580),
.B(n_1551),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1569),
.B(n_1548),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1582),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1582),
.Y(n_1622)
);

BUFx2_ASAP7_75t_L g1623 ( 
.A(n_1593),
.Y(n_1623)
);

INVxp33_ASAP7_75t_L g1624 ( 
.A(n_1592),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1587),
.B(n_1554),
.Y(n_1625)
);

INVx4_ASAP7_75t_L g1626 ( 
.A(n_1594),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1595),
.Y(n_1627)
);

INVxp67_ASAP7_75t_L g1628 ( 
.A(n_1594),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1613),
.Y(n_1629)
);

AOI32xp33_ASAP7_75t_L g1630 ( 
.A1(n_1603),
.A2(n_1602),
.A3(n_1535),
.B1(n_1589),
.B2(n_1596),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1607),
.Y(n_1631)
);

OAI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1607),
.A2(n_1574),
.B(n_1583),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1613),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1613),
.Y(n_1634)
);

NAND2xp33_ASAP7_75t_R g1635 ( 
.A(n_1623),
.B(n_1535),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1606),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1604),
.B(n_1591),
.Y(n_1637)
);

AOI221xp5_ASAP7_75t_L g1638 ( 
.A1(n_1605),
.A2(n_1570),
.B1(n_1581),
.B2(n_1600),
.C(n_1597),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1615),
.B(n_1567),
.Y(n_1639)
);

AOI321xp33_ASAP7_75t_L g1640 ( 
.A1(n_1605),
.A2(n_1570),
.A3(n_1589),
.B1(n_1597),
.B2(n_1596),
.C(n_1600),
.Y(n_1640)
);

INVxp67_ASAP7_75t_SL g1641 ( 
.A(n_1628),
.Y(n_1641)
);

AOI31xp33_ASAP7_75t_L g1642 ( 
.A1(n_1614),
.A2(n_1569),
.A3(n_1577),
.B(n_1563),
.Y(n_1642)
);

OAI21xp33_ASAP7_75t_L g1643 ( 
.A1(n_1603),
.A2(n_1586),
.B(n_1584),
.Y(n_1643)
);

O2A1O1Ixp33_ASAP7_75t_L g1644 ( 
.A1(n_1614),
.A2(n_1577),
.B(n_1549),
.C(n_1597),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1628),
.B(n_1591),
.Y(n_1645)
);

OAI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1616),
.A2(n_1535),
.B(n_1549),
.Y(n_1646)
);

AOI221xp5_ASAP7_75t_L g1647 ( 
.A1(n_1610),
.A2(n_1596),
.B1(n_1522),
.B2(n_1507),
.C(n_1590),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1606),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1631),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1641),
.Y(n_1650)
);

AOI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1632),
.A2(n_1638),
.B1(n_1647),
.B2(n_1635),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1639),
.B(n_1625),
.Y(n_1652)
);

NAND2x1p5_ASAP7_75t_L g1653 ( 
.A(n_1629),
.B(n_1626),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1641),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1631),
.B(n_1625),
.Y(n_1655)
);

NAND2xp33_ASAP7_75t_L g1656 ( 
.A(n_1637),
.B(n_1604),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1642),
.B(n_1612),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1640),
.B(n_1626),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1645),
.Y(n_1659)
);

AOI211xp5_ASAP7_75t_L g1660 ( 
.A1(n_1658),
.A2(n_1646),
.B(n_1644),
.C(n_1643),
.Y(n_1660)
);

OAI211xp5_ASAP7_75t_L g1661 ( 
.A1(n_1658),
.A2(n_1630),
.B(n_1626),
.C(n_1627),
.Y(n_1661)
);

AOI221xp5_ASAP7_75t_L g1662 ( 
.A1(n_1651),
.A2(n_1616),
.B1(n_1633),
.B2(n_1634),
.C(n_1618),
.Y(n_1662)
);

O2A1O1Ixp33_ASAP7_75t_L g1663 ( 
.A1(n_1649),
.A2(n_1618),
.B(n_1648),
.C(n_1636),
.Y(n_1663)
);

NOR3xp33_ASAP7_75t_L g1664 ( 
.A(n_1655),
.B(n_1626),
.C(n_1623),
.Y(n_1664)
);

A2O1A1Ixp33_ASAP7_75t_L g1665 ( 
.A1(n_1657),
.A2(n_1535),
.B(n_1635),
.C(n_1624),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1656),
.A2(n_1627),
.B(n_1620),
.Y(n_1666)
);

OAI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1649),
.A2(n_1571),
.B1(n_1620),
.B2(n_1622),
.C(n_1608),
.Y(n_1667)
);

OAI221xp5_ASAP7_75t_L g1668 ( 
.A1(n_1659),
.A2(n_1571),
.B1(n_1608),
.B2(n_1621),
.C(n_1622),
.Y(n_1668)
);

AOI221xp5_ASAP7_75t_L g1669 ( 
.A1(n_1662),
.A2(n_1660),
.B1(n_1666),
.B2(n_1663),
.C(n_1665),
.Y(n_1669)
);

AOI211xp5_ASAP7_75t_SL g1670 ( 
.A1(n_1661),
.A2(n_1664),
.B(n_1650),
.C(n_1654),
.Y(n_1670)
);

AOI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1668),
.A2(n_1652),
.B(n_1667),
.Y(n_1671)
);

AO21x1_ASAP7_75t_L g1672 ( 
.A1(n_1660),
.A2(n_1653),
.B(n_1621),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1663),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1672),
.B(n_1653),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1673),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1670),
.B(n_1612),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1669),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1671),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1672),
.A2(n_1617),
.B(n_1619),
.Y(n_1679)
);

AND2x4_ASAP7_75t_L g1680 ( 
.A(n_1675),
.B(n_1617),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1677),
.Y(n_1681)
);

NAND2xp33_ASAP7_75t_R g1682 ( 
.A(n_1674),
.B(n_1617),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1676),
.Y(n_1683)
);

AOI31xp33_ASAP7_75t_L g1684 ( 
.A1(n_1678),
.A2(n_1619),
.A3(n_1617),
.B(n_1611),
.Y(n_1684)
);

OAI211xp5_ASAP7_75t_L g1685 ( 
.A1(n_1683),
.A2(n_1679),
.B(n_1681),
.C(n_1682),
.Y(n_1685)
);

NOR4xp75_ASAP7_75t_SL g1686 ( 
.A(n_1684),
.B(n_1541),
.C(n_1373),
.D(n_1376),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1680),
.B(n_1609),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1687),
.Y(n_1688)
);

OAI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1688),
.A2(n_1685),
.B1(n_1686),
.B2(n_1588),
.C(n_1585),
.Y(n_1689)
);

XNOR2x1_ASAP7_75t_L g1690 ( 
.A(n_1689),
.B(n_1680),
.Y(n_1690)
);

AND2x4_ASAP7_75t_L g1691 ( 
.A(n_1689),
.B(n_1609),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1691),
.B(n_1611),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1690),
.Y(n_1693)
);

AO22x2_ASAP7_75t_L g1694 ( 
.A1(n_1693),
.A2(n_1590),
.B1(n_1588),
.B2(n_1585),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1692),
.Y(n_1695)
);

XOR2xp5_ASAP7_75t_L g1696 ( 
.A(n_1695),
.B(n_1571),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1694),
.A2(n_1568),
.B1(n_1567),
.B2(n_1601),
.Y(n_1697)
);

INVx1_ASAP7_75t_SL g1698 ( 
.A(n_1696),
.Y(n_1698)
);

NOR4xp75_ASAP7_75t_L g1699 ( 
.A(n_1698),
.B(n_1697),
.C(n_1568),
.D(n_1598),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1699),
.A2(n_1566),
.B1(n_1565),
.B2(n_1519),
.Y(n_1700)
);

AOI221xp5_ASAP7_75t_L g1701 ( 
.A1(n_1700),
.A2(n_1566),
.B1(n_1565),
.B2(n_1557),
.C(n_1548),
.Y(n_1701)
);

AOI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1701),
.A2(n_1601),
.B1(n_1598),
.B2(n_1565),
.Y(n_1702)
);


endmodule