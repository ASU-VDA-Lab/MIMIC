module fake_jpeg_8731_n_328 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_17),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_1),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_41),
.B(n_47),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_42),
.B(n_25),
.Y(n_80)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_46),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_25),
.Y(n_79)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_30),
.Y(n_69)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_55),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_28),
.B1(n_30),
.B2(n_19),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_52),
.A2(n_26),
.B1(n_29),
.B2(n_34),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_32),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_53),
.B(n_64),
.Y(n_103)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_58),
.Y(n_96)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_62),
.B(n_65),
.Y(n_116)
);

AOI21xp33_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_31),
.B(n_27),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

NAND2xp33_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_31),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_67),
.A2(n_38),
.B1(n_33),
.B2(n_27),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_68),
.Y(n_97)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_18),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_73),
.Y(n_93)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_74),
.B(n_75),
.Y(n_101)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_76),
.B(n_78),
.Y(n_115)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_80),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_18),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_81),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_86),
.B1(n_23),
.B2(n_37),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_24),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_24),
.Y(n_117)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_85),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_43),
.A2(n_21),
.B1(n_23),
.B2(n_36),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_63),
.A2(n_37),
.B1(n_34),
.B2(n_32),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_88),
.A2(n_99),
.B1(n_102),
.B2(n_110),
.Y(n_130)
);

INVx6_ASAP7_75t_SL g89 ( 
.A(n_72),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_89),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_64),
.B1(n_52),
.B2(n_73),
.Y(n_91)
);

AO22x1_ASAP7_75t_L g124 ( 
.A1(n_91),
.A2(n_95),
.B1(n_112),
.B2(n_56),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_105),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_63),
.A2(n_29),
.B1(n_26),
.B2(n_38),
.Y(n_102)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_106),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_109),
.B(n_87),
.Y(n_126)
);

AOI22x1_ASAP7_75t_L g112 ( 
.A1(n_53),
.A2(n_35),
.B1(n_22),
.B2(n_3),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_121),
.Y(n_131)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_61),
.B(n_33),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_20),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_5),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_91),
.A2(n_82),
.B1(n_60),
.B2(n_66),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_123),
.A2(n_146),
.B1(n_152),
.B2(n_155),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_109),
.B1(n_116),
.B2(n_93),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_1),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_125),
.A2(n_136),
.B(n_144),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_126),
.B(n_147),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_108),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_111),
.Y(n_168)
);

INVx2_ASAP7_75t_R g132 ( 
.A(n_112),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_132),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_121),
.B(n_20),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_133),
.B(n_134),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_115),
.Y(n_134)
);

OR2x2_ASAP7_75t_SL g136 ( 
.A(n_103),
.B(n_2),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_142),
.Y(n_165)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_151),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_2),
.Y(n_144)
);

AND2x6_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_2),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_145),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_91),
.A2(n_60),
.B1(n_83),
.B2(n_7),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_3),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_3),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_148),
.B(n_155),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_149),
.B(n_150),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_122),
.B(n_7),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_120),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_153),
.Y(n_184)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_154),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_108),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_156),
.Y(n_190)
);

AO22x1_ASAP7_75t_SL g158 ( 
.A1(n_132),
.A2(n_124),
.B1(n_123),
.B2(n_146),
.Y(n_158)
);

AO22x1_ASAP7_75t_SL g210 ( 
.A1(n_158),
.A2(n_15),
.B1(n_16),
.B2(n_186),
.Y(n_210)
);

O2A1O1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_159),
.A2(n_162),
.B(n_164),
.C(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_160),
.B(n_169),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_118),
.B1(n_119),
.B2(n_117),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_113),
.B1(n_111),
.B2(n_107),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_96),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_166),
.B(n_167),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_92),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_140),
.C(n_129),
.Y(n_196)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_170),
.Y(n_212)
);

AO22x1_ASAP7_75t_L g173 ( 
.A1(n_125),
.A2(n_113),
.B1(n_105),
.B2(n_104),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_148),
.B(n_97),
.Y(n_175)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_178),
.Y(n_217)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

NOR2x1_ASAP7_75t_L g180 ( 
.A(n_125),
.B(n_65),
.Y(n_180)
);

AO21x1_ASAP7_75t_L g207 ( 
.A1(n_180),
.A2(n_182),
.B(n_183),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_145),
.A2(n_65),
.B1(n_58),
.B2(n_11),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_181),
.A2(n_179),
.B1(n_188),
.B2(n_183),
.Y(n_216)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_138),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_185),
.A2(n_187),
.B(n_16),
.Y(n_214)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_147),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_188),
.A2(n_153),
.B1(n_135),
.B2(n_154),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_144),
.B(n_10),
.Y(n_189)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_189),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_180),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_194),
.Y(n_221)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_158),
.A2(n_136),
.B1(n_144),
.B2(n_129),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_195),
.A2(n_202),
.B(n_205),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_201),
.C(n_209),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_197),
.A2(n_204),
.B1(n_210),
.B2(n_173),
.Y(n_230)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_206),
.Y(n_225)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_199),
.B(n_203),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_106),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_174),
.A2(n_135),
.B(n_106),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_174),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_163),
.A2(n_12),
.B(n_14),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_171),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_12),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_208),
.A2(n_215),
.B(n_205),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_100),
.C(n_15),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_161),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_219),
.Y(n_233)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_214),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_163),
.A2(n_186),
.B(n_169),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_216),
.A2(n_176),
.B1(n_173),
.B2(n_160),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_184),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_210),
.Y(n_237)
);

BUFx12_ASAP7_75t_L g223 ( 
.A(n_219),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_226),
.Y(n_248)
);

INVx13_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_224),
.Y(n_252)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_217),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_229),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_228),
.A2(n_232),
.B1(n_236),
.B2(n_243),
.Y(n_264)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_238),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_220),
.A2(n_176),
.B1(n_185),
.B2(n_187),
.Y(n_232)
);

BUFx12f_ASAP7_75t_SL g235 ( 
.A(n_210),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_235),
.A2(n_245),
.B(n_200),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_216),
.A2(n_184),
.B1(n_177),
.B2(n_178),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_237),
.A2(n_238),
.B1(n_191),
.B2(n_208),
.Y(n_246)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_201),
.B(n_157),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_234),
.Y(n_262)
);

BUFx24_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_196),
.B(n_157),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_209),
.C(n_215),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_192),
.A2(n_182),
.B1(n_190),
.B2(n_195),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_200),
.A2(n_212),
.B1(n_204),
.B2(n_208),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_244),
.A2(n_230),
.B1(n_222),
.B2(n_241),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_246),
.A2(n_257),
.B1(n_231),
.B2(n_244),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_225),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_247),
.A2(n_254),
.B(n_258),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_218),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_253),
.C(n_256),
.Y(n_279)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_218),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_224),
.A2(n_214),
.B1(n_203),
.B2(n_197),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_193),
.B(n_235),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_221),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_259),
.B(n_260),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_236),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_261),
.A2(n_265),
.B1(n_243),
.B2(n_232),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_234),
.Y(n_270)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_233),
.Y(n_263)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_263),
.Y(n_283)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_248),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_269),
.Y(n_284)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_268),
.Y(n_295)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_256),
.C(n_262),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_274),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_223),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_276),
.B(n_277),
.Y(n_286)
);

NOR3xp33_ASAP7_75t_SL g274 ( 
.A(n_258),
.B(n_245),
.C(n_228),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_265),
.Y(n_278)
);

INVxp67_ASAP7_75t_SL g287 ( 
.A(n_278),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_281),
.A2(n_282),
.B1(n_249),
.B2(n_276),
.Y(n_293)
);

INVx11_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

NOR2xp67_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_275),
.Y(n_285)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_285),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_291),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_253),
.C(n_250),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_292),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_264),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_281),
.A2(n_251),
.B1(n_249),
.B2(n_223),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_266),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_280),
.C(n_275),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_283),
.Y(n_299)
);

NOR2xp67_ASAP7_75t_SL g296 ( 
.A(n_282),
.B(n_283),
.Y(n_296)
);

NAND2xp33_ASAP7_75t_R g301 ( 
.A(n_296),
.B(n_266),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_289),
.C(n_288),
.Y(n_314)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_300),
.Y(n_313)
);

INVx11_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_268),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_302),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_284),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_304),
.B(n_305),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_295),
.A2(n_297),
.B1(n_287),
.B2(n_286),
.Y(n_305)
);

BUFx4f_ASAP7_75t_SL g307 ( 
.A(n_294),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_291),
.Y(n_308)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_308),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_305),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_312),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_307),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_314),
.A2(n_303),
.B(n_308),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_307),
.B1(n_298),
.B2(n_303),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_319),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_313),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_313),
.B(n_312),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_323),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_318),
.A2(n_311),
.B(n_315),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_322),
.Y(n_325)
);

AOI21x1_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_317),
.B(n_314),
.Y(n_326)
);

NOR3xp33_ASAP7_75t_SL g327 ( 
.A(n_326),
.B(n_309),
.C(n_311),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_316),
.C(n_324),
.Y(n_328)
);


endmodule