module real_aes_4041_n_406 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_401, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_399, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_400, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_398, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_405, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_402, n_87, n_171, n_78, n_1363, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_404, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_403, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_406);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_401;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_399;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_400;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_398;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_405;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_402;
input n_87;
input n_171;
input n_78;
input n_1363;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_404;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_403;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_406;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_592;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_786;
wire n_512;
wire n_795;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1325;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1317;
wire n_417;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_527;
wire n_1342;
wire n_1346;
wire n_552;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_591;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_550;
wire n_966;
wire n_994;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_617;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_807;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1194;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_943;
wire n_977;
wire n_905;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_816;
wire n_625;
wire n_953;
wire n_716;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_1207;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_727;
wire n_1083;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_1139;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_578;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_425;
wire n_879;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_1183;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_698;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_483;
wire n_1352;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1097;
wire n_703;
wire n_601;
wire n_463;
wire n_1236;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_0), .A2(n_384), .B1(n_574), .B2(n_756), .Y(n_755) );
AOI22x1_ASAP7_75t_L g803 ( .A1(n_1), .A2(n_254), .B1(n_563), .B2(n_685), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_2), .A2(n_168), .B1(n_506), .B2(n_507), .Y(n_505) );
AOI22xp33_ASAP7_75t_SL g1341 ( .A1(n_3), .A2(n_284), .B1(n_544), .B2(n_727), .Y(n_1341) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_4), .A2(n_259), .B1(n_499), .B2(n_500), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_5), .B(n_753), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_6), .A2(n_362), .B1(n_599), .B2(n_937), .Y(n_936) );
CKINVDCx5p33_ASAP7_75t_R g714 ( .A(n_7), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_8), .A2(n_361), .B1(n_529), .B2(n_956), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_9), .A2(n_210), .B1(n_556), .B2(n_558), .Y(n_1014) );
INVx1_ASAP7_75t_L g850 ( .A(n_10), .Y(n_850) );
AOI221xp5_ASAP7_75t_L g586 ( .A1(n_11), .A2(n_322), .B1(n_587), .B2(n_588), .C(n_589), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_12), .A2(n_331), .B1(n_615), .B2(n_646), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g933 ( .A1(n_13), .A2(n_113), .B1(n_675), .B2(n_934), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_14), .A2(n_242), .B1(n_685), .B2(n_724), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_15), .A2(n_227), .B1(n_499), .B2(n_500), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_16), .B(n_436), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_17), .A2(n_221), .B1(n_561), .B2(n_563), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_18), .A2(n_305), .B1(n_516), .B2(n_595), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g907 ( .A1(n_19), .A2(n_270), .B1(n_796), .B2(n_908), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_20), .A2(n_36), .B1(n_549), .B2(n_687), .Y(n_838) );
INVx1_ASAP7_75t_L g1311 ( .A(n_21), .Y(n_1311) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_22), .Y(n_436) );
INVx1_ASAP7_75t_L g751 ( .A(n_23), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g1128 ( .A1(n_24), .A2(n_298), .B1(n_1106), .B2(n_1108), .Y(n_1128) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_25), .A2(n_52), .B1(n_544), .B2(n_577), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g940 ( .A1(n_26), .A2(n_375), .B1(n_574), .B2(n_577), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_27), .A2(n_38), .B1(n_502), .B2(n_506), .Y(n_770) );
INVx1_ASAP7_75t_L g869 ( .A(n_28), .Y(n_869) );
AOI22xp5_ASAP7_75t_L g906 ( .A1(n_29), .A2(n_125), .B1(n_516), .B2(n_720), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_30), .A2(n_255), .B1(n_469), .B2(n_494), .Y(n_997) );
AOI22xp5_ASAP7_75t_L g1112 ( .A1(n_31), .A2(n_215), .B1(n_1106), .B2(n_1108), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_32), .A2(n_93), .B1(n_584), .B2(n_633), .Y(n_975) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_33), .B(n_617), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_34), .A2(n_321), .B1(n_805), .B2(n_958), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_35), .A2(n_207), .B1(n_582), .B2(n_584), .Y(n_581) );
AOI221xp5_ASAP7_75t_L g894 ( .A1(n_37), .A2(n_377), .B1(n_455), .B2(n_465), .C(n_895), .Y(n_894) );
AOI21xp33_ASAP7_75t_L g616 ( .A1(n_39), .A2(n_617), .B(n_618), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_40), .A2(n_386), .B1(n_1090), .B2(n_1104), .Y(n_1103) );
INVxp33_ASAP7_75t_SL g1091 ( .A(n_41), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_42), .A2(n_228), .B1(n_1097), .B2(n_1098), .Y(n_1196) );
AOI21xp5_ASAP7_75t_L g1345 ( .A1(n_43), .A2(n_958), .B(n_1346), .Y(n_1345) );
AO22x1_ASAP7_75t_L g1306 ( .A1(n_44), .A2(n_67), .B1(n_806), .B2(n_1307), .Y(n_1306) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_45), .A2(n_72), .B1(n_611), .B2(n_982), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g1197 ( .A1(n_46), .A2(n_61), .B1(n_1075), .B2(n_1095), .Y(n_1197) );
INVx1_ASAP7_75t_L g1347 ( .A(n_47), .Y(n_1347) );
AOI21xp5_ASAP7_75t_L g821 ( .A1(n_48), .A2(n_822), .B(n_824), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_49), .A2(n_217), .B1(n_595), .B2(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g485 ( .A(n_50), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_51), .A2(n_132), .B1(n_549), .B2(n_623), .Y(n_862) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_53), .A2(n_376), .B1(n_625), .B2(n_626), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_54), .A2(n_64), .B1(n_595), .B2(n_614), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_55), .A2(n_123), .B1(n_469), .B2(n_779), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_56), .A2(n_188), .B1(n_573), .B2(n_579), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_57), .A2(n_155), .B1(n_633), .B2(n_1035), .Y(n_1034) );
AOI22xp33_ASAP7_75t_L g1343 ( .A1(n_58), .A2(n_62), .B1(n_563), .B2(n_685), .Y(n_1343) );
AO22x1_ASAP7_75t_L g895 ( .A1(n_59), .A2(n_97), .B1(n_469), .B2(n_483), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_60), .A2(n_277), .B1(n_611), .B2(n_612), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g990 ( .A(n_61), .Y(n_990) );
INVx1_ASAP7_75t_L g527 ( .A(n_63), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_65), .A2(n_332), .B1(n_1040), .B2(n_1041), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_66), .B(n_656), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_68), .A2(n_216), .B1(n_558), .B2(n_682), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_69), .A2(n_191), .B1(n_516), .B2(n_677), .Y(n_676) );
OA22x2_ASAP7_75t_L g442 ( .A1(n_70), .A2(n_179), .B1(n_436), .B2(n_440), .Y(n_442) );
INVx1_ASAP7_75t_L g474 ( .A(n_70), .Y(n_474) );
AOI22xp33_ASAP7_75t_SL g1055 ( .A1(n_71), .A2(n_367), .B1(n_1056), .B2(n_1057), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_73), .A2(n_148), .B1(n_561), .B2(n_563), .Y(n_1012) );
AOI22xp5_ASAP7_75t_L g1129 ( .A1(n_74), .A2(n_318), .B1(n_1104), .B2(n_1114), .Y(n_1129) );
AOI21xp5_ASAP7_75t_L g1045 ( .A1(n_75), .A2(n_1046), .B(n_1047), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_76), .A2(n_334), .B1(n_582), .B2(n_584), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_77), .A2(n_176), .B1(n_561), .B2(n_563), .Y(n_914) );
AOI221x1_ASAP7_75t_L g642 ( .A1(n_78), .A2(n_291), .B1(n_629), .B2(n_633), .C(n_643), .Y(n_642) );
AOI22xp33_ASAP7_75t_SL g543 ( .A1(n_79), .A2(n_366), .B1(n_544), .B2(n_546), .Y(n_543) );
INVxp67_ASAP7_75t_L g835 ( .A(n_80), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_81), .A2(n_167), .B1(n_556), .B2(n_558), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_82), .A2(n_345), .B1(n_549), .B2(n_687), .Y(n_949) );
AOI22xp5_ASAP7_75t_L g1303 ( .A1(n_83), .A2(n_1304), .B1(n_1327), .B2(n_1328), .Y(n_1303) );
CKINVDCx5p33_ASAP7_75t_R g1327 ( .A(n_83), .Y(n_1327) );
AOI221xp5_ASAP7_75t_L g800 ( .A1(n_84), .A2(n_273), .B1(n_682), .B2(n_801), .C(n_802), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_85), .A2(n_314), .B1(n_704), .B2(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g1133 ( .A(n_86), .Y(n_1133) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_87), .A2(n_390), .B1(n_529), .B2(n_679), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_88), .A2(n_400), .B1(n_576), .B2(n_577), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_89), .A2(n_193), .B1(n_561), .B2(n_563), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_90), .A2(n_372), .B1(n_735), .B2(n_737), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g974 ( .A1(n_91), .A2(n_163), .B1(n_551), .B2(n_577), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_92), .A2(n_364), .B1(n_465), .B2(n_469), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_94), .B(n_199), .Y(n_415) );
INVx1_ASAP7_75t_L g439 ( .A(n_94), .Y(n_439) );
OAI21xp33_ASAP7_75t_L g475 ( .A1(n_94), .A2(n_179), .B(n_463), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g1326 ( .A1(n_95), .A2(n_344), .B1(n_682), .B2(n_801), .Y(n_1326) );
AOI221x1_ASAP7_75t_L g901 ( .A1(n_96), .A2(n_378), .B1(n_708), .B2(n_902), .C(n_904), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_98), .A2(n_126), .B1(n_573), .B2(n_579), .Y(n_941) );
INVx1_ASAP7_75t_L g811 ( .A(n_99), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_100), .A2(n_235), .B1(n_431), .B2(n_502), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_101), .A2(n_260), .B1(n_431), .B2(n_507), .Y(n_768) );
NOR3xp33_ASAP7_75t_L g639 ( .A(n_102), .B(n_640), .C(n_644), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_102), .A2(n_644), .B1(n_650), .B2(n_1363), .Y(n_664) );
OAI21xp5_ASAP7_75t_L g665 ( .A1(n_102), .A2(n_640), .B(n_658), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_103), .A2(n_185), .B1(n_499), .B2(n_500), .Y(n_771) );
AOI21xp33_ASAP7_75t_L g775 ( .A1(n_104), .A2(n_494), .B(n_776), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_105), .A2(n_109), .B1(n_546), .B2(n_576), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g1324 ( .A1(n_106), .A2(n_226), .B1(n_735), .B2(n_1325), .Y(n_1324) );
INVxp33_ASAP7_75t_L g1080 ( .A(n_107), .Y(n_1080) );
INVx1_ASAP7_75t_L g1079 ( .A(n_108), .Y(n_1079) );
AND2x4_ASAP7_75t_L g1087 ( .A(n_108), .B(n_301), .Y(n_1087) );
HB1xp67_ASAP7_75t_L g1360 ( .A(n_108), .Y(n_1360) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_110), .A2(n_230), .B1(n_576), .B2(n_660), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_111), .A2(n_117), .B1(n_495), .B2(n_503), .Y(n_769) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_112), .A2(n_672), .B(n_674), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_114), .A2(n_261), .B1(n_587), .B2(n_599), .Y(n_820) );
AOI21xp33_ASAP7_75t_L g482 ( .A1(n_115), .A2(n_483), .B(n_484), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g1018 ( .A1(n_116), .A2(n_652), .B(n_1019), .Y(n_1018) );
XNOR2x2_ASAP7_75t_L g858 ( .A(n_118), .B(n_859), .Y(n_858) );
AOI211xp5_ASAP7_75t_L g789 ( .A1(n_119), .A2(n_790), .B(n_792), .C(n_798), .Y(n_789) );
AOI22xp5_ASAP7_75t_L g793 ( .A1(n_120), .A2(n_214), .B1(n_529), .B2(n_794), .Y(n_793) );
AOI22xp5_ASAP7_75t_L g996 ( .A1(n_121), .A2(n_182), .B1(n_465), .B2(n_982), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_122), .A2(n_256), .B1(n_544), .B2(n_727), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g918 ( .A1(n_124), .A2(n_243), .B1(n_549), .B2(n_799), .Y(n_918) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_127), .A2(n_280), .B1(n_556), .B2(n_558), .Y(n_814) );
INVx1_ASAP7_75t_L g989 ( .A(n_128), .Y(n_989) );
INVx1_ASAP7_75t_L g525 ( .A(n_129), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_130), .A2(n_251), .B1(n_556), .B2(n_558), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_131), .A2(n_153), .B1(n_576), .B2(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g1077 ( .A(n_133), .Y(n_1077) );
AND2x4_ASAP7_75t_L g1082 ( .A(n_133), .B(n_411), .Y(n_1082) );
INVx1_ASAP7_75t_SL g1107 ( .A(n_133), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_134), .A2(n_323), .B1(n_735), .B2(n_799), .Y(n_1340) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_135), .A2(n_395), .B1(n_584), .B2(n_633), .Y(n_1005) );
AOI22xp5_ASAP7_75t_L g1117 ( .A1(n_136), .A2(n_263), .B1(n_1104), .B2(n_1114), .Y(n_1117) );
CKINVDCx16_ASAP7_75t_R g760 ( .A(n_137), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_138), .A2(n_295), .B1(n_595), .B2(n_711), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_139), .A2(n_166), .B1(n_1053), .B2(n_1054), .Y(n_1052) );
XNOR2x1_ASAP7_75t_L g427 ( .A(n_140), .B(n_428), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_141), .A2(n_328), .B1(n_455), .B2(n_465), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_142), .B(n_587), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_143), .A2(n_326), .B1(n_549), .B2(n_551), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g1342 ( .A1(n_144), .A2(n_380), .B1(n_632), .B2(n_682), .Y(n_1342) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_145), .A2(n_257), .B1(n_626), .B2(n_662), .Y(n_994) );
AOI22xp5_ASAP7_75t_L g1025 ( .A1(n_146), .A2(n_308), .B1(n_529), .B2(n_902), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_147), .A2(n_306), .B1(n_1097), .B2(n_1098), .Y(n_1096) );
AO22x1_ASAP7_75t_L g674 ( .A1(n_149), .A2(n_240), .B1(n_612), .B2(n_675), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_150), .A2(n_190), .B1(n_502), .B2(n_503), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_151), .A2(n_184), .B1(n_576), .B2(n_577), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_152), .A2(n_342), .B1(n_516), .B2(n_704), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_154), .B(n_479), .Y(n_478) );
NAND2xp33_ASAP7_75t_L g641 ( .A(n_156), .B(n_623), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_157), .A2(n_392), .B1(n_529), .B2(n_587), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_158), .A2(n_262), .B1(n_576), .B2(n_577), .Y(n_913) );
AOI22xp5_ASAP7_75t_L g1013 ( .A1(n_159), .A2(n_389), .B1(n_544), .B2(n_577), .Y(n_1013) );
AOI22xp5_ASAP7_75t_L g995 ( .A1(n_160), .A2(n_194), .B1(n_579), .B2(n_580), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_161), .A2(n_200), .B1(n_573), .B2(n_630), .Y(n_979) );
INVxp67_ASAP7_75t_SL g945 ( .A(n_162), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_164), .B(n_1350), .Y(n_1349) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_165), .A2(n_399), .B1(n_544), .B2(n_577), .Y(n_950) );
INVx1_ASAP7_75t_L g777 ( .A(n_169), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_170), .A2(n_401), .B1(n_1075), .B2(n_1095), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_171), .A2(n_292), .B1(n_576), .B2(n_577), .Y(n_575) );
INVx1_ASAP7_75t_L g825 ( .A(n_172), .Y(n_825) );
AO22x1_ASAP7_75t_L g807 ( .A1(n_173), .A2(n_253), .B1(n_544), .B2(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g1051 ( .A(n_174), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_175), .A2(n_374), .B1(n_1037), .B2(n_1038), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_177), .A2(n_192), .B1(n_556), .B2(n_801), .Y(n_951) );
INVx1_ASAP7_75t_L g454 ( .A(n_178), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_178), .B(n_237), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_178), .B(n_472), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_179), .B(n_316), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g668 ( .A(n_180), .Y(n_668) );
AND2x2_ASAP7_75t_L g643 ( .A(n_181), .B(n_627), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g1116 ( .A1(n_183), .A2(n_187), .B1(n_1106), .B2(n_1108), .Y(n_1116) );
AOI21xp33_ASAP7_75t_L g867 ( .A1(n_186), .A2(n_479), .B(n_868), .Y(n_867) );
XNOR2x1_ASAP7_75t_L g991 ( .A(n_187), .B(n_992), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_189), .A2(n_320), .B1(n_556), .B2(n_558), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_195), .A2(n_393), .B1(n_727), .B2(n_1043), .Y(n_1042) );
AO22x1_ASAP7_75t_L g798 ( .A1(n_196), .A2(n_340), .B1(n_549), .B2(n_799), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_197), .B(n_711), .Y(n_828) );
AOI22xp5_ASAP7_75t_L g871 ( .A1(n_198), .A2(n_229), .B1(n_584), .B2(n_633), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_199), .B(n_447), .Y(n_446) );
AOI22xp33_ASAP7_75t_SL g631 ( .A1(n_201), .A2(n_368), .B1(n_632), .B2(n_633), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_202), .A2(n_373), .B1(n_629), .B2(n_630), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_203), .A2(n_233), .B1(n_599), .B2(n_648), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_204), .B(n_1024), .Y(n_1023) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_205), .A2(n_336), .B1(n_546), .B2(n_623), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_206), .A2(n_231), .B1(n_561), .B2(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g864 ( .A(n_208), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_209), .A2(n_300), .B1(n_623), .B2(n_629), .Y(n_999) );
AOI21xp33_ASAP7_75t_SL g987 ( .A1(n_211), .A2(n_516), .B(n_988), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_212), .A2(n_351), .B1(n_579), .B2(n_580), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_213), .A2(n_287), .B1(n_611), .B2(n_612), .Y(n_938) );
INVx1_ASAP7_75t_L g780 ( .A(n_215), .Y(n_780) );
OA22x2_ASAP7_75t_L g884 ( .A1(n_218), .A2(n_885), .B1(n_896), .B2(n_897), .Y(n_884) );
INVx1_ASAP7_75t_L g897 ( .A(n_218), .Y(n_897) );
AOI221xp5_ASAP7_75t_L g804 ( .A1(n_219), .A2(n_232), .B1(n_805), .B2(n_806), .C(n_807), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g1316 ( .A1(n_220), .A2(n_224), .B1(n_711), .B2(n_982), .Y(n_1316) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_222), .A2(n_293), .B1(n_1086), .B2(n_1090), .Y(n_1134) );
AOI22xp33_ASAP7_75t_SL g1113 ( .A1(n_223), .A2(n_303), .B1(n_1104), .B2(n_1114), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_225), .A2(n_402), .B1(n_611), .B2(n_612), .Y(n_610) );
INVx1_ASAP7_75t_L g930 ( .A(n_234), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_236), .A2(n_286), .B1(n_876), .B2(n_986), .Y(n_985) );
INVx1_ASAP7_75t_L g437 ( .A(n_237), .Y(n_437) );
OAI22x1_ASAP7_75t_L g1009 ( .A1(n_238), .A2(n_1010), .B1(n_1015), .B2(n_1026), .Y(n_1009) );
NAND5xp2_ASAP7_75t_SL g1010 ( .A(n_238), .B(n_1011), .C(n_1012), .D(n_1013), .E(n_1014), .Y(n_1010) );
AOI22xp5_ASAP7_75t_L g1105 ( .A1(n_238), .A2(n_244), .B1(n_1106), .B2(n_1108), .Y(n_1105) );
INVx1_ASAP7_75t_L g706 ( .A(n_239), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g960 ( .A1(n_241), .A2(n_672), .B(n_961), .Y(n_960) );
AOI22xp5_ASAP7_75t_L g887 ( .A1(n_245), .A2(n_403), .B1(n_495), .B2(n_503), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_246), .A2(n_355), .B1(n_614), .B2(n_615), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_247), .A2(n_387), .B1(n_796), .B2(n_797), .Y(n_795) );
INVx1_ASAP7_75t_L g718 ( .A(n_248), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_249), .A2(n_290), .B1(n_549), .B2(n_687), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_250), .A2(n_365), .B1(n_630), .B2(n_725), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g1348 ( .A1(n_252), .A2(n_311), .B1(n_677), .B2(n_796), .Y(n_1348) );
AOI22xp5_ASAP7_75t_L g890 ( .A1(n_258), .A2(n_354), .B1(n_506), .B2(n_507), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_264), .A2(n_304), .B1(n_538), .B2(n_540), .Y(n_537) );
XNOR2x1_ASAP7_75t_L g606 ( .A(n_265), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g1309 ( .A(n_266), .Y(n_1309) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_267), .A2(n_278), .B1(n_431), .B2(n_455), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_268), .A2(n_352), .B1(n_654), .B2(n_656), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_269), .A2(n_394), .B1(n_682), .B2(n_730), .Y(n_729) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_271), .A2(n_383), .B1(n_632), .B2(n_660), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_272), .A2(n_388), .B1(n_611), .B2(n_876), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_274), .A2(n_357), .B1(n_598), .B2(n_599), .Y(n_597) );
AO22x2_ASAP7_75t_L g1031 ( .A1(n_275), .A2(n_1032), .B1(n_1059), .B2(n_1060), .Y(n_1031) );
INVx1_ASAP7_75t_L g1060 ( .A(n_275), .Y(n_1060) );
AOI22xp5_ASAP7_75t_L g1321 ( .A1(n_276), .A2(n_359), .B1(n_577), .B2(n_1322), .Y(n_1321) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_279), .A2(n_302), .B1(n_573), .B2(n_574), .Y(n_572) );
INVx1_ASAP7_75t_L g1004 ( .A(n_281), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_282), .B(n_753), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_283), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g532 ( .A(n_285), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g1319 ( .A1(n_288), .A2(n_324), .B1(n_1043), .B2(n_1320), .Y(n_1319) );
AOI221xp5_ASAP7_75t_SL g891 ( .A1(n_289), .A2(n_347), .B1(n_479), .B2(n_494), .C(n_892), .Y(n_891) );
AOI22xp5_ASAP7_75t_L g943 ( .A1(n_294), .A2(n_397), .B1(n_576), .B2(n_841), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_296), .A2(n_341), .B1(n_549), .B2(n_687), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_297), .A2(n_313), .B1(n_549), .B2(n_687), .Y(n_815) );
INVx1_ASAP7_75t_L g740 ( .A(n_298), .Y(n_740) );
CKINVDCx5p33_ASAP7_75t_R g701 ( .A(n_299), .Y(n_701) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_301), .Y(n_416) );
AND2x4_ASAP7_75t_L g1078 ( .A(n_301), .B(n_1079), .Y(n_1078) );
AOI22xp5_ASAP7_75t_L g845 ( .A1(n_307), .A2(n_333), .B1(n_598), .B2(n_846), .Y(n_845) );
CKINVDCx5p33_ASAP7_75t_R g700 ( .A(n_309), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g1351 ( .A1(n_310), .A2(n_396), .B1(n_720), .B2(n_794), .Y(n_1351) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_312), .A2(n_358), .B1(n_579), .B2(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g590 ( .A(n_315), .Y(n_590) );
INVx1_ASAP7_75t_L g452 ( .A(n_316), .Y(n_452) );
INVxp67_ASAP7_75t_L g462 ( .A(n_316), .Y(n_462) );
AOI21xp33_ASAP7_75t_L g848 ( .A1(n_317), .A2(n_516), .B(n_849), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_319), .B(n_794), .Y(n_935) );
INVx2_ASAP7_75t_L g411 ( .A(n_325), .Y(n_411) );
INVx1_ASAP7_75t_L g518 ( .A(n_327), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_329), .A2(n_382), .B1(n_563), .B2(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g619 ( .A(n_330), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_335), .A2(n_353), .B1(n_561), .B2(n_660), .Y(n_816) );
INVx1_ASAP7_75t_L g1083 ( .A(n_337), .Y(n_1083) );
INVx1_ASAP7_75t_L g905 ( .A(n_338), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_339), .A2(n_379), .B1(n_582), .B2(n_584), .Y(n_758) );
AOI221xp5_ASAP7_75t_L g1000 ( .A1(n_343), .A2(n_370), .B1(n_986), .B2(n_1001), .C(n_1003), .Y(n_1000) );
INVx2_ASAP7_75t_R g510 ( .A(n_346), .Y(n_510) );
CKINVDCx5p33_ASAP7_75t_R g893 ( .A(n_348), .Y(n_893) );
CKINVDCx14_ASAP7_75t_R g787 ( .A(n_349), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_350), .B(n_708), .Y(n_844) );
INVx1_ASAP7_75t_L g964 ( .A(n_356), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_360), .A2(n_398), .B1(n_494), .B2(n_495), .Y(n_493) );
INVx1_ASAP7_75t_L g1020 ( .A(n_363), .Y(n_1020) );
INVx1_ASAP7_75t_L g514 ( .A(n_369), .Y(n_514) );
INVx1_ASAP7_75t_L g1088 ( .A(n_371), .Y(n_1088) );
AOI22xp5_ASAP7_75t_L g1334 ( .A1(n_371), .A2(n_1335), .B1(n_1355), .B2(n_1357), .Y(n_1334) );
OAI21xp5_ASAP7_75t_L g1337 ( .A1(n_371), .A2(n_1338), .B(n_1352), .Y(n_1337) );
INVx1_ASAP7_75t_L g1049 ( .A(n_381), .Y(n_1049) );
INVx1_ASAP7_75t_L g1314 ( .A(n_385), .Y(n_1314) );
OAI21x1_ASAP7_75t_L g898 ( .A1(n_391), .A2(n_899), .B(n_919), .Y(n_898) );
INVx1_ASAP7_75t_L g922 ( .A(n_391), .Y(n_922) );
XNOR2x1_ASAP7_75t_L g569 ( .A(n_404), .B(n_570), .Y(n_569) );
AOI21xp33_ASAP7_75t_L g747 ( .A1(n_405), .A2(n_748), .B(n_750), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_417), .B(n_1066), .Y(n_406) );
INVx2_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
NAND3xp33_ASAP7_75t_L g408 ( .A(n_409), .B(n_412), .C(n_416), .Y(n_408) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_409), .B(n_1333), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_409), .B(n_1356), .Y(n_1355) );
AOI21xp5_ASAP7_75t_L g1361 ( .A1(n_409), .A2(n_416), .B(n_1107), .Y(n_1361) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AO21x1_ASAP7_75t_L g1358 ( .A1(n_410), .A2(n_1359), .B(n_1361), .Y(n_1358) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_411), .B(n_1077), .Y(n_1076) );
AND3x4_ASAP7_75t_L g1106 ( .A(n_411), .B(n_1078), .C(n_1107), .Y(n_1106) );
NOR2xp33_ASAP7_75t_L g1356 ( .A(n_412), .B(n_1333), .Y(n_1356) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AO21x2_ASAP7_75t_L g488 ( .A1(n_413), .A2(n_489), .B(n_490), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVx1_ASAP7_75t_L g1333 ( .A(n_416), .Y(n_1333) );
XNOR2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_829), .Y(n_417) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B1(n_691), .B2(n_692), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AO22x2_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_422), .B1(n_602), .B2(n_603), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OAI22x1_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_424), .B1(n_567), .B2(n_601), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AO22x2_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_508), .B1(n_509), .B2(n_566), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g566 ( .A(n_427), .Y(n_566) );
NOR2x1_ASAP7_75t_L g428 ( .A(n_429), .B(n_492), .Y(n_428) );
NAND4xp25_ASAP7_75t_L g429 ( .A(n_430), .B(n_464), .C(n_478), .D(n_482), .Y(n_429) );
AND2x4_ASAP7_75t_L g431 ( .A(n_432), .B(n_443), .Y(n_431) );
AND2x4_ASAP7_75t_L g499 ( .A(n_432), .B(n_467), .Y(n_499) );
AND2x4_ASAP7_75t_L g500 ( .A(n_432), .B(n_476), .Y(n_500) );
AND2x4_ASAP7_75t_L g502 ( .A(n_432), .B(n_496), .Y(n_502) );
AND2x4_ASAP7_75t_L g550 ( .A(n_432), .B(n_504), .Y(n_550) );
AND2x4_ASAP7_75t_L g557 ( .A(n_432), .B(n_467), .Y(n_557) );
AND2x2_ASAP7_75t_L g559 ( .A(n_432), .B(n_476), .Y(n_559) );
AND2x4_ASAP7_75t_L g562 ( .A(n_432), .B(n_496), .Y(n_562) );
AND2x4_ASAP7_75t_L g432 ( .A(n_433), .B(n_441), .Y(n_432) );
AND2x2_ASAP7_75t_L g481 ( .A(n_433), .B(n_442), .Y(n_481) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g466 ( .A(n_434), .B(n_442), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_438), .Y(n_434) );
NAND2xp33_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx2_ASAP7_75t_L g440 ( .A(n_436), .Y(n_440) );
INVx3_ASAP7_75t_L g447 ( .A(n_436), .Y(n_447) );
NAND2xp33_ASAP7_75t_L g453 ( .A(n_436), .B(n_454), .Y(n_453) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_436), .Y(n_458) );
INVx1_ASAP7_75t_L g463 ( .A(n_436), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_437), .B(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_439), .A2(n_462), .B(n_463), .Y(n_461) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g460 ( .A(n_442), .B(n_461), .Y(n_460) );
AND2x4_ASAP7_75t_L g547 ( .A(n_443), .B(n_466), .Y(n_547) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g504 ( .A(n_444), .Y(n_504) );
OR2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_449), .Y(n_444) );
AND2x2_ASAP7_75t_L g456 ( .A(n_445), .B(n_457), .Y(n_456) );
AND2x4_ASAP7_75t_L g467 ( .A(n_445), .B(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g477 ( .A(n_445), .Y(n_477) );
AND2x4_ASAP7_75t_L g496 ( .A(n_445), .B(n_497), .Y(n_496) );
AND2x4_ASAP7_75t_L g445 ( .A(n_446), .B(n_448), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_447), .B(n_452), .Y(n_451) );
INVxp67_ASAP7_75t_L g472 ( .A(n_447), .Y(n_472) );
NAND3xp33_ASAP7_75t_L g490 ( .A(n_448), .B(n_471), .C(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g497 ( .A(n_449), .Y(n_497) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g468 ( .A(n_450), .Y(n_468) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_453), .Y(n_450) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_460), .Y(n_455) );
AND2x4_ASAP7_75t_L g539 ( .A(n_456), .B(n_460), .Y(n_539) );
AND2x4_ASAP7_75t_L g827 ( .A(n_456), .B(n_460), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
INVx1_ASAP7_75t_L g489 ( .A(n_458), .Y(n_489) );
AND2x4_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
AND2x2_ASAP7_75t_L g483 ( .A(n_466), .B(n_476), .Y(n_483) );
AND2x4_ASAP7_75t_L g495 ( .A(n_466), .B(n_496), .Y(n_495) );
AND2x4_ASAP7_75t_L g503 ( .A(n_466), .B(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g523 ( .A(n_466), .B(n_467), .Y(n_523) );
AND2x2_ASAP7_75t_L g536 ( .A(n_466), .B(n_476), .Y(n_536) );
AND2x2_ASAP7_75t_L g545 ( .A(n_466), .B(n_496), .Y(n_545) );
AND2x2_ASAP7_75t_L g627 ( .A(n_466), .B(n_496), .Y(n_627) );
AND2x4_ASAP7_75t_L g494 ( .A(n_467), .B(n_481), .Y(n_494) );
AND2x4_ASAP7_75t_L g517 ( .A(n_467), .B(n_481), .Y(n_517) );
AND2x4_ASAP7_75t_L g476 ( .A(n_468), .B(n_477), .Y(n_476) );
AND2x4_ASAP7_75t_L g469 ( .A(n_470), .B(n_476), .Y(n_469) );
AND2x4_ASAP7_75t_L g506 ( .A(n_470), .B(n_496), .Y(n_506) );
AND2x4_ASAP7_75t_L g507 ( .A(n_470), .B(n_504), .Y(n_507) );
AND2x4_ASAP7_75t_L g530 ( .A(n_470), .B(n_476), .Y(n_530) );
AND2x4_ASAP7_75t_L g553 ( .A(n_470), .B(n_504), .Y(n_553) );
AND2x4_ASAP7_75t_L g565 ( .A(n_470), .B(n_496), .Y(n_565) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_475), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
AND2x4_ASAP7_75t_L g480 ( .A(n_476), .B(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g779 ( .A(n_476), .B(n_481), .Y(n_779) );
BUFx3_ASAP7_75t_L g956 ( .A(n_479), .Y(n_956) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g526 ( .A(n_480), .Y(n_526) );
BUFx8_ASAP7_75t_SL g587 ( .A(n_480), .Y(n_587) );
BUFx3_ASAP7_75t_L g648 ( .A(n_480), .Y(n_648) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_480), .Y(n_717) );
INVx2_ASAP7_75t_L g903 ( .A(n_480), .Y(n_903) );
INVx2_ASAP7_75t_L g1002 ( .A(n_483), .Y(n_1002) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
INVx1_ASAP7_75t_L g540 ( .A(n_486), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_486), .B(n_751), .Y(n_750) );
INVx4_ASAP7_75t_L g797 ( .A(n_486), .Y(n_797) );
NOR2xp33_ASAP7_75t_L g904 ( .A(n_486), .B(n_905), .Y(n_904) );
NOR2xp33_ASAP7_75t_L g1019 ( .A(n_486), .B(n_1020), .Y(n_1019) );
INVx4_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx3_ASAP7_75t_L g712 ( .A(n_487), .Y(n_712) );
INVx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_488), .Y(n_593) );
NAND4xp25_ASAP7_75t_L g492 ( .A(n_493), .B(n_498), .C(n_501), .D(n_505), .Y(n_492) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
XNOR2x1_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_541), .Y(n_511) );
NOR3xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_524), .C(n_531), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B1(n_518), .B2(n_519), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_515), .A2(n_700), .B1(n_701), .B2(n_702), .Y(n_699) );
INVx4_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx3_ASAP7_75t_L g614 ( .A(n_517), .Y(n_614) );
BUFx3_ASAP7_75t_L g652 ( .A(n_517), .Y(n_652) );
INVx1_ASAP7_75t_L g749 ( .A(n_517), .Y(n_749) );
INVxp67_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g598 ( .A(n_521), .Y(n_598) );
INVx1_ASAP7_75t_L g677 ( .A(n_521), .Y(n_677) );
INVx2_ASAP7_75t_L g1307 ( .A(n_521), .Y(n_1307) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g646 ( .A(n_522), .Y(n_646) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_523), .Y(n_611) );
BUFx3_ASAP7_75t_L g704 ( .A(n_523), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_526), .B1(n_527), .B2(n_528), .Y(n_524) );
INVx2_ASAP7_75t_L g679 ( .A(n_526), .Y(n_679) );
INVx3_ASAP7_75t_L g794 ( .A(n_526), .Y(n_794) );
INVx4_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx3_ASAP7_75t_L g1054 ( .A(n_529), .Y(n_1054) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx3_ASAP7_75t_L g600 ( .A(n_530), .Y(n_600) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_530), .Y(n_615) );
OAI21xp33_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B(n_537), .Y(n_531) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g588 ( .A(n_535), .Y(n_588) );
INVx3_ASAP7_75t_SL g753 ( .A(n_535), .Y(n_753) );
INVx2_ASAP7_75t_L g791 ( .A(n_535), .Y(n_791) );
INVx2_ASAP7_75t_L g934 ( .A(n_535), .Y(n_934) );
INVx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx3_ASAP7_75t_L g617 ( .A(n_536), .Y(n_617) );
INVx2_ASAP7_75t_L g655 ( .A(n_536), .Y(n_655) );
BUFx4f_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx5_ASAP7_75t_L g596 ( .A(n_539), .Y(n_596) );
BUFx2_ASAP7_75t_L g612 ( .A(n_539), .Y(n_612) );
BUFx2_ASAP7_75t_L g963 ( .A(n_539), .Y(n_963) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_554), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_548), .Y(n_542) );
BUFx8_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_545), .Y(n_576) );
BUFx3_ASAP7_75t_L g727 ( .A(n_546), .Y(n_727) );
BUFx12f_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_547), .Y(n_577) );
BUFx6f_ASAP7_75t_L g662 ( .A(n_547), .Y(n_662) );
BUFx6f_ASAP7_75t_L g756 ( .A(n_547), .Y(n_756) );
BUFx3_ASAP7_75t_L g808 ( .A(n_547), .Y(n_808) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
BUFx6f_ASAP7_75t_L g573 ( .A(n_550), .Y(n_573) );
BUFx6f_ASAP7_75t_L g629 ( .A(n_550), .Y(n_629) );
BUFx6f_ASAP7_75t_L g736 ( .A(n_550), .Y(n_736) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx3_ASAP7_75t_L g574 ( .A(n_552), .Y(n_574) );
INVx5_ASAP7_75t_L g623 ( .A(n_552), .Y(n_623) );
INVx2_ASAP7_75t_L g739 ( .A(n_552), .Y(n_739) );
INVx1_ASAP7_75t_L g799 ( .A(n_552), .Y(n_799) );
INVx6_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx12f_ASAP7_75t_L g687 ( .A(n_553), .Y(n_687) );
NAND2xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_560), .Y(n_554) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx3_ASAP7_75t_L g583 ( .A(n_557), .Y(n_583) );
BUFx12f_ASAP7_75t_L g633 ( .A(n_557), .Y(n_633) );
BUFx3_ASAP7_75t_L g1035 ( .A(n_558), .Y(n_1035) );
BUFx5_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_559), .Y(n_584) );
BUFx3_ASAP7_75t_L g632 ( .A(n_559), .Y(n_632) );
INVx1_ASAP7_75t_L g733 ( .A(n_559), .Y(n_733) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx12f_ASAP7_75t_L g579 ( .A(n_562), .Y(n_579) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_562), .Y(n_630) );
INVx4_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_SL g580 ( .A(n_564), .Y(n_580) );
INVx2_ASAP7_75t_L g625 ( .A(n_564), .Y(n_625) );
INVx4_ASAP7_75t_L g660 ( .A(n_564), .Y(n_660) );
INVx4_ASAP7_75t_L g725 ( .A(n_564), .Y(n_725) );
INVx2_ASAP7_75t_L g841 ( .A(n_564), .Y(n_841) );
INVx1_ASAP7_75t_L g978 ( .A(n_564), .Y(n_978) );
INVx8_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g601 ( .A(n_567), .Y(n_601) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NOR2x1_ASAP7_75t_L g570 ( .A(n_571), .B(n_585), .Y(n_570) );
NAND4xp25_ASAP7_75t_L g571 ( .A(n_572), .B(n_575), .C(n_578), .D(n_581), .Y(n_571) );
BUFx3_ASAP7_75t_L g1037 ( .A(n_573), .Y(n_1037) );
BUFx3_ASAP7_75t_L g1043 ( .A(n_576), .Y(n_1043) );
BUFx12f_ASAP7_75t_L g685 ( .A(n_579), .Y(n_685) );
BUFx6f_ASAP7_75t_L g1325 ( .A(n_579), .Y(n_1325) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g683 ( .A(n_583), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g585 ( .A(n_586), .B(n_594), .C(n_597), .Y(n_585) );
HB1xp67_ASAP7_75t_L g1053 ( .A(n_587), .Y(n_1053) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_591), .B(n_869), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g1346 ( .A(n_591), .B(n_1347), .Y(n_1346) );
INVx3_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
BUFx6f_ASAP7_75t_L g620 ( .A(n_593), .Y(n_620) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_593), .Y(n_657) );
INVx1_ASAP7_75t_L g675 ( .A(n_593), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g892 ( .A(n_593), .B(n_893), .Y(n_892) );
INVx4_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx3_ASAP7_75t_L g796 ( .A(n_596), .Y(n_796) );
INVx2_ASAP7_75t_L g846 ( .A(n_596), .Y(n_846) );
INVx2_ASAP7_75t_L g982 ( .A(n_596), .Y(n_982) );
INVx2_ASAP7_75t_L g1022 ( .A(n_596), .Y(n_1022) );
INVx3_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g876 ( .A(n_600), .Y(n_876) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AO22x1_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_634), .B1(n_635), .B2(n_689), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
BUFx4_ASAP7_75t_SL g690 ( .A(n_606), .Y(n_690) );
NOR2x1_ASAP7_75t_L g607 ( .A(n_608), .B(n_621), .Y(n_607) );
NAND4xp25_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .C(n_613), .D(n_616), .Y(n_608) );
BUFx2_ASAP7_75t_L g1056 ( .A(n_614), .Y(n_1056) );
BUFx3_ASAP7_75t_L g720 ( .A(n_615), .Y(n_720) );
INVx3_ASAP7_75t_L g1310 ( .A(n_615), .Y(n_1310) );
INVx1_ASAP7_75t_L g673 ( .A(n_617), .Y(n_673) );
INVx2_ASAP7_75t_L g823 ( .A(n_617), .Y(n_823) );
BUFx3_ASAP7_75t_L g1350 ( .A(n_617), .Y(n_1350) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g1003 ( .A(n_620), .B(n_1004), .Y(n_1003) );
NAND4xp25_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .C(n_628), .D(n_631), .Y(n_621) );
HB1xp67_ASAP7_75t_L g1322 ( .A(n_623), .Y(n_1322) );
BUFx2_ASAP7_75t_SL g1041 ( .A(n_625), .Y(n_1041) );
BUFx4f_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
BUFx2_ASAP7_75t_SL g1040 ( .A(n_630), .Y(n_1040) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B1(n_666), .B2(n_667), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g783 ( .A(n_638), .Y(n_783) );
AO21x2_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_649), .B(n_663), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_645), .B(n_647), .Y(n_644) );
BUFx3_ASAP7_75t_L g805 ( .A(n_646), .Y(n_805) );
INVx1_ASAP7_75t_L g909 ( .A(n_646), .Y(n_909) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_650), .B(n_658), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .Y(n_650) );
HB1xp67_ASAP7_75t_L g806 ( .A(n_652), .Y(n_806) );
INVx2_ASAP7_75t_L g959 ( .A(n_652), .Y(n_959) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
BUFx6f_ASAP7_75t_L g709 ( .A(n_655), .Y(n_709) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g988 ( .A(n_657), .B(n_989), .Y(n_988) );
NAND2x1_ASAP7_75t_SL g658 ( .A(n_659), .B(n_661), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
XNOR2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
NOR2xp67_ASAP7_75t_L g669 ( .A(n_670), .B(n_680), .Y(n_669) );
NAND3xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_676), .C(n_678), .Y(n_670) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g851 ( .A(n_675), .Y(n_851) );
NAND4xp25_ASAP7_75t_L g680 ( .A(n_681), .B(n_684), .C(n_686), .D(n_688), .Y(n_680) );
BUFx4f_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
BUFx3_ASAP7_75t_L g1038 ( .A(n_687), .Y(n_1038) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
XNOR2xp5_ASAP7_75t_L g692 ( .A(n_693), .B(n_781), .Y(n_692) );
XNOR2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_762), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B1(n_741), .B2(n_761), .Y(n_694) );
INVx2_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
XOR2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_740), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_698), .B(n_721), .Y(n_697) );
NOR3xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_705), .C(n_713), .Y(n_698) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
BUFx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g1058 ( .A(n_704), .Y(n_1058) );
OAI21xp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_707), .B(n_710), .Y(n_705) );
INVx2_ASAP7_75t_SL g1046 ( .A(n_707), .Y(n_1046) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g866 ( .A(n_709), .Y(n_866) );
INVx2_ASAP7_75t_L g1024 ( .A(n_709), .Y(n_1024) );
INVx1_ASAP7_75t_L g1050 ( .A(n_711), .Y(n_1050) );
INVx4_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g776 ( .A(n_712), .B(n_777), .Y(n_776) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B1(n_718), .B2(n_719), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
BUFx3_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NOR2xp67_ASAP7_75t_L g721 ( .A(n_722), .B(n_728), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_726), .Y(n_722) );
BUFx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_734), .Y(n_728) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
BUFx6f_ASAP7_75t_L g801 ( .A(n_732), .Y(n_801) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
BUFx3_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g761 ( .A(n_741), .Y(n_761) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
XNOR2x1_ASAP7_75t_L g742 ( .A(n_743), .B(n_760), .Y(n_742) );
OR2x2_ASAP7_75t_L g743 ( .A(n_744), .B(n_754), .Y(n_743) );
NAND4xp25_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .C(n_747), .D(n_752), .Y(n_744) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g937 ( .A(n_749), .Y(n_937) );
INVx1_ASAP7_75t_L g1315 ( .A(n_753), .Y(n_1315) );
NAND4xp25_ASAP7_75t_L g754 ( .A(n_755), .B(n_757), .C(n_758), .D(n_759), .Y(n_754) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVxp33_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g1030 ( .A(n_765), .Y(n_1030) );
XOR2x2_ASAP7_75t_L g765 ( .A(n_766), .B(n_780), .Y(n_765) );
NOR2xp67_ASAP7_75t_L g766 ( .A(n_767), .B(n_772), .Y(n_766) );
NAND4xp25_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .C(n_770), .D(n_771), .Y(n_767) );
NAND4xp25_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .C(n_775), .D(n_778), .Y(n_772) );
XNOR2x1_ASAP7_75t_L g781 ( .A(n_782), .B(n_784), .Y(n_781) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_786), .B1(n_809), .B2(n_810), .Y(n_784) );
INVxp67_ASAP7_75t_SL g785 ( .A(n_786), .Y(n_785) );
XNOR2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
NAND3xp33_ASAP7_75t_L g788 ( .A(n_789), .B(n_800), .C(n_804), .Y(n_788) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_793), .B(n_795), .Y(n_792) );
INVx2_ASAP7_75t_L g1312 ( .A(n_794), .Y(n_1312) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
XNOR2x1_ASAP7_75t_L g810 ( .A(n_811), .B(n_812), .Y(n_810) );
NOR2x1_ASAP7_75t_L g812 ( .A(n_813), .B(n_818), .Y(n_812) );
NAND4xp25_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .C(n_816), .D(n_817), .Y(n_813) );
NAND3xp33_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .C(n_821), .Y(n_818) );
INVx2_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
OAI21xp5_ASAP7_75t_L g824 ( .A1(n_825), .A2(n_826), .B(n_828), .Y(n_824) );
INVx4_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
XNOR2x1_ASAP7_75t_L g829 ( .A(n_830), .B(n_968), .Y(n_829) );
XNOR2xp5_ASAP7_75t_L g830 ( .A(n_831), .B(n_879), .Y(n_830) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_858), .B1(n_877), .B2(n_878), .Y(n_831) );
INVx1_ASAP7_75t_L g877 ( .A(n_832), .Y(n_877) );
HB1xp67_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
HB1xp67_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
OAI21xp5_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_836), .B(n_852), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_835), .B(n_845), .Y(n_855) );
NOR2xp67_ASAP7_75t_L g836 ( .A(n_837), .B(n_843), .Y(n_836) );
INVx1_ASAP7_75t_L g853 ( .A(n_837), .Y(n_853) );
NAND4xp25_ASAP7_75t_L g837 ( .A(n_838), .B(n_839), .C(n_840), .D(n_842), .Y(n_837) );
NAND4xp25_ASAP7_75t_L g843 ( .A(n_844), .B(n_845), .C(n_847), .D(n_848), .Y(n_843) );
INVx1_ASAP7_75t_L g856 ( .A(n_844), .Y(n_856) );
INVx1_ASAP7_75t_L g1048 ( .A(n_846), .Y(n_1048) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_847), .B(n_848), .Y(n_857) );
NOR2xp33_ASAP7_75t_L g849 ( .A(n_850), .B(n_851), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_853), .B(n_854), .Y(n_852) );
NOR3xp33_ASAP7_75t_L g854 ( .A(n_855), .B(n_856), .C(n_857), .Y(n_854) );
INVx2_ASAP7_75t_L g878 ( .A(n_858), .Y(n_878) );
NAND4xp75_ASAP7_75t_L g859 ( .A(n_860), .B(n_863), .C(n_870), .D(n_873), .Y(n_859) );
AND2x2_ASAP7_75t_L g860 ( .A(n_861), .B(n_862), .Y(n_860) );
OA21x2_ASAP7_75t_L g863 ( .A1(n_864), .A2(n_865), .B(n_867), .Y(n_863) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
AND2x2_ASAP7_75t_L g870 ( .A(n_871), .B(n_872), .Y(n_870) );
AND2x2_ASAP7_75t_L g873 ( .A(n_874), .B(n_875), .Y(n_873) );
AOI22xp5_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_881), .B1(n_944), .B2(n_967), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_882), .A2(n_883), .B1(n_926), .B2(n_927), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
XNOR2xp5_ASAP7_75t_L g883 ( .A(n_884), .B(n_898), .Y(n_883) );
INVx1_ASAP7_75t_L g896 ( .A(n_885), .Y(n_896) );
NAND3xp33_ASAP7_75t_L g885 ( .A(n_886), .B(n_891), .C(n_894), .Y(n_885) );
AND4x1_ASAP7_75t_L g886 ( .A(n_887), .B(n_888), .C(n_889), .D(n_890), .Y(n_886) );
NOR2x1_ASAP7_75t_L g899 ( .A(n_900), .B(n_910), .Y(n_899) );
NAND3xp33_ASAP7_75t_L g900 ( .A(n_901), .B(n_906), .C(n_907), .Y(n_900) );
INVx1_ASAP7_75t_L g924 ( .A(n_901), .Y(n_924) );
INVx2_ASAP7_75t_SL g902 ( .A(n_903), .Y(n_902) );
INVx2_ASAP7_75t_SL g986 ( .A(n_903), .Y(n_986) );
INVxp67_ASAP7_75t_SL g925 ( .A(n_906), .Y(n_925) );
INVx1_ASAP7_75t_L g921 ( .A(n_907), .Y(n_921) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_911), .B(n_915), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
NOR3xp33_ASAP7_75t_L g920 ( .A(n_912), .B(n_921), .C(n_922), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_913), .B(n_914), .Y(n_912) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
NOR3xp33_ASAP7_75t_L g923 ( .A(n_916), .B(n_924), .C(n_925), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_917), .B(n_918), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_920), .B(n_923), .Y(n_919) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
XNOR2xp5_ASAP7_75t_L g928 ( .A(n_929), .B(n_931), .Y(n_928) );
CKINVDCx5p33_ASAP7_75t_R g929 ( .A(n_930), .Y(n_929) );
NOR2x1_ASAP7_75t_L g931 ( .A(n_932), .B(n_939), .Y(n_931) );
NAND4xp25_ASAP7_75t_L g932 ( .A(n_933), .B(n_935), .C(n_936), .D(n_938), .Y(n_932) );
NAND4xp25_ASAP7_75t_L g939 ( .A(n_940), .B(n_941), .C(n_942), .D(n_943), .Y(n_939) );
INVx2_ASAP7_75t_L g967 ( .A(n_944), .Y(n_967) );
AO21x2_ASAP7_75t_L g944 ( .A1(n_945), .A2(n_946), .B(n_966), .Y(n_944) );
NOR3xp33_ASAP7_75t_L g966 ( .A(n_945), .B(n_948), .C(n_954), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_947), .B(n_953), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
NAND4xp25_ASAP7_75t_SL g948 ( .A(n_949), .B(n_950), .C(n_951), .D(n_952), .Y(n_948) );
INVx1_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
NAND3xp33_ASAP7_75t_L g954 ( .A(n_955), .B(n_957), .C(n_960), .Y(n_954) );
INVx2_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
OAI21xp5_ASAP7_75t_SL g961 ( .A1(n_962), .A2(n_964), .B(n_965), .Y(n_961) );
INVxp67_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
OA22x2_ASAP7_75t_L g968 ( .A1(n_969), .A2(n_1006), .B1(n_1062), .B2(n_1063), .Y(n_968) );
INVx1_ASAP7_75t_L g1062 ( .A(n_969), .Y(n_1062) );
HB1xp67_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
XNOR2xp5_ASAP7_75t_L g970 ( .A(n_971), .B(n_991), .Y(n_970) );
XNOR2x1_ASAP7_75t_L g971 ( .A(n_972), .B(n_990), .Y(n_971) );
NOR4xp75_ASAP7_75t_L g972 ( .A(n_973), .B(n_976), .C(n_980), .D(n_984), .Y(n_972) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_974), .B(n_975), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g976 ( .A(n_977), .B(n_979), .Y(n_976) );
BUFx2_ASAP7_75t_L g1320 ( .A(n_978), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_981), .B(n_983), .Y(n_980) );
NAND2xp5_ASAP7_75t_SL g984 ( .A(n_985), .B(n_987), .Y(n_984) );
NOR2x1_ASAP7_75t_L g992 ( .A(n_993), .B(n_998), .Y(n_992) );
NAND4xp25_ASAP7_75t_L g993 ( .A(n_994), .B(n_995), .C(n_996), .D(n_997), .Y(n_993) );
NAND3xp33_ASAP7_75t_L g998 ( .A(n_999), .B(n_1000), .C(n_1005), .Y(n_998) );
INVx2_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
AOI22xp5_ASAP7_75t_L g1006 ( .A1(n_1007), .A2(n_1008), .B1(n_1031), .B2(n_1061), .Y(n_1006) );
OAI22xp5_ASAP7_75t_L g1063 ( .A1(n_1007), .A2(n_1061), .B1(n_1064), .B2(n_1065), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1007), .Y(n_1064) );
INVx2_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
XNOR2x1_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1030), .Y(n_1008) );
NAND4xp25_ASAP7_75t_L g1027 ( .A(n_1011), .B(n_1012), .C(n_1014), .D(n_1023), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_1013), .B(n_1025), .Y(n_1029) );
NAND3xp33_ASAP7_75t_L g1015 ( .A(n_1016), .B(n_1023), .C(n_1025), .Y(n_1015) );
INVxp67_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
OR2x2_ASAP7_75t_L g1028 ( .A(n_1017), .B(n_1029), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1021), .Y(n_1017) );
NOR2x1_ASAP7_75t_L g1026 ( .A(n_1027), .B(n_1028), .Y(n_1026) );
INVx4_ASAP7_75t_L g1061 ( .A(n_1031), .Y(n_1061) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1032), .Y(n_1059) );
NOR2x1_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1044), .Y(n_1032) );
NAND4xp25_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1036), .C(n_1039), .D(n_1042), .Y(n_1033) );
NAND3xp33_ASAP7_75t_L g1044 ( .A(n_1045), .B(n_1052), .C(n_1055), .Y(n_1044) );
OAI22xp5_ASAP7_75t_L g1047 ( .A1(n_1048), .A2(n_1049), .B1(n_1050), .B2(n_1051), .Y(n_1047) );
INVx2_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
OAI221xp5_ASAP7_75t_L g1132 ( .A1(n_1060), .A2(n_1074), .B1(n_1081), .B2(n_1133), .C(n_1134), .Y(n_1132) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1061), .Y(n_1065) );
OAI221xp5_ASAP7_75t_L g1066 ( .A1(n_1067), .A2(n_1301), .B1(n_1303), .B2(n_1329), .C(n_1334), .Y(n_1066) );
AND5x1_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1248), .C(n_1287), .D(n_1291), .E(n_1294), .Y(n_1067) );
AOI321xp33_ASAP7_75t_L g1068 ( .A1(n_1069), .A2(n_1130), .A3(n_1162), .B1(n_1191), .B2(n_1198), .C(n_1219), .Y(n_1068) );
A2O1A1Ixp33_ASAP7_75t_L g1069 ( .A1(n_1070), .A2(n_1135), .B(n_1140), .C(n_1150), .Y(n_1069) );
AOI211xp5_ASAP7_75t_L g1070 ( .A1(n_1071), .A2(n_1099), .B(n_1118), .C(n_1125), .Y(n_1070) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1071), .Y(n_1216) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1092), .Y(n_1071) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1072), .Y(n_1136) );
INVx2_ASAP7_75t_L g1143 ( .A(n_1072), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1072), .B(n_1127), .Y(n_1161) );
OR2x2_ASAP7_75t_L g1188 ( .A(n_1072), .B(n_1127), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1072), .B(n_1093), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1072), .B(n_1213), .Y(n_1271) );
OR2x2_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1084), .Y(n_1072) );
OAI22xp5_ASAP7_75t_L g1073 ( .A1(n_1074), .A2(n_1080), .B1(n_1081), .B2(n_1083), .Y(n_1073) );
INVx3_ASAP7_75t_L g1074 ( .A(n_1075), .Y(n_1074) );
AND2x4_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1078), .Y(n_1075) );
AND2x4_ASAP7_75t_L g1086 ( .A(n_1076), .B(n_1087), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1076), .B(n_1087), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1104 ( .A(n_1076), .B(n_1087), .Y(n_1104) );
NAND2xp5_ASAP7_75t_L g1081 ( .A(n_1078), .B(n_1082), .Y(n_1081) );
AND2x4_ASAP7_75t_L g1095 ( .A(n_1078), .B(n_1082), .Y(n_1095) );
AND2x4_ASAP7_75t_L g1108 ( .A(n_1078), .B(n_1082), .Y(n_1108) );
AND2x4_ASAP7_75t_L g1090 ( .A(n_1082), .B(n_1087), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_1082), .B(n_1087), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1082), .B(n_1087), .Y(n_1114) );
OAI22xp5_ASAP7_75t_L g1084 ( .A1(n_1085), .A2(n_1088), .B1(n_1089), .B2(n_1091), .Y(n_1084) );
INVx3_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
BUFx2_ASAP7_75t_L g1302 ( .A(n_1086), .Y(n_1302) );
NOR2xp33_ASAP7_75t_L g1353 ( .A(n_1088), .B(n_1344), .Y(n_1353) );
INVx2_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
INVx2_ASAP7_75t_L g1120 ( .A(n_1092), .Y(n_1120) );
NOR2x1_ASAP7_75t_L g1138 ( .A(n_1092), .B(n_1139), .Y(n_1138) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_1092), .B(n_1146), .Y(n_1145) );
BUFx6f_ASAP7_75t_L g1153 ( .A(n_1092), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1092), .B(n_1123), .Y(n_1159) );
NAND2xp5_ASAP7_75t_SL g1182 ( .A(n_1092), .B(n_1183), .Y(n_1182) );
NAND2xp5_ASAP7_75t_SL g1206 ( .A(n_1092), .B(n_1207), .Y(n_1206) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1092), .Y(n_1230) );
INVx2_ASAP7_75t_L g1238 ( .A(n_1092), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1092), .B(n_1136), .Y(n_1262) );
INVx4_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
OR2x2_ASAP7_75t_L g1172 ( .A(n_1093), .B(n_1100), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1096), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1099), .B(n_1120), .Y(n_1266) );
NAND2xp5_ASAP7_75t_L g1268 ( .A(n_1099), .B(n_1269), .Y(n_1268) );
INVx2_ASAP7_75t_SL g1286 ( .A(n_1099), .Y(n_1286) );
AND2x4_ASAP7_75t_L g1099 ( .A(n_1100), .B(n_1109), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1100), .B(n_1155), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1100), .B(n_1115), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1100), .B(n_1123), .Y(n_1251) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
INVx1_ASAP7_75t_SL g1101 ( .A(n_1102), .Y(n_1101) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1102), .Y(n_1122) );
OR2x2_ASAP7_75t_L g1176 ( .A(n_1102), .B(n_1110), .Y(n_1176) );
OR2x2_ASAP7_75t_L g1179 ( .A(n_1102), .B(n_1139), .Y(n_1179) );
NAND2xp5_ASAP7_75t_L g1190 ( .A(n_1102), .B(n_1183), .Y(n_1190) );
NAND2xp5_ASAP7_75t_L g1200 ( .A(n_1102), .B(n_1159), .Y(n_1200) );
NAND2xp5_ASAP7_75t_L g1208 ( .A(n_1102), .B(n_1111), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1102), .B(n_1124), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1105), .Y(n_1102) );
NAND2xp5_ASAP7_75t_L g1263 ( .A(n_1109), .B(n_1264), .Y(n_1263) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
NAND2xp5_ASAP7_75t_L g1280 ( .A(n_1110), .B(n_1215), .Y(n_1280) );
OR2x2_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1115), .Y(n_1110) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1111), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1111), .B(n_1115), .Y(n_1155) );
AOI322xp5_ASAP7_75t_L g1294 ( .A1(n_1111), .A2(n_1209), .A3(n_1221), .B1(n_1264), .B2(n_1295), .C1(n_1297), .C2(n_1298), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1112), .B(n_1113), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_1115), .B(n_1124), .Y(n_1123) );
OR2x2_ASAP7_75t_L g1139 ( .A(n_1115), .B(n_1124), .Y(n_1139) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1115), .Y(n_1147) );
NAND2xp5_ASAP7_75t_L g1244 ( .A(n_1115), .B(n_1122), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1116), .B(n_1117), .Y(n_1115) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
NOR2xp33_ASAP7_75t_L g1290 ( .A(n_1119), .B(n_1141), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1121), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1120), .B(n_1175), .Y(n_1174) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1120), .Y(n_1269) );
NOR2xp33_ASAP7_75t_L g1165 ( .A(n_1121), .B(n_1166), .Y(n_1165) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1121), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1123), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1122), .B(n_1138), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1122), .B(n_1147), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1122), .B(n_1155), .Y(n_1154) );
NOR2x1_ASAP7_75t_R g1255 ( .A(n_1122), .B(n_1182), .Y(n_1255) );
NOR2xp33_ASAP7_75t_L g1279 ( .A(n_1122), .B(n_1280), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1122), .B(n_1124), .Y(n_1300) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1123), .Y(n_1171) );
NAND2xp5_ASAP7_75t_L g1253 ( .A(n_1123), .B(n_1229), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1130), .Y(n_1125) );
AOI211xp5_ASAP7_75t_L g1140 ( .A1(n_1126), .A2(n_1141), .B(n_1144), .C(n_1148), .Y(n_1140) );
CKINVDCx14_ASAP7_75t_R g1185 ( .A(n_1126), .Y(n_1185) );
OAI221xp5_ASAP7_75t_L g1219 ( .A1(n_1126), .A2(n_1173), .B1(n_1220), .B2(n_1227), .C(n_1228), .Y(n_1219) );
OAI21xp5_ASAP7_75t_L g1287 ( .A1(n_1126), .A2(n_1288), .B(n_1290), .Y(n_1287) );
INVx2_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1127), .B(n_1143), .Y(n_1167) );
HB1xp67_ASAP7_75t_L g1180 ( .A(n_1127), .Y(n_1180) );
OR2x2_ASAP7_75t_L g1210 ( .A(n_1127), .B(n_1195), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1127), .B(n_1194), .Y(n_1213) );
OR2x2_ASAP7_75t_L g1231 ( .A(n_1127), .B(n_1143), .Y(n_1231) );
OR2x2_ASAP7_75t_L g1242 ( .A(n_1127), .B(n_1194), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1127), .B(n_1193), .Y(n_1277) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_1128), .B(n_1129), .Y(n_1127) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
NOR2xp33_ASAP7_75t_L g1297 ( .A(n_1131), .B(n_1227), .Y(n_1297) );
INVx2_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
HB1xp67_ASAP7_75t_L g1149 ( .A(n_1132), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1132), .B(n_1241), .Y(n_1240) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_1132), .B(n_1227), .Y(n_1245) );
NAND2xp5_ASAP7_75t_L g1135 ( .A(n_1136), .B(n_1137), .Y(n_1135) );
INVx2_ASAP7_75t_L g1169 ( .A(n_1136), .Y(n_1169) );
O2A1O1Ixp33_ASAP7_75t_SL g1283 ( .A1(n_1136), .A2(n_1245), .B(n_1284), .C(n_1286), .Y(n_1283) );
NAND2xp5_ASAP7_75t_L g1293 ( .A(n_1136), .B(n_1266), .Y(n_1293) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1138), .Y(n_1199) );
AOI22xp5_ASAP7_75t_L g1270 ( .A1(n_1138), .A2(n_1236), .B1(n_1271), .B2(n_1272), .Y(n_1270) );
INVx3_ASAP7_75t_SL g1183 ( .A(n_1139), .Y(n_1183) );
AOI21xp5_ASAP7_75t_L g1220 ( .A1(n_1141), .A2(n_1221), .B(n_1224), .Y(n_1220) );
INVx2_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
AOI21xp5_ASAP7_75t_L g1150 ( .A1(n_1142), .A2(n_1151), .B(n_1156), .Y(n_1150) );
NAND2xp5_ASAP7_75t_L g1173 ( .A(n_1142), .B(n_1174), .Y(n_1173) );
NOR2xp67_ASAP7_75t_SL g1249 ( .A(n_1142), .B(n_1250), .Y(n_1249) );
INVx2_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1143), .B(n_1203), .Y(n_1202) );
NOR2xp33_ASAP7_75t_L g1272 ( .A(n_1143), .B(n_1210), .Y(n_1272) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
NOR2xp33_ASAP7_75t_L g1211 ( .A(n_1145), .B(n_1212), .Y(n_1211) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1146), .Y(n_1233) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1148), .B(n_1192), .Y(n_1191) );
AOI221xp5_ASAP7_75t_L g1248 ( .A1(n_1148), .A2(n_1241), .B1(n_1249), .B2(n_1252), .C(n_1273), .Y(n_1248) );
INVx2_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
AOI221xp5_ASAP7_75t_L g1177 ( .A1(n_1149), .A2(n_1178), .B1(n_1180), .B2(n_1181), .C(n_1184), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1154), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g1296 ( .A(n_1152), .B(n_1167), .Y(n_1296) );
INVx2_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
OAI321xp33_ASAP7_75t_L g1256 ( .A1(n_1153), .A2(n_1201), .A3(n_1257), .B1(n_1259), .B2(n_1260), .C(n_1261), .Y(n_1256) );
OAI21xp5_ASAP7_75t_L g1284 ( .A1(n_1153), .A2(n_1227), .B(n_1285), .Y(n_1284) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1154), .Y(n_1157) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1155), .Y(n_1215) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1155), .B(n_1223), .Y(n_1222) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_1155), .B(n_1238), .Y(n_1237) );
AOI21xp33_ASAP7_75t_L g1156 ( .A1(n_1157), .A2(n_1158), .B(n_1160), .Y(n_1156) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
OAI21xp5_ASAP7_75t_SL g1267 ( .A1(n_1160), .A2(n_1268), .B(n_1270), .Y(n_1267) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
NAND2xp5_ASAP7_75t_L g1282 ( .A(n_1161), .B(n_1238), .Y(n_1282) );
NAND4xp25_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1173), .C(n_1177), .D(n_1186), .Y(n_1162) );
AOI21xp5_ASAP7_75t_L g1163 ( .A1(n_1164), .A2(n_1167), .B(n_1168), .Y(n_1163) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
O2A1O1Ixp33_ASAP7_75t_L g1265 ( .A1(n_1167), .A2(n_1226), .B(n_1266), .C(n_1267), .Y(n_1265) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1168), .Y(n_1275) );
NOR2xp33_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1170), .Y(n_1168) );
NAND2xp5_ASAP7_75t_L g1225 ( .A(n_1169), .B(n_1226), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1259 ( .A(n_1169), .B(n_1192), .Y(n_1259) );
NOR2xp33_ASAP7_75t_L g1288 ( .A(n_1169), .B(n_1289), .Y(n_1288) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1170), .Y(n_1226) );
OR2x2_ASAP7_75t_L g1170 ( .A(n_1171), .B(n_1172), .Y(n_1170) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1172), .Y(n_1223) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1174), .Y(n_1274) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
NAND2xp33_ASAP7_75t_L g1298 ( .A(n_1179), .B(n_1299), .Y(n_1298) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
CKINVDCx14_ASAP7_75t_R g1184 ( .A(n_1185), .Y(n_1184) );
NAND2xp5_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1189), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_1187), .B(n_1218), .Y(n_1264) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1190), .Y(n_1189) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1195), .Y(n_1203) );
NAND2xp5_ASAP7_75t_L g1195 ( .A(n_1196), .B(n_1197), .Y(n_1195) );
A2O1A1Ixp33_ASAP7_75t_L g1198 ( .A1(n_1199), .A2(n_1200), .B(n_1201), .C(n_1204), .Y(n_1198) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
BUFx3_ASAP7_75t_L g1218 ( .A(n_1203), .Y(n_1218) );
INVx2_ASAP7_75t_L g1227 ( .A(n_1203), .Y(n_1227) );
AOI211xp5_ASAP7_75t_L g1204 ( .A1(n_1205), .A2(n_1209), .B(n_1211), .C(n_1214), .Y(n_1204) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1206), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g1261 ( .A(n_1207), .B(n_1262), .Y(n_1261) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
NOR2xp33_ASAP7_75t_L g1292 ( .A(n_1212), .B(n_1293), .Y(n_1292) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
AOI21xp5_ASAP7_75t_L g1254 ( .A1(n_1213), .A2(n_1255), .B(n_1256), .Y(n_1254) );
NOR3xp33_ASAP7_75t_L g1214 ( .A(n_1215), .B(n_1216), .C(n_1217), .Y(n_1214) );
AOI211xp5_ASAP7_75t_SL g1243 ( .A1(n_1215), .A2(n_1244), .B(n_1245), .C(n_1246), .Y(n_1243) );
INVx2_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
AOI21xp5_ASAP7_75t_L g1232 ( .A1(n_1218), .A2(n_1233), .B(n_1234), .Y(n_1232) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
AOI31xp33_ASAP7_75t_L g1278 ( .A1(n_1227), .A2(n_1279), .A3(n_1281), .B(n_1283), .Y(n_1278) );
AOI221xp5_ASAP7_75t_L g1228 ( .A1(n_1229), .A2(n_1232), .B1(n_1236), .B2(n_1239), .C(n_1243), .Y(n_1228) );
NOR2xp33_ASAP7_75t_L g1229 ( .A(n_1230), .B(n_1231), .Y(n_1229) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1231), .Y(n_1285) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
NAND2xp67_ASAP7_75t_L g1250 ( .A(n_1238), .B(n_1251), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1299 ( .A(n_1238), .B(n_1300), .Y(n_1299) );
INVxp67_ASAP7_75t_SL g1239 ( .A(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
NAND4xp25_ASAP7_75t_L g1252 ( .A(n_1253), .B(n_1254), .C(n_1263), .D(n_1265), .Y(n_1252) );
INVxp67_ASAP7_75t_SL g1289 ( .A(n_1255), .Y(n_1289) );
CKINVDCx20_ASAP7_75t_R g1257 ( .A(n_1258), .Y(n_1257) );
A2O1A1Ixp33_ASAP7_75t_L g1273 ( .A1(n_1274), .A2(n_1275), .B(n_1276), .C(n_1278), .Y(n_1273) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
INVxp67_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
CKINVDCx5p33_ASAP7_75t_R g1301 ( .A(n_1302), .Y(n_1301) );
INVxp67_ASAP7_75t_SL g1328 ( .A(n_1304), .Y(n_1328) );
AND2x4_ASAP7_75t_L g1304 ( .A(n_1305), .B(n_1317), .Y(n_1304) );
NOR3xp33_ASAP7_75t_L g1305 ( .A(n_1306), .B(n_1308), .C(n_1313), .Y(n_1305) );
OAI22xp5_ASAP7_75t_L g1308 ( .A1(n_1309), .A2(n_1310), .B1(n_1311), .B2(n_1312), .Y(n_1308) );
OAI21xp33_ASAP7_75t_L g1313 ( .A1(n_1314), .A2(n_1315), .B(n_1316), .Y(n_1313) );
NOR2x1_ASAP7_75t_L g1317 ( .A(n_1318), .B(n_1323), .Y(n_1317) );
NAND2xp5_ASAP7_75t_L g1318 ( .A(n_1319), .B(n_1321), .Y(n_1318) );
NAND2xp5_ASAP7_75t_L g1323 ( .A(n_1324), .B(n_1326), .Y(n_1323) );
CKINVDCx5p33_ASAP7_75t_R g1329 ( .A(n_1330), .Y(n_1329) );
HB1xp67_ASAP7_75t_SL g1330 ( .A(n_1331), .Y(n_1330) );
BUFx2_ASAP7_75t_SL g1331 ( .A(n_1332), .Y(n_1331) );
BUFx2_ASAP7_75t_L g1335 ( .A(n_1336), .Y(n_1335) );
HB1xp67_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
NOR2xp33_ASAP7_75t_L g1338 ( .A(n_1339), .B(n_1344), .Y(n_1338) );
INVxp67_ASAP7_75t_L g1354 ( .A(n_1339), .Y(n_1354) );
NAND4xp25_ASAP7_75t_L g1339 ( .A(n_1340), .B(n_1341), .C(n_1342), .D(n_1343), .Y(n_1339) );
NAND4xp25_ASAP7_75t_L g1344 ( .A(n_1345), .B(n_1348), .C(n_1349), .D(n_1351), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1352 ( .A(n_1353), .B(n_1354), .Y(n_1352) );
BUFx3_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
CKINVDCx5p33_ASAP7_75t_R g1359 ( .A(n_1360), .Y(n_1359) );
endmodule