module fake_jpeg_17503_n_331 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_331);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx8_ASAP7_75t_SL g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_38),
.B(n_39),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_14),
.B(n_1),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_40),
.B(n_3),
.Y(n_116)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_43),
.Y(n_71)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_11),
.B1(n_9),
.B2(n_3),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_46),
.A2(n_18),
.B1(n_22),
.B2(n_13),
.Y(n_90)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_21),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_53),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_16),
.B(n_11),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_60),
.Y(n_81)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_16),
.B(n_1),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_22),
.B1(n_13),
.B2(n_31),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_64),
.Y(n_87)
);

NAND2xp33_ASAP7_75t_SL g63 ( 
.A(n_36),
.B(n_33),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_63),
.A2(n_29),
.B(n_37),
.C(n_34),
.Y(n_106)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_33),
.B(n_1),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_67),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_30),
.Y(n_101)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_69),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_70),
.A2(n_72),
.B1(n_75),
.B2(n_85),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_42),
.A2(n_19),
.B1(n_24),
.B2(n_35),
.Y(n_72)
);

AOI32xp33_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_27),
.A3(n_35),
.B1(n_17),
.B2(n_23),
.Y(n_73)
);

AOI32xp33_ASAP7_75t_L g140 ( 
.A1(n_73),
.A2(n_6),
.A3(n_8),
.B1(n_90),
.B2(n_91),
.Y(n_140)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_74),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_58),
.A2(n_24),
.B1(n_35),
.B2(n_23),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_24),
.C(n_22),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_92),
.Y(n_121)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_82),
.A2(n_100),
.B1(n_8),
.B2(n_98),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_50),
.A2(n_24),
.B1(n_23),
.B2(n_20),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_64),
.A2(n_27),
.B1(n_17),
.B2(n_20),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_86),
.A2(n_96),
.B1(n_111),
.B2(n_112),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_90),
.A2(n_4),
.B(n_5),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_46),
.B(n_20),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_91),
.B(n_97),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_18),
.C(n_17),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_56),
.A2(n_16),
.B1(n_18),
.B2(n_37),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_93),
.A2(n_113),
.B1(n_114),
.B2(n_30),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_34),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_99),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_43),
.A2(n_26),
.B1(n_34),
.B2(n_31),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_38),
.B(n_26),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_48),
.B(n_37),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_110),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_106),
.Y(n_139)
);

CKINVDCx12_ASAP7_75t_R g110 ( 
.A(n_67),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_49),
.A2(n_25),
.B1(n_29),
.B2(n_28),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_54),
.A2(n_25),
.B1(n_29),
.B2(n_28),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_45),
.A2(n_25),
.B1(n_28),
.B2(n_26),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_53),
.A2(n_31),
.B1(n_30),
.B2(n_5),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_116),
.B(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_118),
.Y(n_188)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_119),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_4),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_136),
.Y(n_165)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_122),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_80),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_123),
.B(n_127),
.Y(n_166)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_124),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_125),
.B(n_146),
.Y(n_189)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_126),
.B(n_132),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_62),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_129),
.B(n_130),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_77),
.B(n_4),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_116),
.B(n_81),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_87),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_135),
.Y(n_181)
);

O2A1O1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_134),
.A2(n_157),
.B(n_136),
.C(n_144),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_89),
.B(n_8),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_5),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_92),
.B(n_6),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_137),
.B(n_138),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_102),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_SL g173 ( 
.A(n_140),
.B(n_155),
.C(n_120),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_142),
.B(n_149),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_79),
.B(n_8),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_146),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_70),
.A2(n_105),
.B1(n_100),
.B2(n_98),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_145),
.A2(n_157),
.B1(n_152),
.B2(n_148),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_103),
.B(n_78),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_147),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_88),
.B(n_71),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_148),
.A2(n_152),
.B(n_161),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_69),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_88),
.B(n_71),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_94),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_154),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_69),
.B(n_109),
.Y(n_154)
);

NOR2xp67_ASAP7_75t_R g155 ( 
.A(n_69),
.B(n_83),
.Y(n_155)
);

AO22x1_ASAP7_75t_L g157 ( 
.A1(n_109),
.A2(n_107),
.B1(n_108),
.B2(n_83),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_74),
.A2(n_82),
.B1(n_107),
.B2(n_108),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_159),
.A2(n_118),
.B1(n_119),
.B2(n_126),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_83),
.B(n_94),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_121),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_91),
.A2(n_46),
.B(n_75),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_80),
.Y(n_162)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_123),
.C(n_128),
.Y(n_190)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_158),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_167),
.Y(n_213)
);

INVxp33_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_121),
.A2(n_143),
.B(n_151),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_171),
.A2(n_200),
.B(n_174),
.Y(n_203)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_172),
.B(n_187),
.Y(n_219)
);

OR2x4_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_189),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_121),
.A2(n_139),
.B1(n_131),
.B2(n_140),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_174),
.A2(n_179),
.B1(n_183),
.B2(n_195),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_175),
.B(n_165),
.Y(n_216)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_177),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_117),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_182),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_134),
.B1(n_124),
.B2(n_150),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_180),
.A2(n_171),
.B(n_166),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_131),
.B(n_150),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_145),
.A2(n_127),
.B1(n_142),
.B2(n_122),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_184),
.A2(n_168),
.B(n_198),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_189),
.B(n_164),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_190),
.B(n_176),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_148),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_198),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_152),
.B(n_157),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_156),
.A2(n_139),
.B1(n_161),
.B2(n_140),
.Y(n_199)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_172),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_117),
.B(n_124),
.C(n_144),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_164),
.C(n_200),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_203),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_204),
.B(n_220),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_194),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_205),
.B(n_207),
.Y(n_254)
);

INVx13_ASAP7_75t_L g207 ( 
.A(n_201),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_208),
.A2(n_216),
.B1(n_222),
.B2(n_206),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_202),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_217),
.C(n_226),
.Y(n_240)
);

OAI32xp33_ASAP7_75t_L g212 ( 
.A1(n_182),
.A2(n_179),
.A3(n_178),
.B1(n_165),
.B2(n_169),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_215),
.Y(n_237)
);

INVxp67_ASAP7_75t_SL g214 ( 
.A(n_163),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_214),
.B(n_228),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_169),
.B(n_187),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_180),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_234),
.Y(n_248)
);

AND2x6_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_173),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_221),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_188),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_227),
.Y(n_241)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_177),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_192),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_188),
.Y(n_227)
);

AND2x6_ASAP7_75t_L g229 ( 
.A(n_186),
.B(n_195),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_229),
.Y(n_244)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_231),
.B(n_233),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_185),
.B(n_183),
.C(n_193),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_236),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_181),
.B(n_170),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_196),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_168),
.A2(n_197),
.B(n_191),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_215),
.B(n_194),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_238),
.B(n_252),
.Y(n_272)
);

AND2x2_ASAP7_75t_SL g242 ( 
.A(n_210),
.B(n_218),
.Y(n_242)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_243),
.B(n_253),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_225),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_245),
.B(n_246),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_230),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_234),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_261),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_211),
.A2(n_216),
.B1(n_210),
.B2(n_229),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_250),
.A2(n_253),
.B1(n_252),
.B2(n_243),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_206),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_211),
.A2(n_216),
.B1(n_232),
.B2(n_224),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_209),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_256),
.Y(n_267)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_257),
.Y(n_281)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_219),
.Y(n_261)
);

NOR3xp33_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_208),
.C(n_221),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_262),
.B(n_268),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_256),
.C(n_247),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_264),
.B(n_265),
.C(n_276),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_217),
.C(n_203),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_259),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_223),
.Y(n_270)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_270),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_258),
.A2(n_222),
.B1(n_236),
.B2(n_220),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_271),
.A2(n_248),
.B(n_244),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_260),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_273),
.B(n_274),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_227),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_245),
.Y(n_275)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_275),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_224),
.C(n_213),
.Y(n_276)
);

NAND3xp33_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_207),
.C(n_239),
.Y(n_277)
);

OAI322xp33_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_246),
.A3(n_255),
.B1(n_251),
.B2(n_241),
.C1(n_242),
.C2(n_238),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_237),
.B(n_250),
.Y(n_278)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_278),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_237),
.B(n_244),
.Y(n_279)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_279),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_242),
.C(n_241),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_242),
.Y(n_293)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_275),
.Y(n_283)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

AO21x1_ASAP7_75t_L g284 ( 
.A1(n_272),
.A2(n_248),
.B(n_255),
.Y(n_284)
);

AO21x1_ASAP7_75t_L g307 ( 
.A1(n_284),
.A2(n_285),
.B(n_293),
.Y(n_307)
);

BUFx12_ASAP7_75t_L g287 ( 
.A(n_275),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_281),
.Y(n_301)
);

NAND4xp25_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_284),
.C(n_269),
.D(n_290),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_271),
.Y(n_305)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_266),
.Y(n_296)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_296),
.Y(n_306)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_297),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_266),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_290),
.A2(n_282),
.B1(n_263),
.B2(n_276),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_300),
.B(n_304),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_301),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_280),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_305),
.Y(n_315)
);

NAND4xp25_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_286),
.C(n_285),
.D(n_295),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_268),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_288),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_309),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_264),
.Y(n_309)
);

NAND2xp33_ASAP7_75t_R g319 ( 
.A(n_310),
.B(n_307),
.Y(n_319)
);

OAI22xp33_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_283),
.B1(n_296),
.B2(n_293),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_316),
.Y(n_320)
);

NAND4xp25_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_281),
.C(n_287),
.D(n_288),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_314),
.A2(n_312),
.B(n_263),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_307),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_318),
.A2(n_299),
.B(n_298),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_321),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_322),
.A2(n_316),
.B(n_314),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_309),
.C(n_302),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_323),
.B(n_315),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_320),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_325),
.B(n_317),
.Y(n_327)
);

AOI322xp5_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_328),
.A3(n_311),
.B1(n_313),
.B2(n_289),
.C1(n_326),
.C2(n_251),
.Y(n_329)
);

A2O1A1Ixp33_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_272),
.B(n_289),
.C(n_267),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_300),
.Y(n_331)
);


endmodule