module fake_jpeg_400_n_61 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_7),
.B(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_8),
.A2(n_0),
.B(n_1),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_17),
.A2(n_23),
.B(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_13),
.Y(n_18)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_0),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_19),
.B(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_25),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_12),
.A2(n_16),
.B1(n_9),
.B2(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_26),
.B(n_27),
.Y(n_38)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_23),
.A2(n_15),
.B1(n_11),
.B2(n_4),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_30),
.A2(n_32),
.B1(n_34),
.B2(n_39),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_19),
.A2(n_3),
.B1(n_6),
.B2(n_27),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_26),
.B1(n_30),
.B2(n_32),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_18),
.A2(n_6),
.B(n_21),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_34),
.B(n_38),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_44),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_26),
.C(n_6),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_45),
.C(n_31),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_33),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_47),
.B(n_48),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_31),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_37),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_51),
.Y(n_57)
);

BUFx12f_ASAP7_75t_SL g51 ( 
.A(n_48),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_45),
.C(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_56),
.Y(n_58)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_57),
.A2(n_51),
.B(n_52),
.Y(n_59)
);

AOI321xp33_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_55),
.A3(n_54),
.B1(n_50),
.B2(n_44),
.C(n_37),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_58),
.Y(n_61)
);


endmodule