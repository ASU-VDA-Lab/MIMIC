module fake_jpeg_8755_n_71 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_71);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_71;

wire n_61;
wire n_45;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_59;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_39;
wire n_42;
wire n_49;
wire n_38;
wire n_56;
wire n_50;
wire n_67;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_69;
wire n_40;
wire n_35;
wire n_48;
wire n_46;
wire n_44;
wire n_36;
wire n_62;
wire n_37;
wire n_43;
wire n_70;
wire n_66;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_20),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_46),
.B(n_50),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_51),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_45),
.B1(n_36),
.B2(n_37),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_43),
.B1(n_7),
.B2(n_10),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_45),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_1),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_2),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_44),
.C(n_41),
.Y(n_54)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_3),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_14),
.B1(n_17),
.B2(n_19),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_55),
.Y(n_63)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_62),
.B1(n_57),
.B2(n_22),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_63),
.B(n_64),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_56),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_21),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_67),
.A2(n_25),
.B(n_26),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_27),
.C(n_28),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_SL g70 ( 
.A1(n_69),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_32),
.Y(n_71)
);


endmodule