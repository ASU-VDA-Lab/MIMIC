module fake_jpeg_8746_n_171 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_171);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_18),
.Y(n_28)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_41),
.B(n_44),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_17),
.B1(n_12),
.B2(n_27),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_12),
.B1(n_21),
.B2(n_20),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_17),
.B1(n_22),
.B2(n_12),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_12),
.B1(n_17),
.B2(n_24),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_13),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_29),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_46),
.B(n_50),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_13),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_24),
.C(n_29),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_18),
.B(n_28),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_49),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_19),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_51),
.B(n_52),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_63),
.B1(n_69),
.B2(n_39),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_55),
.B(n_19),
.Y(n_81)
);

O2A1O1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_51),
.A2(n_28),
.B(n_26),
.C(n_36),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_66),
.B(n_28),
.Y(n_79)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_67),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_22),
.B1(n_36),
.B2(n_19),
.Y(n_63)
);

NOR3xp33_ASAP7_75t_SL g67 ( 
.A(n_41),
.B(n_21),
.C(n_14),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_48),
.A2(n_26),
.B1(n_28),
.B2(n_32),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_71),
.Y(n_97)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_72),
.A2(n_78),
.B(n_79),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_64),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_75),
.B(n_76),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_46),
.Y(n_74)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_68),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_53),
.Y(n_77)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_49),
.Y(n_78)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_83),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_26),
.C(n_49),
.Y(n_83)
);

NAND2x1_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_69),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_86),
.A2(n_93),
.B(n_95),
.Y(n_105)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_62),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_82),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_91),
.B(n_92),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp67_ASAP7_75t_SL g93 ( 
.A(n_83),
.B(n_67),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_59),
.B1(n_54),
.B2(n_61),
.Y(n_95)
);

NAND3xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_60),
.C(n_10),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_9),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_79),
.B(n_76),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_81),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_76),
.A2(n_83),
.B1(n_82),
.B2(n_71),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_74),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_110),
.C(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_108),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_103),
.A2(n_116),
.B(n_94),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_112),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_75),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_109),
.B(n_113),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_73),
.C(n_61),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_11),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_11),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_114),
.Y(n_123)
);

XNOR2x1_ASAP7_75t_SL g115 ( 
.A(n_86),
.B(n_11),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_115),
.B(n_26),
.Y(n_126)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_87),
.B(n_90),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_104),
.B(n_102),
.Y(n_131)
);

BUFx12_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_124),
.B(n_65),
.Y(n_134)
);

AO21x1_ASAP7_75t_L g125 ( 
.A1(n_115),
.A2(n_87),
.B(n_11),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_111),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_126),
.B(n_128),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_102),
.A2(n_62),
.B1(n_65),
.B2(n_45),
.Y(n_127)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_105),
.B(n_26),
.Y(n_128)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_139),
.Y(n_144)
);

OAI31xp33_ASAP7_75t_L g143 ( 
.A1(n_133),
.A2(n_136),
.A3(n_125),
.B(n_126),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_107),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_40),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_128),
.Y(n_142)
);

BUFx24_ASAP7_75t_SL g139 ( 
.A(n_122),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_123),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_141),
.B(n_1),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_147),
.Y(n_153)
);

AOI31xp67_ASAP7_75t_L g149 ( 
.A1(n_143),
.A2(n_136),
.A3(n_124),
.B(n_3),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_137),
.A2(n_119),
.B1(n_121),
.B2(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_146),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_119),
.Y(n_147)
);

AOI21x1_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_5),
.B(n_6),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_9),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_152),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_L g152 ( 
.A1(n_140),
.A2(n_19),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_1),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_2),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_154),
.Y(n_160)
);

NOR2x1_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_141),
.Y(n_155)
);

NOR4xp25_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_7),
.C(n_16),
.D(n_160),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_142),
.Y(n_156)
);

NAND3xp33_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_158),
.C(n_5),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_159),
.A2(n_147),
.B1(n_153),
.B2(n_8),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_161),
.B(n_162),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_16),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_164),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_16),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_165),
.A2(n_7),
.B(n_16),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_163),
.C(n_7),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_170),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_16),
.C(n_168),
.Y(n_170)
);


endmodule