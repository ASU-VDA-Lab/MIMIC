module fake_jpeg_6548_n_176 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_8),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g30 ( 
.A(n_27),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_36),
.Y(n_47)
);

HAxp5_ASAP7_75t_SL g32 ( 
.A(n_13),
.B(n_0),
.CON(n_32),
.SN(n_32)
);

OAI21xp33_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_33),
.B(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_24),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_51),
.B1(n_15),
.B2(n_16),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_48),
.Y(n_59)
);

CKINVDCx6p67_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_44),
.Y(n_67)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_43),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_17),
.B1(n_25),
.B2(n_16),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_13),
.B1(n_25),
.B2(n_19),
.Y(n_58)
);

NOR2x1_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_21),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_24),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_22),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_30),
.B(n_17),
.C(n_26),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_26),
.B(n_15),
.Y(n_55)
);

OAI21xp33_ASAP7_75t_SL g69 ( 
.A1(n_54),
.A2(n_39),
.B(n_19),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_11),
.Y(n_84)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_61),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_60),
.B1(n_22),
.B2(n_53),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_35),
.B1(n_29),
.B2(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_62),
.Y(n_73)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_63),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_65),
.Y(n_76)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_57),
.B(n_55),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_69),
.A2(n_73),
.B1(n_77),
.B2(n_63),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

NAND3xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_84),
.C(n_18),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_74),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_35),
.B1(n_47),
.B2(n_48),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_80),
.B1(n_83),
.B2(n_82),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_54),
.A2(n_47),
.B1(n_36),
.B2(n_29),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_40),
.B1(n_45),
.B2(n_31),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_92),
.Y(n_104)
);

AOI221xp5_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_91),
.B1(n_18),
.B2(n_67),
.C(n_37),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_79),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_40),
.B1(n_45),
.B2(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_98),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_66),
.B(n_67),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_34),
.B(n_37),
.Y(n_107)
);

OAI211xp5_ASAP7_75t_SL g110 ( 
.A1(n_96),
.A2(n_41),
.B(n_42),
.C(n_34),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_84),
.B(n_28),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_97),
.Y(n_103)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_64),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_71),
.B(n_28),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_18),
.Y(n_109)
);

NOR2xp67_ASAP7_75t_SL g101 ( 
.A(n_91),
.B(n_76),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_105),
.B(n_111),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_114),
.B(n_116),
.Y(n_127)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_110),
.A2(n_42),
.B1(n_41),
.B2(n_46),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_92),
.C(n_97),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_85),
.B1(n_98),
.B2(n_87),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_34),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_78),
.C(n_64),
.Y(n_116)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_86),
.B(n_85),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_119),
.B1(n_118),
.B2(n_120),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_106),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_125),
.Y(n_141)
);

XNOR2x1_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_94),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_103),
.C(n_108),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_104),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_110),
.A2(n_88),
.B1(n_37),
.B2(n_20),
.Y(n_126)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_107),
.Y(n_128)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_42),
.B1(n_46),
.B2(n_41),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_130),
.B1(n_102),
.B2(n_114),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_116),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_134),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_132),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_137),
.C(n_18),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_109),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_112),
.C(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_140),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_18),
.Y(n_140)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_138),
.A2(n_118),
.B(n_120),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_143),
.A2(n_149),
.B1(n_150),
.B2(n_137),
.Y(n_154)
);

NAND4xp25_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_126),
.C(n_127),
.D(n_130),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_152),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_134),
.C(n_3),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_20),
.B1(n_46),
.B2(n_4),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_136),
.A2(n_2),
.B(n_3),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_131),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_155),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_154),
.B(n_159),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_158),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_5),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_6),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_6),
.C(n_7),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_7),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_163),
.B(n_8),
.Y(n_170)
);

OAI221xp5_ASAP7_75t_L g164 ( 
.A1(n_157),
.A2(n_146),
.B1(n_143),
.B2(n_150),
.C(n_9),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_166),
.Y(n_168)
);

OAI221xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.C(n_155),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_162),
.B(n_160),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_167),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_161),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_169),
.A2(n_165),
.B(n_10),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_170),
.B(n_165),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_173),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_172),
.A2(n_168),
.B(n_10),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_174),
.Y(n_176)
);


endmodule