module fake_jpeg_32143_n_186 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_186);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_154;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_4),
.B(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_35),
.B(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_1),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_48),
.Y(n_58)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_38),
.Y(n_66)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_45),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_25),
.B(n_2),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_25),
.B(n_3),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_34),
.Y(n_72)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_49),
.B1(n_46),
.B2(n_37),
.Y(n_53)
);

OAI32xp33_ASAP7_75t_L g86 ( 
.A1(n_53),
.A2(n_55),
.A3(n_74),
.B1(n_33),
.B2(n_30),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_29),
.B1(n_32),
.B2(n_16),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_26),
.B1(n_21),
.B2(n_32),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_59),
.A2(n_67),
.B1(n_3),
.B2(n_4),
.Y(n_96)
);

OR2x2_ASAP7_75t_SL g60 ( 
.A(n_51),
.B(n_34),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_47),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_63),
.Y(n_90)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_27),
.C(n_20),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_26),
.B1(n_21),
.B2(n_23),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_20),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_L g74 ( 
.A1(n_36),
.A2(n_17),
.B(n_24),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_70),
.B(n_48),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_84),
.C(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_79),
.B(n_87),
.Y(n_103)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_35),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_83),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_18),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_43),
.C(n_41),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_85),
.Y(n_102)
);

NOR2x1p5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_98),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_27),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_23),
.B1(n_41),
.B2(n_30),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_95),
.B1(n_66),
.B2(n_60),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_92),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_55),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_24),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_66),
.B1(n_73),
.B2(n_69),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_55),
.A2(n_33),
.B1(n_17),
.B2(n_5),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_96),
.A2(n_97),
.B(n_99),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_106),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_55),
.B1(n_53),
.B2(n_57),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_110),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_53),
.B1(n_57),
.B2(n_56),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_84),
.A2(n_53),
.B1(n_56),
.B2(n_62),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_83),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_90),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_125),
.Y(n_128)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_78),
.C(n_81),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_124),
.C(n_79),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_127),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_78),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

INVx6_ASAP7_75t_SL g127 ( 
.A(n_102),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_127),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_129),
.B(n_131),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_116),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_132),
.B(n_139),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_120),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_134),
.A2(n_120),
.B(n_119),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_123),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_79),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_113),
.C(n_107),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_141),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_102),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_104),
.B(n_118),
.Y(n_155)
);

OAI32xp33_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_107),
.A3(n_119),
.B1(n_111),
.B2(n_110),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_148),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_120),
.B1(n_101),
.B2(n_112),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_147),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_133),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_139),
.B(n_103),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_149),
.B(n_117),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_101),
.B1(n_137),
.B2(n_130),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_155),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_132),
.C(n_136),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_98),
.C(n_99),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_143),
.A2(n_135),
.B(n_138),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_153),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_SL g154 ( 
.A1(n_148),
.A2(n_138),
.B(n_121),
.Y(n_154)
);

OAI322xp33_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_97),
.A3(n_89),
.B1(n_77),
.B2(n_80),
.C1(n_69),
.C2(n_76),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_3),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_164),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_158),
.A2(n_140),
.B1(n_146),
.B2(n_145),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_4),
.C(n_6),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_166),
.C(n_155),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_163),
.A2(n_82),
.B1(n_7),
.B2(n_8),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_13),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_11),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_91),
.C(n_76),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_171),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_166),
.A2(n_64),
.B(n_82),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_169),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_15),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_175),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_170),
.A2(n_159),
.B1(n_162),
.B2(n_14),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_177),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_174),
.A2(n_15),
.B(n_7),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_178),
.A2(n_6),
.B(n_8),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_173),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_182),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_179),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_183),
.B(n_6),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_184),
.Y(n_186)
);


endmodule