module real_jpeg_6176_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_1),
.B(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_1),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_2),
.B(n_34),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_2),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_2),
.B(n_60),
.Y(n_149)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_3),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_3),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_3),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_3),
.B(n_218),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_3),
.B(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_4),
.Y(n_216)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_4),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_5),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_5),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_5),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_5),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_5),
.B(n_47),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_6),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_6),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_6),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_6),
.B(n_134),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_6),
.B(n_227),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_6),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_6),
.B(n_274),
.Y(n_273)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_8),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_8),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_8),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_8),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_8),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_8),
.B(n_243),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_8),
.B(n_276),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_9),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_9),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_9),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_10),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_10),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_10),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_10),
.B(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_11),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_11),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_11),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_11),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_11),
.B(n_45),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_11),
.B(n_134),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_12),
.Y(n_77)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_13),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_14),
.B(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_15),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_15),
.Y(n_117)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_15),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_16),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_16),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_16),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_16),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_16),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_16),
.B(n_213),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_16),
.B(n_250),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_16),
.B(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_17),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_188),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_187),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_157),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_22),
.B(n_157),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_98),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_63),
.C(n_78),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_24),
.B(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_40),
.C(n_48),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_25),
.A2(n_26),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_31),
.Y(n_26)
);

MAJx2_ASAP7_75t_L g143 ( 
.A(n_27),
.B(n_32),
.C(n_39),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_28),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_30),
.B(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_37),
.B2(n_39),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_36),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_36),
.Y(n_198)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_38),
.Y(n_108)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_41),
.B(n_49),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_46),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_42),
.B(n_46),
.Y(n_291)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJx2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_54),
.C(n_59),
.Y(n_49)
);

FAx1_ASAP7_75t_SL g288 ( 
.A(n_50),
.B(n_54),
.CI(n_59),
.CON(n_288),
.SN(n_288)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_53),
.Y(n_277)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_57),
.Y(n_243)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_58),
.Y(n_228)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_58),
.Y(n_271)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_61),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_63),
.B(n_78),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_64),
.B(n_69),
.C(n_74),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_74),
.Y(n_68)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_72),
.Y(n_248)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_77),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_87),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

MAJx2_ASAP7_75t_L g145 ( 
.A(n_80),
.B(n_83),
.C(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_82),
.Y(n_261)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_86),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_87),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.C(n_94),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_88),
.B(n_182),
.Y(n_181)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_91),
.A2(n_94),
.B1(n_95),
.B2(n_183),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_91),
.Y(n_183)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_93),
.Y(n_224)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_93),
.Y(n_250)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_125),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_109),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.Y(n_103)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_121),
.B1(n_122),
.B2(n_124),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_119),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_144),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_136),
.C(n_143),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_127),
.A2(n_128),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_132),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_133),
.C(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_136),
.A2(n_137),
.B(n_139),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_136),
.B(n_143),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_138),
.Y(n_201)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_138),
.Y(n_219)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_147),
.B1(n_155),
.B2(n_156),
.Y(n_144)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_153),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.C(n_184),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_159),
.B(n_311),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_161),
.B(n_184),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_179),
.C(n_180),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_162),
.B(n_304),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_168),
.C(n_174),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_163),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_262)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_169),
.B(n_175),
.Y(n_285)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_173),
.Y(n_274)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_179),
.Y(n_305)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_185),
.Y(n_186)
);

AOI21x1_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_309),
.B(n_313),
.Y(n_188)
);

OAI21x1_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_296),
.B(n_308),
.Y(n_189)
);

AOI21x1_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_281),
.B(n_295),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_253),
.B(n_280),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_230),
.B(n_252),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_207),
.B(n_229),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_204),
.B(n_206),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_202),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_202),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_199),
.Y(n_208)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_209),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_220),
.B2(n_221),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_210),
.B(n_223),
.C(n_225),
.Y(n_251)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_217),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_217),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_225),
.B2(n_226),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_251),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_251),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_241),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_240),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_240),
.C(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_239),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_239),
.Y(n_258)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_265),
.C(n_266),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_249),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_249),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_256),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_263),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_257),
.B(n_264),
.C(n_267),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_260),
.C(n_262),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_267),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_272),
.Y(n_267)
);

MAJx2_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_275),
.C(n_278),
.Y(n_293)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_275),
.B1(n_278),
.B2(n_279),
.Y(n_272)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_273),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_275),
.Y(n_279)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_294),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_294),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_287),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_286),
.C(n_307),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_291),
.C(n_292),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g315 ( 
.A(n_288),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_293),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_306),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_306),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_303),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_300),
.C(n_303),
.Y(n_312)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_312),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_312),
.Y(n_313)
);


endmodule