module fake_jpeg_15492_n_277 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_277);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_175;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_258;
wire n_96;

INVx4_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_3),
.B(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_7),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_40),
.B(n_44),
.Y(n_101)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_19),
.A2(n_0),
.B(n_1),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_58),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_1),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_1),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_3),
.Y(n_49)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_26),
.B(n_31),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_56),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_34),
.Y(n_55)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_29),
.B(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_5),
.C(n_6),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_21),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_37),
.Y(n_105)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_75),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_72),
.B(n_74),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_29),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_66),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_78),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_40),
.B(n_17),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_17),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_85),
.Y(n_118)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_42),
.A2(n_24),
.B1(n_32),
.B2(n_16),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_88),
.A2(n_21),
.B1(n_28),
.B2(n_59),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_39),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_90),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_39),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_91),
.Y(n_144)
);

CKINVDCx6p67_ASAP7_75t_R g95 ( 
.A(n_50),
.Y(n_95)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_54),
.A2(n_36),
.B1(n_24),
.B2(n_38),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_99),
.A2(n_102),
.B1(n_65),
.B2(n_30),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_48),
.A2(n_63),
.B1(n_38),
.B2(n_25),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_52),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_103),
.B(n_30),
.Y(n_110)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_27),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_41),
.A2(n_32),
.B1(n_37),
.B2(n_30),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_133)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_117),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_79),
.A2(n_101),
.B(n_67),
.C(n_69),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_113),
.B(n_137),
.Y(n_150)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_115),
.Y(n_174)
);

INVx4_ASAP7_75t_SL g116 ( 
.A(n_76),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_116),
.Y(n_164)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_119),
.A2(n_131),
.B(n_133),
.Y(n_168)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_130),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_57),
.C(n_33),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_132),
.C(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_123),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_129),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_83),
.B(n_5),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_68),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_82),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_98),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_92),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_33),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_133),
.A2(n_68),
.B1(n_87),
.B2(n_80),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_73),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_145),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_27),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_138),
.Y(n_147)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_8),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_139),
.A2(n_114),
.B(n_144),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_95),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_71),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_140),
.B(n_109),
.C(n_123),
.Y(n_167)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_108),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_98),
.B(n_14),
.C(n_82),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_140),
.Y(n_172)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_122),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_148),
.B(n_176),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_149),
.A2(n_154),
.B1(n_129),
.B2(n_112),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_95),
.B(n_80),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_153),
.A2(n_157),
.B(n_163),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_155),
.B(n_158),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_124),
.B(n_100),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_160),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_137),
.A2(n_85),
.B(n_98),
.Y(n_157)
);

FAx1_ASAP7_75t_SL g158 ( 
.A(n_118),
.B(n_70),
.CI(n_104),
.CON(n_158),
.SN(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_96),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_113),
.B(n_70),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_162),
.Y(n_189)
);

NOR3xp33_ASAP7_75t_SL g203 ( 
.A(n_167),
.B(n_171),
.C(n_177),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_135),
.Y(n_169)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_115),
.A2(n_126),
.B1(n_136),
.B2(n_138),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_170),
.A2(n_174),
.B1(n_155),
.B2(n_156),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g171 ( 
.A(n_111),
.B(n_139),
.C(n_130),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_141),
.C(n_120),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_117),
.B(n_139),
.Y(n_173)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_140),
.B(n_143),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_125),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_178),
.A2(n_200),
.B1(n_174),
.B2(n_168),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_180),
.B(n_172),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_195),
.Y(n_206)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_159),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_186),
.B(n_198),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_128),
.C(n_145),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_192),
.C(n_193),
.Y(n_216)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_128),
.C(n_116),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_125),
.C(n_112),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_158),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_162),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_199),
.Y(n_212)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_202),
.Y(n_221)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_146),
.Y(n_202)
);

AO21x1_ASAP7_75t_L g210 ( 
.A1(n_203),
.A2(n_150),
.B(n_173),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_194),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_213),
.Y(n_227)
);

A2O1A1O1Ixp25_ASAP7_75t_L g205 ( 
.A1(n_203),
.A2(n_185),
.B(n_167),
.C(n_190),
.D(n_153),
.Y(n_205)
);

AOI21xp33_ASAP7_75t_L g239 ( 
.A1(n_205),
.A2(n_210),
.B(n_179),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_208),
.B(n_181),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_195),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_220),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_154),
.B1(n_161),
.B2(n_160),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_218),
.B1(n_223),
.B2(n_224),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_183),
.A2(n_154),
.B1(n_170),
.B2(n_149),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_190),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_191),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_157),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_225),
.C(n_180),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_178),
.A2(n_150),
.B1(n_158),
.B2(n_146),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_188),
.A2(n_148),
.B1(n_164),
.B2(n_175),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_163),
.C(n_164),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_228),
.C(n_236),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_192),
.C(n_193),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

BUFx12_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_230),
.B(n_238),
.Y(n_242)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_240),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_215),
.A2(n_189),
.B(n_196),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_233),
.A2(n_209),
.B(n_217),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_237),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_181),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_218),
.A2(n_188),
.B1(n_189),
.B2(n_200),
.Y(n_238)
);

A2O1A1O1Ixp25_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_219),
.B(n_225),
.C(n_224),
.D(n_182),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_212),
.B(n_199),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_220),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_243),
.Y(n_256)
);

AOI322xp5_ASAP7_75t_L g245 ( 
.A1(n_234),
.A2(n_231),
.A3(n_205),
.B1(n_235),
.B2(n_233),
.C1(n_210),
.C2(n_238),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_247),
.Y(n_257)
);

AO21x1_ASAP7_75t_L g261 ( 
.A1(n_246),
.A2(n_232),
.B(n_241),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_216),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_222),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_226),
.C(n_228),
.Y(n_255)
);

AOI31xp67_ASAP7_75t_L g260 ( 
.A1(n_250),
.A2(n_206),
.A3(n_211),
.B(n_230),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_243),
.A2(n_231),
.B(n_227),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_253),
.A2(n_242),
.B(n_250),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_244),
.B(n_217),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_254),
.B(n_259),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_255),
.A2(n_260),
.B(n_248),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_251),
.B(n_211),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_258),
.B(n_261),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_230),
.Y(n_259)
);

AOI322xp5_ASAP7_75t_L g271 ( 
.A1(n_262),
.A2(n_263),
.A3(n_267),
.B1(n_248),
.B2(n_252),
.C1(n_147),
.C2(n_184),
.Y(n_271)
);

BUFx24_ASAP7_75t_SL g264 ( 
.A(n_257),
.Y(n_264)
);

BUFx24_ASAP7_75t_SL g270 ( 
.A(n_264),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_255),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_256),
.Y(n_268)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_268),
.Y(n_273)
);

NAND4xp25_ASAP7_75t_SL g269 ( 
.A(n_265),
.B(n_261),
.C(n_256),
.D(n_147),
.Y(n_269)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_269),
.Y(n_274)
);

NAND3xp33_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_252),
.C(n_147),
.Y(n_272)
);

AO21x1_ASAP7_75t_L g275 ( 
.A1(n_272),
.A2(n_270),
.B(n_162),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_276),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_274),
.Y(n_276)
);


endmodule