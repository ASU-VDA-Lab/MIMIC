module real_jpeg_22085_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

OAI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_0),
.A2(n_32),
.B1(n_38),
.B2(n_39),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_0),
.A2(n_32),
.B1(n_58),
.B2(n_59),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_0),
.A2(n_32),
.B1(n_53),
.B2(n_54),
.Y(n_105)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_3),
.B(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_3),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_3),
.B(n_31),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_3),
.B(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_5),
.A2(n_53),
.B1(n_54),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_5),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_5),
.A2(n_58),
.B1(n_59),
.B2(n_67),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_67),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_67),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_6),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_42),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_8),
.A2(n_53),
.B(n_55),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_8),
.B(n_53),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_8),
.A2(n_26),
.B1(n_58),
.B2(n_59),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_8),
.A2(n_26),
.B1(n_38),
.B2(n_39),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_8),
.B(n_56),
.Y(n_162)
);

AOI21xp33_ASAP7_75t_L g179 ( 
.A1(n_8),
.A2(n_10),
.B(n_25),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_8),
.B(n_125),
.Y(n_200)
);

O2A1O1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_8),
.A2(n_58),
.B(n_73),
.C(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_9),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_57)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_9),
.A2(n_53),
.B(n_57),
.C(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_9),
.B(n_53),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_10),
.Y(n_36)
);

O2A1O1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_10),
.A2(n_35),
.B(n_38),
.C(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_10),
.B(n_38),
.Y(n_46)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_11),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_136),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_134),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_106),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_15),
.B(n_106),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_91),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_82),
.B2(n_83),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_47),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_33),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_20),
.B(n_33),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_21),
.B(n_188),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_22),
.B(n_28),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_23),
.A2(n_29),
.B(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_24),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_30),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_26),
.A2(n_36),
.B(n_39),
.C(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_26),
.B(n_34),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_26),
.B(n_86),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_L g211 ( 
.A1(n_26),
.A2(n_38),
.B(n_75),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_27),
.A2(n_30),
.B(n_94),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_27),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_28),
.B(n_175),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_29),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.B(n_43),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_34),
.A2(n_88),
.B(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_35),
.B(n_44),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_35),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_35),
.B(n_98),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_37),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_38),
.A2(n_39),
.B1(n_73),
.B2(n_75),
.Y(n_72)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_43),
.B(n_182),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_45),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_45),
.B(n_183),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_68),
.B2(n_81),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_61),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_56),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_52),
.B(n_63),
.Y(n_143)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_56),
.B(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_66),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_72),
.B(n_73),
.C(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_73),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_58),
.B(n_60),
.Y(n_119)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_59),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_61),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_105),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_76),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_70),
.B(n_127),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_71),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_72),
.A2(n_79),
.B(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_76),
.B(n_149),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_77),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_77),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_78),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_79),
.B(n_128),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_87),
.B2(n_90),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_84),
.A2(n_85),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_85),
.B(n_210),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_87),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_89),
.B(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_99),
.C(n_102),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_96),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_95),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_95),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_97),
.B(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_99),
.A2(n_100),
.B1(n_102),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.C(n_111),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_107),
.B(n_110),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_111),
.A2(n_112),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_122),
.C(n_130),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_113),
.A2(n_114),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_122),
.A2(n_123),
.B1(n_130),
.B2(n_131),
.Y(n_153)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_129),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_166),
.B(n_243),
.C(n_248),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_155),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_138),
.B(n_155),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_152),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_140),
.B(n_141),
.C(n_152),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.C(n_147),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_159),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_156),
.B(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_158),
.Y(n_240)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.C(n_163),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_161),
.B(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_162),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_174),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_242),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_236),
.B(n_241),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_221),
.B(n_235),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_206),
.B(n_220),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_195),
.B(n_205),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_184),
.B(n_194),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_176),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_178),
.B(n_180),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_189),
.B(n_193),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_187),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_197),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_204),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_202),
.C(n_204),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_208),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_213),
.B1(n_214),
.B2(n_219),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_209),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_210),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_215),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_218),
.C(n_219),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_222),
.B(n_223),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_228),
.B2(n_229),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_230),
.C(n_234),
.Y(n_237)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_230),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_232),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_237),
.B(n_238),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_244),
.B(n_245),
.Y(n_248)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);


endmodule