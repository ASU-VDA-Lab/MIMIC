module fake_netlist_6_1016_n_2062 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2062);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2062;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_405;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_1094;
wire n_953;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_811;
wire n_683;
wire n_527;
wire n_474;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g217 ( 
.A(n_64),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_90),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_87),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_177),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_216),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_154),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_93),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_98),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_180),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_163),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_84),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_156),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_173),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_186),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_126),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_147),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_134),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_151),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_205),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_38),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_111),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_46),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_12),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_189),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_77),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_179),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_165),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_85),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_32),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_164),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_124),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_97),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_51),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_178),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_181),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_168),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_100),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_182),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_116),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_210),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_36),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_45),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_75),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_56),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_24),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_209),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_136),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_196),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_198),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_174),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_121),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_148),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_204),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_137),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_203),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_47),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_20),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_128),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_105),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_10),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_78),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_91),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_32),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_120),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_28),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_96),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_14),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_59),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_46),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_11),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_117),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_150),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_58),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_153),
.Y(n_293)
);

BUFx10_ASAP7_75t_L g294 ( 
.A(n_26),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_94),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_73),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_40),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_34),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_56),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_5),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_61),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_6),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_79),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_62),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_88),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_13),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_3),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_25),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_48),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_59),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_17),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_57),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_51),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_7),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_24),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_99),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_43),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_72),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_135),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_81),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_12),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_187),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_161),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_143),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_206),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_155),
.Y(n_326)
);

BUFx5_ASAP7_75t_L g327 ( 
.A(n_197),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_140),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_60),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_6),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_172),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_130),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_101),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_144),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_138),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_125),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_67),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_191),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_8),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_157),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_76),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_167),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_74),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_119),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_53),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_112),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_36),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_60),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_40),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_170),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_45),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_29),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_113),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_141),
.Y(n_354)
);

BUFx8_ASAP7_75t_SL g355 ( 
.A(n_190),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_110),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_11),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_1),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_127),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_21),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_18),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_31),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_89),
.Y(n_363)
);

INVxp33_ASAP7_75t_L g364 ( 
.A(n_65),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_28),
.Y(n_365)
);

BUFx2_ASAP7_75t_SL g366 ( 
.A(n_49),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_42),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_44),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_103),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_21),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_146),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_131),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_129),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_58),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_15),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_194),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_65),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_159),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_16),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_122),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_118),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_4),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_53),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_42),
.Y(n_384)
);

BUFx5_ASAP7_75t_L g385 ( 
.A(n_64),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_31),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g387 ( 
.A(n_66),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_176),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_35),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_30),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_67),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_215),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_44),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_71),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_5),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_8),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_109),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_213),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_192),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_86),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_62),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_175),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_39),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_2),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_27),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_43),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_49),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_19),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_171),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_37),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_30),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_16),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_184),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_142),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_188),
.Y(n_415)
);

BUFx8_ASAP7_75t_SL g416 ( 
.A(n_114),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_17),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_29),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_95),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_7),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_106),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_166),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_199),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_195),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_0),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_15),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_149),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_139),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_169),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_80),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_385),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_302),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_271),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_355),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_385),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_385),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_352),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_385),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_385),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_386),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_416),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_385),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_257),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_368),
.Y(n_444)
);

INVxp33_ASAP7_75t_SL g445 ( 
.A(n_242),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_258),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_385),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_426),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_259),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_267),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_249),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_385),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_285),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_268),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_312),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_269),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_312),
.Y(n_457)
);

INVxp33_ASAP7_75t_SL g458 ( 
.A(n_242),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_312),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_272),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_274),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_294),
.Y(n_462)
);

INVxp33_ASAP7_75t_SL g463 ( 
.A(n_248),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_294),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_312),
.Y(n_465)
);

INVxp67_ASAP7_75t_SL g466 ( 
.A(n_415),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_312),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_314),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_314),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_280),
.Y(n_470)
);

INVxp67_ASAP7_75t_SL g471 ( 
.A(n_220),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_277),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_293),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_370),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_226),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_370),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_384),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_384),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_412),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_327),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_281),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_226),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_412),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_337),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_337),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_367),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_367),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_356),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_375),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_375),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_217),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_327),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_241),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_252),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_264),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_286),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_296),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_327),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_311),
.Y(n_499)
);

INVxp67_ASAP7_75t_SL g500 ( 
.A(n_429),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_283),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_290),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_327),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_291),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_315),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_327),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_248),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_329),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_305),
.Y(n_509)
);

INVxp67_ASAP7_75t_SL g510 ( 
.A(n_429),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g511 ( 
.A(n_266),
.Y(n_511)
);

INVxp67_ASAP7_75t_SL g512 ( 
.A(n_218),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_402),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_224),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_327),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_294),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_339),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_327),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_360),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_319),
.Y(n_520)
);

INVxp33_ASAP7_75t_SL g521 ( 
.A(n_401),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_327),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_365),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_374),
.Y(n_524)
);

INVxp33_ASAP7_75t_SL g525 ( 
.A(n_401),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_379),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_391),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_393),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_408),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_425),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_403),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_325),
.Y(n_532)
);

INVxp33_ASAP7_75t_L g533 ( 
.A(n_364),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_238),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_232),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_238),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_276),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_276),
.Y(n_538)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_306),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_233),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_387),
.Y(n_541)
);

INVxp33_ASAP7_75t_L g542 ( 
.A(n_235),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_320),
.Y(n_543)
);

INVxp67_ASAP7_75t_SL g544 ( 
.A(n_239),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_323),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_387),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_326),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_431),
.A2(n_397),
.B(n_245),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_455),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_455),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_457),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_457),
.Y(n_552)
);

AND2x4_ASAP7_75t_L g553 ( 
.A(n_512),
.B(n_254),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_459),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_459),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_465),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_465),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_467),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_467),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_431),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_435),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_435),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_436),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_436),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_443),
.B(n_446),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_544),
.B(n_245),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_475),
.B(n_318),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_438),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_449),
.B(n_397),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_438),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_482),
.B(n_236),
.Y(n_571)
);

INVxp67_ASAP7_75t_SL g572 ( 
.A(n_500),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_450),
.B(n_278),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_439),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_454),
.B(n_244),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_439),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_442),
.Y(n_577)
);

OAI21x1_ASAP7_75t_L g578 ( 
.A1(n_442),
.A2(n_251),
.B(n_250),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_447),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_456),
.B(n_262),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_514),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_514),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_447),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_452),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_452),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_480),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_480),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_492),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_SL g589 ( 
.A(n_511),
.B(n_378),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_524),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_524),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_492),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_530),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_498),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_498),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_503),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_507),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_503),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_530),
.Y(n_599)
);

NOR2xp67_ASAP7_75t_L g600 ( 
.A(n_506),
.B(n_270),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_491),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_506),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_515),
.Y(n_603)
);

CKINVDCx16_ASAP7_75t_R g604 ( 
.A(n_440),
.Y(n_604)
);

AND2x2_ASAP7_75t_SL g605 ( 
.A(n_511),
.B(n_228),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_515),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_491),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_518),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_493),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_510),
.B(n_219),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_518),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_533),
.B(n_219),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_460),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_493),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_522),
.Y(n_615)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_531),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_461),
.B(n_273),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_494),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_522),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_535),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_494),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_470),
.B(n_295),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_495),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_495),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_496),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_468),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_L g627 ( 
.A(n_481),
.B(n_403),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_501),
.B(n_303),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_468),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_532),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_433),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_496),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_469),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_535),
.Y(n_634)
);

NOR3xp33_ASAP7_75t_L g635 ( 
.A(n_440),
.B(n_420),
.C(n_288),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_432),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_469),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_540),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_484),
.B(n_221),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_497),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_497),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_587),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_554),
.Y(n_643)
);

NOR2x1p5_ASAP7_75t_L g644 ( 
.A(n_613),
.B(n_434),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_587),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_563),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_556),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_605),
.A2(n_471),
.B1(n_472),
.B2(n_543),
.Y(n_648)
);

INVx4_ASAP7_75t_L g649 ( 
.A(n_563),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_556),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_592),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_561),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_572),
.B(n_502),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_563),
.Y(n_654)
);

NOR3xp33_ASAP7_75t_L g655 ( 
.A(n_604),
.B(n_437),
.C(n_451),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_581),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_587),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_610),
.Y(n_658)
);

AND3x2_ASAP7_75t_L g659 ( 
.A(n_589),
.B(n_432),
.C(n_462),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_581),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_610),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_561),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_587),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_592),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_587),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_631),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_605),
.B(n_504),
.Y(n_667)
);

AND3x2_ASAP7_75t_L g668 ( 
.A(n_573),
.B(n_516),
.C(n_464),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_605),
.B(n_509),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_562),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_592),
.Y(n_671)
);

NAND2xp33_ASAP7_75t_L g672 ( 
.A(n_569),
.B(n_228),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_639),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_562),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_594),
.Y(n_675)
);

INVxp33_ASAP7_75t_L g676 ( 
.A(n_612),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_564),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_594),
.Y(n_678)
);

AND2x6_ASAP7_75t_L g679 ( 
.A(n_553),
.B(n_228),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_587),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_594),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_602),
.Y(n_682)
);

AOI21x1_ASAP7_75t_L g683 ( 
.A1(n_600),
.A2(n_322),
.B(n_316),
.Y(n_683)
);

INVx5_ASAP7_75t_L g684 ( 
.A(n_563),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_564),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_588),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_639),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_602),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_602),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_627),
.A2(n_545),
.B1(n_466),
.B2(n_520),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_568),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_588),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_571),
.Y(n_693)
);

AO22x2_ASAP7_75t_L g694 ( 
.A1(n_636),
.A2(n_444),
.B1(n_366),
.B2(n_448),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_571),
.Y(n_695)
);

OAI22xp33_ASAP7_75t_L g696 ( 
.A1(n_636),
.A2(n_542),
.B1(n_263),
.B2(n_275),
.Y(n_696)
);

INVxp67_ASAP7_75t_SL g697 ( 
.A(n_620),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_606),
.Y(n_698)
);

AND2x2_ASAP7_75t_SL g699 ( 
.A(n_553),
.B(n_228),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_606),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_606),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_553),
.B(n_547),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_575),
.B(n_445),
.Y(n_703)
);

INVx6_ASAP7_75t_L g704 ( 
.A(n_620),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_581),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_553),
.B(n_540),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_568),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_588),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_611),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_574),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_611),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_574),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_582),
.Y(n_713)
);

BUFx16f_ASAP7_75t_R g714 ( 
.A(n_604),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_L g715 ( 
.A(n_580),
.B(n_228),
.Y(n_715)
);

AO22x1_ASAP7_75t_L g716 ( 
.A1(n_635),
.A2(n_405),
.B1(n_406),
.B2(n_404),
.Y(n_716)
);

INVx5_ASAP7_75t_L g717 ( 
.A(n_563),
.Y(n_717)
);

BUFx10_ASAP7_75t_L g718 ( 
.A(n_566),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_582),
.B(n_620),
.Y(n_719)
);

OA22x2_ASAP7_75t_L g720 ( 
.A1(n_567),
.A2(n_536),
.B1(n_537),
.B2(n_534),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_560),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_617),
.B(n_328),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_567),
.B(n_484),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_579),
.Y(n_724)
);

AO22x2_ASAP7_75t_L g725 ( 
.A1(n_597),
.A2(n_333),
.B1(n_338),
.B2(n_334),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_588),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_566),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_560),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_579),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_585),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_622),
.B(n_336),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_585),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_628),
.B(n_620),
.Y(n_733)
);

CKINVDCx20_ASAP7_75t_R g734 ( 
.A(n_630),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_566),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_588),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_620),
.B(n_340),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_620),
.B(n_341),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_560),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_570),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_583),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_634),
.B(n_499),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_588),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_583),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_595),
.Y(n_745)
);

OR2x6_ASAP7_75t_L g746 ( 
.A(n_565),
.B(n_485),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_570),
.Y(n_747)
);

INVx4_ASAP7_75t_L g748 ( 
.A(n_563),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_634),
.B(n_458),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_570),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_630),
.Y(n_751)
);

INVx5_ASAP7_75t_L g752 ( 
.A(n_576),
.Y(n_752)
);

INVxp33_ASAP7_75t_L g753 ( 
.A(n_601),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_616),
.A2(n_521),
.B1(n_525),
.B2(n_463),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_577),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_634),
.B(n_441),
.Y(n_756)
);

NAND2xp33_ASAP7_75t_L g757 ( 
.A(n_576),
.B(n_265),
.Y(n_757)
);

OR2x6_ASAP7_75t_L g758 ( 
.A(n_566),
.B(n_485),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_634),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_577),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_634),
.B(n_539),
.Y(n_761)
);

AOI21x1_ASAP7_75t_L g762 ( 
.A1(n_600),
.A2(n_548),
.B(n_577),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_634),
.B(n_638),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_638),
.B(n_499),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_638),
.B(n_343),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_584),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_601),
.B(n_486),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_584),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_584),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_638),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_550),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_638),
.B(n_221),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_638),
.B(n_222),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_548),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_576),
.B(n_344),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_550),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_595),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_576),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_551),
.Y(n_779)
);

NAND3xp33_ASAP7_75t_L g780 ( 
.A(n_607),
.B(n_487),
.C(n_486),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_607),
.B(n_487),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_576),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_576),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_595),
.B(n_346),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_595),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_552),
.Y(n_786)
);

NAND2xp33_ASAP7_75t_L g787 ( 
.A(n_595),
.B(n_265),
.Y(n_787)
);

INVx4_ASAP7_75t_L g788 ( 
.A(n_595),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_596),
.B(n_350),
.Y(n_789)
);

NOR2x1p5_ASAP7_75t_L g790 ( 
.A(n_609),
.B(n_404),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_609),
.B(n_222),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_552),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_555),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_555),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_614),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_614),
.B(n_223),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_596),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_557),
.Y(n_798)
);

NOR3xp33_ASAP7_75t_L g799 ( 
.A(n_667),
.B(n_490),
.C(n_489),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_719),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_719),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_727),
.B(n_596),
.Y(n_802)
);

INVxp33_ASAP7_75t_L g803 ( 
.A(n_754),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_699),
.A2(n_578),
.B1(n_261),
.B2(n_299),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_790),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_651),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_693),
.B(n_223),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_735),
.B(n_699),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_693),
.B(n_225),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_695),
.B(n_658),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_735),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_695),
.B(n_225),
.Y(n_812)
);

NAND3xp33_ASAP7_75t_L g813 ( 
.A(n_658),
.B(n_661),
.C(n_648),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_661),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_673),
.B(n_596),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_702),
.B(n_227),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_795),
.B(n_489),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_767),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_673),
.B(n_596),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_767),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_781),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_687),
.B(n_227),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_718),
.B(n_265),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_664),
.Y(n_824)
);

O2A1O1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_687),
.A2(n_618),
.B(n_623),
.C(n_621),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_781),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_771),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_652),
.B(n_596),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_652),
.B(n_598),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_718),
.B(n_229),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_753),
.B(n_229),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_670),
.B(n_598),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_670),
.B(n_598),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_758),
.Y(n_834)
);

NAND2xp33_ASAP7_75t_L g835 ( 
.A(n_679),
.B(n_353),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_718),
.B(n_265),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_671),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_792),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_674),
.B(n_677),
.Y(n_839)
);

INVx6_ASAP7_75t_L g840 ( 
.A(n_719),
.Y(n_840)
);

NAND2xp33_ASAP7_75t_L g841 ( 
.A(n_679),
.B(n_354),
.Y(n_841)
);

OR2x2_ASAP7_75t_L g842 ( 
.A(n_746),
.B(n_490),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_674),
.B(n_598),
.Y(n_843)
);

OR2x2_ASAP7_75t_L g844 ( 
.A(n_746),
.B(n_641),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_653),
.B(n_230),
.Y(n_845)
);

BUFx5_ASAP7_75t_L g846 ( 
.A(n_774),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_656),
.B(n_231),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_792),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_677),
.B(n_685),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_723),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_734),
.Y(n_851)
);

NAND2xp33_ASAP7_75t_L g852 ( 
.A(n_679),
.B(n_363),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_675),
.Y(n_853)
);

AO22x1_ASAP7_75t_L g854 ( 
.A1(n_676),
.A2(n_406),
.B1(n_410),
.B2(n_405),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_675),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_710),
.B(n_598),
.Y(n_856)
);

OAI221xp5_ASAP7_75t_L g857 ( 
.A1(n_706),
.A2(n_641),
.B1(n_640),
.B2(n_618),
.C(n_632),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_712),
.B(n_598),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_656),
.B(n_231),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_733),
.B(n_265),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_703),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_774),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_669),
.B(n_234),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_723),
.A2(n_578),
.B1(n_307),
.B2(n_308),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_725),
.A2(n_321),
.B1(n_351),
.B2(n_282),
.Y(n_865)
);

OAI22xp33_ASAP7_75t_L g866 ( 
.A1(n_758),
.A2(n_746),
.B1(n_720),
.B2(n_690),
.Y(n_866)
);

O2A1O1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_712),
.A2(n_623),
.B(n_624),
.C(n_621),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_724),
.B(n_608),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_784),
.A2(n_615),
.B(n_608),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_724),
.B(n_608),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_729),
.B(n_608),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_729),
.B(n_730),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_SL g873 ( 
.A1(n_694),
.A2(n_473),
.B1(n_488),
.B2(n_453),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_730),
.B(n_732),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_732),
.B(n_608),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_662),
.B(n_324),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_691),
.B(n_608),
.Y(n_877)
);

INVx8_ASAP7_75t_L g878 ( 
.A(n_746),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_678),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_707),
.B(n_324),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_722),
.B(n_731),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_678),
.Y(n_882)
);

OR2x2_ASAP7_75t_L g883 ( 
.A(n_758),
.B(n_640),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_713),
.B(n_615),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_681),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_758),
.B(n_624),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_713),
.B(n_615),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_660),
.B(n_513),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_742),
.B(n_615),
.Y(n_889)
);

OAI21xp33_ASAP7_75t_L g890 ( 
.A1(n_720),
.A2(n_536),
.B(n_534),
.Y(n_890)
);

INVxp67_ASAP7_75t_L g891 ( 
.A(n_791),
.Y(n_891)
);

OAI221xp5_ASAP7_75t_L g892 ( 
.A1(n_720),
.A2(n_625),
.B1(n_632),
.B2(n_359),
.C(n_373),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_759),
.B(n_324),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_759),
.B(n_324),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_666),
.Y(n_895)
);

AND2x6_ASAP7_75t_SL g896 ( 
.A(n_714),
.B(n_505),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_764),
.B(n_615),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_764),
.B(n_615),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_660),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_679),
.B(n_776),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_776),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_679),
.B(n_619),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_679),
.B(n_619),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_779),
.B(n_619),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_770),
.Y(n_905)
);

AND2x2_ASAP7_75t_SL g906 ( 
.A(n_715),
.B(n_324),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_779),
.B(n_619),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_786),
.Y(n_908)
);

O2A1O1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_672),
.A2(n_625),
.B(n_558),
.C(n_559),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_705),
.A2(n_371),
.B1(n_398),
.B2(n_381),
.Y(n_910)
);

OAI221xp5_ASAP7_75t_L g911 ( 
.A1(n_780),
.A2(n_342),
.B1(n_388),
.B2(n_414),
.C(n_430),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_786),
.B(n_619),
.Y(n_912)
);

OA21x2_ASAP7_75t_L g913 ( 
.A1(n_762),
.A2(n_558),
.B(n_557),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_705),
.B(n_331),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_793),
.B(n_619),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_794),
.B(n_586),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_794),
.B(n_586),
.Y(n_917)
);

AND2x2_ASAP7_75t_SL g918 ( 
.A(n_715),
.B(n_672),
.Y(n_918)
);

NAND2x1p5_ASAP7_75t_L g919 ( 
.A(n_770),
.B(n_331),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_798),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_798),
.B(n_586),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_749),
.A2(n_369),
.B1(n_372),
.B2(n_376),
.Y(n_922)
);

INVxp67_ASAP7_75t_L g923 ( 
.A(n_796),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_741),
.B(n_603),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_682),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_696),
.B(n_234),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_761),
.B(n_237),
.Y(n_927)
);

INVxp67_ASAP7_75t_L g928 ( 
.A(n_694),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_688),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_744),
.B(n_603),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_775),
.B(n_603),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_642),
.B(n_603),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_642),
.B(n_559),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_642),
.B(n_626),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_659),
.B(n_237),
.Y(n_935)
);

NOR3xp33_ASAP7_75t_SL g936 ( 
.A(n_751),
.B(n_411),
.C(n_410),
.Y(n_936)
);

NOR3xp33_ASAP7_75t_L g937 ( 
.A(n_716),
.B(n_538),
.C(n_537),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_778),
.B(n_331),
.Y(n_938)
);

OR2x2_ASAP7_75t_L g939 ( 
.A(n_716),
.B(n_538),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_L g940 ( 
.A1(n_725),
.A2(n_382),
.B1(n_417),
.B2(n_361),
.Y(n_940)
);

NOR2xp67_ASAP7_75t_L g941 ( 
.A(n_737),
.B(n_738),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_756),
.B(n_772),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_689),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_773),
.B(n_240),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_698),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_668),
.B(n_240),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_765),
.B(n_243),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_645),
.B(n_626),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_655),
.A2(n_380),
.B1(n_392),
.B2(n_243),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_657),
.B(n_549),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_810),
.B(n_751),
.Y(n_951)
);

AOI22xp33_ASAP7_75t_L g952 ( 
.A1(n_926),
.A2(n_725),
.B1(n_750),
.B2(n_694),
.Y(n_952)
);

AND2x6_ASAP7_75t_SL g953 ( 
.A(n_946),
.B(n_541),
.Y(n_953)
);

OAI21xp33_ASAP7_75t_L g954 ( 
.A1(n_926),
.A2(n_694),
.B(n_725),
.Y(n_954)
);

NAND3xp33_ASAP7_75t_L g955 ( 
.A(n_810),
.B(n_789),
.C(n_768),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_850),
.B(n_666),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_901),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_899),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_881),
.B(n_760),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_908),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_920),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_862),
.Y(n_962)
);

INVx2_ASAP7_75t_SL g963 ( 
.A(n_817),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_839),
.B(n_760),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_827),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_814),
.B(n_763),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_861),
.B(n_734),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_806),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_849),
.B(n_768),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_803),
.B(n_407),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_862),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_899),
.B(n_418),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_838),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_872),
.B(n_721),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_942),
.A2(n_697),
.B1(n_783),
.B2(n_782),
.Y(n_975)
);

NAND2x1p5_ASAP7_75t_L g976 ( 
.A(n_800),
.B(n_646),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_862),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_814),
.B(n_644),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_848),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_862),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_SL g981 ( 
.A1(n_873),
.A2(n_865),
.B1(n_940),
.B2(n_895),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_834),
.B(n_505),
.Y(n_982)
);

BUFx4f_ASAP7_75t_L g983 ( 
.A(n_878),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_804),
.A2(n_411),
.B1(n_279),
.B2(n_284),
.Y(n_984)
);

AOI21x1_ASAP7_75t_L g985 ( 
.A1(n_860),
.A2(n_874),
.B(n_902),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_831),
.B(n_541),
.Y(n_986)
);

AND2x6_ASAP7_75t_SL g987 ( 
.A(n_946),
.B(n_546),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_811),
.B(n_721),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_891),
.B(n_646),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_818),
.B(n_728),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_800),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_800),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_942),
.A2(n_863),
.B1(n_866),
.B2(n_816),
.Y(n_993)
);

AO21x1_ASAP7_75t_L g994 ( 
.A1(n_863),
.A2(n_757),
.B(n_762),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_820),
.B(n_728),
.Y(n_995)
);

INVxp67_ASAP7_75t_L g996 ( 
.A(n_831),
.Y(n_996)
);

NAND3xp33_ASAP7_75t_L g997 ( 
.A(n_813),
.B(n_711),
.C(n_709),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_824),
.Y(n_998)
);

AND3x1_ASAP7_75t_SL g999 ( 
.A(n_911),
.B(n_517),
.C(n_508),
.Y(n_999)
);

INVxp67_ASAP7_75t_SL g1000 ( 
.A(n_800),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_821),
.B(n_739),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_851),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_815),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_804),
.A2(n_711),
.B1(n_709),
.B2(n_766),
.Y(n_1004)
);

NAND2x1p5_ASAP7_75t_L g1005 ( 
.A(n_801),
.B(n_646),
.Y(n_1005)
);

CKINVDCx20_ASAP7_75t_R g1006 ( 
.A(n_888),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_819),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_834),
.B(n_508),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_807),
.B(n_546),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_923),
.B(n_649),
.Y(n_1010)
);

BUFx4f_ASAP7_75t_L g1011 ( 
.A(n_878),
.Y(n_1011)
);

NAND3xp33_ASAP7_75t_SL g1012 ( 
.A(n_865),
.B(n_287),
.C(n_260),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_801),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_R g1014 ( 
.A(n_805),
.B(n_246),
.Y(n_1014)
);

NAND2x1p5_ASAP7_75t_L g1015 ( 
.A(n_801),
.B(n_649),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_864),
.A2(n_301),
.B1(n_300),
.B2(n_298),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_826),
.B(n_739),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_864),
.A2(n_292),
.B1(n_289),
.B2(n_297),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_807),
.B(n_306),
.Y(n_1019)
);

INVx4_ASAP7_75t_L g1020 ( 
.A(n_801),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_896),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_808),
.A2(n_766),
.B1(n_747),
.B2(n_755),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_874),
.B(n_740),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_840),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_816),
.B(n_657),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_840),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_822),
.B(n_306),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_844),
.B(n_883),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_837),
.Y(n_1029)
);

NOR2x1p5_ASAP7_75t_L g1030 ( 
.A(n_842),
.B(n_304),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_846),
.B(n_740),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_828),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_886),
.B(n_517),
.Y(n_1033)
);

INVx4_ASAP7_75t_L g1034 ( 
.A(n_840),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_802),
.A2(n_788),
.B(n_654),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_939),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_829),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_832),
.Y(n_1038)
);

XOR2xp5_ASAP7_75t_L g1039 ( 
.A(n_949),
.B(n_246),
.Y(n_1039)
);

NAND3xp33_ASAP7_75t_SL g1040 ( 
.A(n_940),
.B(n_310),
.C(n_309),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_833),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_905),
.Y(n_1042)
);

INVx5_ASAP7_75t_L g1043 ( 
.A(n_905),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_853),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_846),
.B(n_747),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_846),
.B(n_755),
.Y(n_1046)
);

INVx2_ASAP7_75t_SL g1047 ( 
.A(n_809),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_855),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_843),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_879),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_846),
.B(n_769),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_822),
.B(n_918),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_944),
.A2(n_704),
.B1(n_680),
.B2(n_708),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_856),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_882),
.Y(n_1055)
);

NOR2x1p5_ASAP7_75t_L g1056 ( 
.A(n_854),
.B(n_313),
.Y(n_1056)
);

INVxp67_ASAP7_75t_SL g1057 ( 
.A(n_846),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_812),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_SL g1059 ( 
.A1(n_928),
.A2(n_317),
.B1(n_330),
.B2(n_345),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_858),
.Y(n_1060)
);

INVxp67_ASAP7_75t_SL g1061 ( 
.A(n_846),
.Y(n_1061)
);

AOI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_944),
.A2(n_704),
.B1(n_680),
.B2(n_708),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_889),
.A2(n_788),
.B(n_748),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_885),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_941),
.B(n_698),
.Y(n_1065)
);

NOR2x1_ASAP7_75t_R g1066 ( 
.A(n_847),
.B(n_247),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_868),
.Y(n_1067)
);

OR2x2_ASAP7_75t_SL g1068 ( 
.A(n_936),
.B(n_519),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_927),
.B(n_247),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_878),
.Y(n_1070)
);

NAND2x1p5_ASAP7_75t_L g1071 ( 
.A(n_823),
.B(n_654),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_927),
.B(n_253),
.Y(n_1072)
);

OR2x6_ASAP7_75t_L g1073 ( 
.A(n_825),
.B(n_519),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_870),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_799),
.A2(n_643),
.B1(n_647),
.B2(n_650),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_859),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_871),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_913),
.B(n_700),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_914),
.Y(n_1079)
);

INVxp67_ASAP7_75t_L g1080 ( 
.A(n_935),
.Y(n_1080)
);

NAND2x1p5_ASAP7_75t_L g1081 ( 
.A(n_823),
.B(n_836),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_937),
.B(n_523),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_913),
.B(n_700),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_845),
.B(n_253),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_875),
.Y(n_1085)
);

XNOR2xp5_ASAP7_75t_L g1086 ( 
.A(n_910),
.B(n_255),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_867),
.Y(n_1087)
);

AOI22x1_ASAP7_75t_SL g1088 ( 
.A1(n_935),
.A2(n_347),
.B1(n_348),
.B2(n_349),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_914),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_925),
.Y(n_1090)
);

INVx5_ASAP7_75t_L g1091 ( 
.A(n_929),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_890),
.B(n_523),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_830),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_922),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_900),
.Y(n_1095)
);

NAND2xp33_ASAP7_75t_L g1096 ( 
.A(n_903),
.B(n_663),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_943),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_947),
.B(n_526),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_918),
.B(n_893),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_897),
.A2(n_788),
.B(n_748),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_892),
.A2(n_357),
.B1(n_358),
.B2(n_362),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_893),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_945),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_933),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_913),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_894),
.B(n_526),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_884),
.B(n_527),
.Y(n_1107)
);

NAND2x1p5_ASAP7_75t_L g1108 ( 
.A(n_836),
.B(n_654),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_SL g1109 ( 
.A1(n_906),
.A2(n_331),
.B1(n_428),
.B2(n_256),
.Y(n_1109)
);

OAI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_857),
.A2(n_877),
.B1(n_894),
.B2(n_898),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_904),
.A2(n_797),
.B(n_708),
.C(n_692),
.Y(n_1111)
);

OR2x2_ASAP7_75t_SL g1112 ( 
.A(n_924),
.B(n_527),
.Y(n_1112)
);

BUFx3_ASAP7_75t_L g1113 ( 
.A(n_919),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_916),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_917),
.B(n_701),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_921),
.B(n_701),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_887),
.B(n_934),
.Y(n_1117)
);

CKINVDCx16_ASAP7_75t_R g1118 ( 
.A(n_930),
.Y(n_1118)
);

INVx2_ASAP7_75t_SL g1119 ( 
.A(n_958),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_996),
.B(n_948),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_970),
.B(n_931),
.Y(n_1121)
);

NAND3xp33_ASAP7_75t_L g1122 ( 
.A(n_993),
.B(n_909),
.C(n_880),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_962),
.Y(n_1123)
);

INVx3_ASAP7_75t_SL g1124 ( 
.A(n_1021),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_962),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_965),
.Y(n_1126)
);

INVx4_ASAP7_75t_L g1127 ( 
.A(n_991),
.Y(n_1127)
);

INVx2_ASAP7_75t_SL g1128 ( 
.A(n_1002),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_1118),
.B(n_907),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1035),
.A2(n_869),
.B(n_950),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_959),
.B(n_912),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1052),
.A2(n_915),
.B(n_932),
.C(n_876),
.Y(n_1132)
);

OAI22x1_ASAP7_75t_L g1133 ( 
.A1(n_1039),
.A2(n_377),
.B1(n_383),
.B2(n_389),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_959),
.A2(n_748),
.B(n_835),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_R g1135 ( 
.A(n_1006),
.B(n_841),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1099),
.A2(n_880),
.B1(n_876),
.B2(n_394),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1009),
.B(n_665),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1043),
.A2(n_1045),
.B(n_1031),
.Y(n_1138)
);

BUFx8_ASAP7_75t_L g1139 ( 
.A(n_978),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_SL g1140 ( 
.A1(n_981),
.A2(n_332),
.B1(n_256),
.B2(n_335),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_986),
.B(n_665),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1109),
.A2(n_396),
.B1(n_390),
.B2(n_395),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1003),
.B(n_665),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1043),
.A2(n_852),
.B(n_745),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_962),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_1070),
.B(n_590),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1007),
.B(n_1104),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1102),
.B(n_686),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_952),
.A2(n_938),
.B1(n_528),
.B2(n_529),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_963),
.B(n_528),
.Y(n_1150)
);

O2A1O1Ixp5_ASAP7_75t_L g1151 ( 
.A1(n_994),
.A2(n_938),
.B(n_683),
.C(n_736),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_964),
.A2(n_529),
.B1(n_332),
.B2(n_335),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1012),
.A2(n_1040),
.B1(n_1094),
.B2(n_1082),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_1080),
.B(n_797),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_971),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_971),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_1036),
.Y(n_1157)
);

AOI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1025),
.A2(n_683),
.B(n_647),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_964),
.A2(n_969),
.B1(n_979),
.B2(n_973),
.Y(n_1159)
);

O2A1O1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_1069),
.A2(n_787),
.B(n_643),
.C(n_650),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_1047),
.B(n_399),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1106),
.B(n_686),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_953),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1107),
.B(n_692),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1043),
.A2(n_745),
.B(n_785),
.Y(n_1165)
);

NOR2xp67_ASAP7_75t_L g1166 ( 
.A(n_1093),
.B(n_399),
.Y(n_1166)
);

AND2x6_ASAP7_75t_L g1167 ( 
.A(n_971),
.B(n_331),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1028),
.A2(n_1058),
.B1(n_1076),
.B2(n_951),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1078),
.A2(n_797),
.B(n_692),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_1070),
.B(n_590),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1031),
.A2(n_785),
.B(n_777),
.Y(n_1171)
);

NOR3xp33_ASAP7_75t_SL g1172 ( 
.A(n_954),
.B(n_400),
.C(n_409),
.Y(n_1172)
);

NOR2xp67_ASAP7_75t_SL g1173 ( 
.A(n_992),
.B(n_400),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_972),
.B(n_736),
.Y(n_1174)
);

INVxp67_ASAP7_75t_L g1175 ( 
.A(n_967),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1046),
.A2(n_785),
.B(n_777),
.Y(n_1176)
);

NOR3xp33_ASAP7_75t_SL g1177 ( 
.A(n_1059),
.B(n_409),
.C(n_413),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_988),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_982),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_988),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1019),
.B(n_743),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1079),
.A2(n_743),
.B1(n_704),
.B2(n_663),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1046),
.A2(n_785),
.B(n_777),
.Y(n_1183)
);

NOR2xp67_ASAP7_75t_L g1184 ( 
.A(n_1027),
.B(n_413),
.Y(n_1184)
);

AOI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1072),
.A2(n_419),
.B1(n_421),
.B2(n_428),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1051),
.A2(n_777),
.B(n_745),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1055),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1086),
.B(n_422),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_989),
.B(n_629),
.Y(n_1189)
);

CKINVDCx14_ASAP7_75t_R g1190 ( 
.A(n_1014),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_990),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1051),
.A2(n_745),
.B(n_726),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1033),
.B(n_591),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_969),
.A2(n_423),
.B1(n_427),
.B2(n_424),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1057),
.A2(n_423),
.B1(n_427),
.B2(n_424),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_984),
.A2(n_599),
.B(n_593),
.C(n_591),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1090),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_990),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1078),
.A2(n_637),
.B(n_629),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1065),
.A2(n_1061),
.B(n_1096),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1090),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_992),
.B(n_663),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_R g1203 ( 
.A(n_983),
.B(n_82),
.Y(n_1203)
);

A2O1A1Ixp33_ASAP7_75t_SL g1204 ( 
.A1(n_1010),
.A2(n_593),
.B(n_599),
.C(n_633),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_956),
.B(n_663),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_982),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_992),
.B(n_726),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_995),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1032),
.B(n_633),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1065),
.A2(n_745),
.B(n_726),
.Y(n_1210)
);

BUFx2_ASAP7_75t_L g1211 ( 
.A(n_1008),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1037),
.B(n_726),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_977),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_957),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_1013),
.B(n_684),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_977),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_995),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1066),
.B(n_984),
.Y(n_1218)
);

INVxp67_ASAP7_75t_L g1219 ( 
.A(n_1008),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1033),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1089),
.B(n_0),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_974),
.A2(n_752),
.B(n_717),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1001),
.Y(n_1223)
);

INVx4_ASAP7_75t_L g1224 ( 
.A(n_1013),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1084),
.B(n_1),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_974),
.A2(n_483),
.B1(n_476),
.B2(n_477),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_977),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1038),
.B(n_637),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1087),
.A2(n_479),
.B1(n_476),
.B2(n_477),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1004),
.A2(n_474),
.B1(n_478),
.B2(n_479),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1041),
.B(n_637),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_968),
.Y(n_1232)
);

AOI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1030),
.A2(n_478),
.B1(n_474),
.B2(n_549),
.Y(n_1233)
);

OAI22x1_ASAP7_75t_L g1234 ( 
.A1(n_1056),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_1234)
);

OR2x2_ASAP7_75t_L g1235 ( 
.A(n_1112),
.B(n_1098),
.Y(n_1235)
);

INVx4_ASAP7_75t_L g1236 ( 
.A(n_980),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1083),
.A2(n_752),
.B(n_717),
.Y(n_1237)
);

AOI222xp33_ASAP7_75t_L g1238 ( 
.A1(n_1016),
.A2(n_9),
.B1(n_10),
.B2(n_14),
.C1(n_18),
.C2(n_19),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1001),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1070),
.B(n_83),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1049),
.B(n_549),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_SL g1242 ( 
.A1(n_1018),
.A2(n_9),
.B1(n_20),
.B2(n_22),
.Y(n_1242)
);

OA21x2_ASAP7_75t_L g1243 ( 
.A1(n_1111),
.A2(n_1083),
.B(n_955),
.Y(n_1243)
);

O2A1O1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1018),
.A2(n_22),
.B(n_23),
.C(n_25),
.Y(n_1244)
);

O2A1O1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1101),
.A2(n_23),
.B(n_26),
.C(n_27),
.Y(n_1245)
);

NOR3xp33_ASAP7_75t_SL g1246 ( 
.A(n_1101),
.B(n_33),
.C(n_34),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_1114),
.A2(n_549),
.B(n_717),
.C(n_684),
.Y(n_1247)
);

OAI21xp33_ASAP7_75t_L g1248 ( 
.A1(n_1092),
.A2(n_549),
.B(n_35),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_966),
.B(n_33),
.Y(n_1249)
);

O2A1O1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1017),
.A2(n_38),
.B(n_39),
.C(n_41),
.Y(n_1250)
);

CKINVDCx16_ASAP7_75t_R g1251 ( 
.A(n_1088),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1054),
.B(n_1060),
.Y(n_1252)
);

CKINVDCx16_ASAP7_75t_R g1253 ( 
.A(n_1068),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_998),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1067),
.B(n_752),
.Y(n_1255)
);

INVx4_ASAP7_75t_L g1256 ( 
.A(n_980),
.Y(n_1256)
);

A2O1A1Ixp33_ASAP7_75t_L g1257 ( 
.A1(n_955),
.A2(n_752),
.B(n_717),
.C(n_684),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_983),
.B(n_1011),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1034),
.B(n_123),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1074),
.B(n_684),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1063),
.A2(n_115),
.B(n_211),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1029),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1134),
.A2(n_1110),
.B(n_1100),
.Y(n_1263)
);

AOI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1218),
.A2(n_1073),
.B1(n_961),
.B2(n_960),
.Y(n_1264)
);

AO32x2_ASAP7_75t_L g1265 ( 
.A1(n_1159),
.A2(n_1149),
.A3(n_1152),
.B1(n_1136),
.B2(n_1229),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_1128),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1147),
.A2(n_1011),
.B1(n_1081),
.B2(n_980),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1131),
.A2(n_1015),
.B(n_976),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1126),
.Y(n_1269)
);

A2O1A1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1121),
.A2(n_1077),
.B(n_1085),
.C(n_997),
.Y(n_1270)
);

BUFx12f_ASAP7_75t_L g1271 ( 
.A(n_1139),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1237),
.A2(n_985),
.B(n_1023),
.Y(n_1272)
);

AO31x2_ASAP7_75t_L g1273 ( 
.A1(n_1247),
.A2(n_1105),
.A3(n_1023),
.B(n_1116),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1188),
.A2(n_1024),
.B1(n_1026),
.B2(n_1095),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1122),
.A2(n_997),
.B(n_1116),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1122),
.A2(n_1115),
.B(n_1117),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1178),
.B(n_1180),
.Y(n_1277)
);

NAND3xp33_ASAP7_75t_SL g1278 ( 
.A(n_1238),
.B(n_1153),
.C(n_1140),
.Y(n_1278)
);

NAND3xp33_ASAP7_75t_L g1279 ( 
.A(n_1225),
.B(n_1073),
.C(n_975),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1119),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1139),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1191),
.B(n_1198),
.Y(n_1282)
);

INVxp67_ASAP7_75t_L g1283 ( 
.A(n_1157),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1200),
.A2(n_1138),
.B(n_1144),
.Y(n_1284)
);

OAI22x1_ASAP7_75t_L g1285 ( 
.A1(n_1168),
.A2(n_1081),
.B1(n_987),
.B2(n_1062),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1123),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1252),
.B(n_1000),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1259),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1130),
.A2(n_1108),
.B(n_1071),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1181),
.A2(n_976),
.B(n_1005),
.Y(n_1290)
);

AOI221x1_ASAP7_75t_L g1291 ( 
.A1(n_1248),
.A2(n_1117),
.B1(n_1095),
.B2(n_1103),
.C(n_1097),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1259),
.Y(n_1292)
);

A2O1A1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1184),
.A2(n_1053),
.B(n_1042),
.C(n_1050),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1211),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1208),
.A2(n_1073),
.B1(n_1042),
.B2(n_1091),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1217),
.B(n_1095),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1223),
.B(n_1026),
.Y(n_1297)
);

AO31x2_ASAP7_75t_L g1298 ( 
.A1(n_1132),
.A2(n_1044),
.A3(n_1064),
.B(n_1048),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1239),
.B(n_1026),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1171),
.A2(n_1071),
.B(n_1022),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1189),
.A2(n_1005),
.B(n_1015),
.Y(n_1301)
);

OA22x2_ASAP7_75t_L g1302 ( 
.A1(n_1234),
.A2(n_1034),
.B1(n_1020),
.B2(n_999),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1120),
.B(n_1193),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1150),
.B(n_1020),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1258),
.B(n_1113),
.Y(n_1305)
);

AO31x2_ASAP7_75t_L g1306 ( 
.A1(n_1257),
.A2(n_1091),
.A3(n_1075),
.B(n_48),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1124),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1176),
.A2(n_1091),
.B(n_132),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_1219),
.B(n_1091),
.Y(n_1309)
);

OA21x2_ASAP7_75t_L g1310 ( 
.A1(n_1169),
.A2(n_108),
.B(n_207),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1175),
.B(n_41),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1183),
.A2(n_107),
.B(n_202),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1137),
.A2(n_1141),
.B(n_1210),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1146),
.B(n_214),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1235),
.B(n_47),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1186),
.A2(n_104),
.B(n_193),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1151),
.A2(n_200),
.B(n_102),
.Y(n_1317)
);

A2O1A1Ixp33_ASAP7_75t_L g1318 ( 
.A1(n_1249),
.A2(n_50),
.B(n_52),
.C(n_54),
.Y(n_1318)
);

OA21x2_ASAP7_75t_L g1319 ( 
.A1(n_1192),
.A2(n_133),
.B(n_185),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1214),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1243),
.A2(n_92),
.B(n_183),
.Y(n_1321)
);

AO31x2_ASAP7_75t_L g1322 ( 
.A1(n_1136),
.A2(n_52),
.A3(n_54),
.B(n_55),
.Y(n_1322)
);

AO31x2_ASAP7_75t_L g1323 ( 
.A1(n_1149),
.A2(n_55),
.A3(n_57),
.B(n_61),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1232),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1174),
.B(n_63),
.Y(n_1325)
);

BUFx10_ASAP7_75t_L g1326 ( 
.A(n_1221),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1254),
.Y(n_1327)
);

A2O1A1Ixp33_ASAP7_75t_L g1328 ( 
.A1(n_1244),
.A2(n_63),
.B(n_66),
.C(n_68),
.Y(n_1328)
);

OAI22x1_ASAP7_75t_L g1329 ( 
.A1(n_1233),
.A2(n_1129),
.B1(n_1161),
.B2(n_1163),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1152),
.B(n_68),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1262),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1162),
.A2(n_145),
.B(n_160),
.Y(n_1332)
);

INVxp67_ASAP7_75t_L g1333 ( 
.A(n_1179),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1209),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1165),
.A2(n_162),
.B(n_158),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1222),
.A2(n_152),
.B(n_70),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1220),
.B(n_73),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_SL g1338 ( 
.A1(n_1240),
.A2(n_69),
.B(n_70),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1241),
.A2(n_1228),
.B(n_1231),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1206),
.B(n_69),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_SL g1341 ( 
.A(n_1245),
.B(n_71),
.Y(n_1341)
);

OA21x2_ASAP7_75t_L g1342 ( 
.A1(n_1212),
.A2(n_72),
.B(n_1261),
.Y(n_1342)
);

AO31x2_ASAP7_75t_L g1343 ( 
.A1(n_1229),
.A2(n_1182),
.A3(n_1230),
.B(n_1255),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1187),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1253),
.B(n_1133),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1146),
.B(n_1170),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1194),
.B(n_1154),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_1194),
.B(n_1201),
.Y(n_1348)
);

OAI22x1_ASAP7_75t_L g1349 ( 
.A1(n_1238),
.A2(n_1205),
.B1(n_1240),
.B2(n_1170),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1143),
.A2(n_1160),
.B(n_1243),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1197),
.B(n_1172),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1166),
.B(n_1148),
.Y(n_1352)
);

AOI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1202),
.A2(n_1207),
.B(n_1260),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1164),
.A2(n_1204),
.B(n_1215),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1135),
.B(n_1177),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1230),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1190),
.B(n_1142),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1185),
.B(n_1203),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_SL g1359 ( 
.A(n_1123),
.B(n_1213),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1142),
.B(n_1242),
.Y(n_1360)
);

AOI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1173),
.A2(n_1226),
.B(n_1195),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1127),
.A2(n_1224),
.B(n_1196),
.Y(n_1362)
);

OAI21xp33_ASAP7_75t_SL g1363 ( 
.A1(n_1127),
.A2(n_1224),
.B(n_1256),
.Y(n_1363)
);

AOI221xp5_ASAP7_75t_SL g1364 ( 
.A1(n_1250),
.A2(n_1195),
.B1(n_1246),
.B2(n_1125),
.C(n_1145),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1167),
.A2(n_1236),
.B(n_1123),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1125),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1145),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1155),
.B(n_1156),
.Y(n_1368)
);

INVx4_ASAP7_75t_L g1369 ( 
.A(n_1155),
.Y(n_1369)
);

NOR4xp25_ASAP7_75t_L g1370 ( 
.A(n_1167),
.B(n_1251),
.C(n_1156),
.D(n_1213),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1213),
.A2(n_1216),
.B(n_1227),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1216),
.B(n_1227),
.Y(n_1372)
);

AOI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1158),
.A2(n_1134),
.B(n_1200),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1119),
.Y(n_1374)
);

OA21x2_ASAP7_75t_L g1375 ( 
.A1(n_1199),
.A2(n_1169),
.B(n_1151),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1237),
.A2(n_1199),
.B(n_1130),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1235),
.B(n_693),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_SL g1378 ( 
.A(n_1175),
.B(n_1118),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1175),
.B(n_970),
.Y(n_1379)
);

AO32x2_ASAP7_75t_L g1380 ( 
.A1(n_1159),
.A2(n_981),
.A3(n_1149),
.B1(n_1152),
.B2(n_1136),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1134),
.A2(n_1131),
.B(n_959),
.Y(n_1381)
);

AOI21xp33_ASAP7_75t_L g1382 ( 
.A1(n_1121),
.A2(n_993),
.B(n_1052),
.Y(n_1382)
);

AOI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1218),
.A2(n_993),
.B1(n_981),
.B2(n_1012),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1121),
.B(n_996),
.Y(n_1384)
);

NAND2xp33_ASAP7_75t_R g1385 ( 
.A(n_1135),
.B(n_666),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1126),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_SL g1387 ( 
.A(n_1218),
.B(n_981),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1121),
.B(n_996),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1126),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1122),
.A2(n_993),
.B(n_1052),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_1175),
.B(n_970),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1150),
.B(n_693),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1124),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1124),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1237),
.A2(n_1199),
.B(n_1130),
.Y(n_1395)
);

BUFx6f_ASAP7_75t_L g1396 ( 
.A(n_1123),
.Y(n_1396)
);

OR2x6_ASAP7_75t_L g1397 ( 
.A(n_1258),
.B(n_1128),
.Y(n_1397)
);

AO31x2_ASAP7_75t_L g1398 ( 
.A1(n_1247),
.A2(n_994),
.A3(n_1159),
.B(n_1132),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1258),
.B(n_1070),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1235),
.B(n_693),
.Y(n_1400)
);

OAI21xp33_ASAP7_75t_L g1401 ( 
.A1(n_1188),
.A2(n_993),
.B(n_1218),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_1124),
.Y(n_1402)
);

INVx2_ASAP7_75t_SL g1403 ( 
.A(n_1128),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1258),
.B(n_1070),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1237),
.A2(n_1199),
.B(n_1130),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1237),
.A2(n_1199),
.B(n_1130),
.Y(n_1406)
);

AOI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1218),
.A2(n_993),
.B1(n_981),
.B2(n_1012),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1259),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1147),
.A2(n_993),
.B1(n_804),
.B2(n_1191),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1237),
.A2(n_1199),
.B(n_1130),
.Y(n_1410)
);

CKINVDCx11_ASAP7_75t_R g1411 ( 
.A(n_1124),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1134),
.A2(n_1131),
.B(n_959),
.Y(n_1412)
);

OAI22x1_ASAP7_75t_L g1413 ( 
.A1(n_1218),
.A2(n_993),
.B1(n_1188),
.B2(n_1039),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1147),
.A2(n_993),
.B1(n_804),
.B2(n_1191),
.Y(n_1414)
);

CKINVDCx16_ASAP7_75t_R g1415 ( 
.A(n_1385),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1269),
.Y(n_1416)
);

NOR2xp67_ASAP7_75t_L g1417 ( 
.A(n_1283),
.B(n_1403),
.Y(n_1417)
);

INVx5_ASAP7_75t_L g1418 ( 
.A(n_1286),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1278),
.A2(n_1401),
.B1(n_1387),
.B2(n_1360),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1401),
.B(n_1387),
.Y(n_1420)
);

INVxp67_ASAP7_75t_SL g1421 ( 
.A(n_1282),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1289),
.A2(n_1395),
.B(n_1376),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1405),
.A2(n_1410),
.B(n_1406),
.Y(n_1423)
);

INVx1_ASAP7_75t_SL g1424 ( 
.A(n_1374),
.Y(n_1424)
);

AOI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1373),
.A2(n_1354),
.B(n_1263),
.Y(n_1425)
);

AOI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1361),
.A2(n_1412),
.B(n_1381),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1384),
.A2(n_1388),
.B1(n_1407),
.B2(n_1383),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1306),
.Y(n_1428)
);

AO31x2_ASAP7_75t_L g1429 ( 
.A1(n_1284),
.A2(n_1291),
.A3(n_1313),
.B(n_1295),
.Y(n_1429)
);

AO21x2_ASAP7_75t_L g1430 ( 
.A1(n_1317),
.A2(n_1390),
.B(n_1275),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1280),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1272),
.A2(n_1308),
.B(n_1350),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1288),
.B(n_1292),
.Y(n_1433)
);

OR2x6_ASAP7_75t_L g1434 ( 
.A(n_1349),
.B(n_1397),
.Y(n_1434)
);

INVx1_ASAP7_75t_SL g1435 ( 
.A(n_1294),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_1303),
.B(n_1378),
.Y(n_1436)
);

AOI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1301),
.A2(n_1295),
.B(n_1290),
.Y(n_1437)
);

OR2x6_ASAP7_75t_L g1438 ( 
.A(n_1397),
.B(n_1338),
.Y(n_1438)
);

AOI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1339),
.A2(n_1353),
.B(n_1268),
.Y(n_1439)
);

AOI21xp33_ASAP7_75t_L g1440 ( 
.A1(n_1413),
.A2(n_1279),
.B(n_1409),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_SL g1441 ( 
.A1(n_1264),
.A2(n_1321),
.B(n_1362),
.Y(n_1441)
);

AO21x2_ASAP7_75t_L g1442 ( 
.A1(n_1390),
.A2(n_1275),
.B(n_1321),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1266),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1379),
.B(n_1391),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1392),
.B(n_1334),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1300),
.A2(n_1312),
.B(n_1336),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1377),
.B(n_1400),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1282),
.B(n_1277),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1382),
.A2(n_1330),
.B1(n_1341),
.B2(n_1279),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1304),
.B(n_1347),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1264),
.A2(n_1274),
.B1(n_1288),
.B2(n_1292),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1414),
.B(n_1341),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1287),
.B(n_1346),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1276),
.A2(n_1316),
.B(n_1375),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1358),
.A2(n_1311),
.B1(n_1325),
.B2(n_1357),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1270),
.A2(n_1352),
.B(n_1276),
.Y(n_1456)
);

INVx4_ASAP7_75t_SL g1457 ( 
.A(n_1323),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1375),
.A2(n_1335),
.B(n_1319),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1397),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1306),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1319),
.A2(n_1332),
.B(n_1267),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1315),
.A2(n_1285),
.B1(n_1326),
.B2(n_1302),
.Y(n_1462)
);

INVx1_ASAP7_75t_SL g1463 ( 
.A(n_1372),
.Y(n_1463)
);

OA21x2_ASAP7_75t_L g1464 ( 
.A1(n_1364),
.A2(n_1356),
.B(n_1293),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1310),
.A2(n_1342),
.B(n_1267),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1346),
.B(n_1305),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1310),
.A2(n_1342),
.B(n_1365),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1326),
.A2(n_1329),
.B1(n_1345),
.B2(n_1348),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1306),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1367),
.Y(n_1470)
);

OA21x2_ASAP7_75t_L g1471 ( 
.A1(n_1364),
.A2(n_1328),
.B(n_1296),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1305),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_SL g1473 ( 
.A(n_1408),
.B(n_1370),
.Y(n_1473)
);

INVx1_ASAP7_75t_SL g1474 ( 
.A(n_1307),
.Y(n_1474)
);

NAND3xp33_ASAP7_75t_L g1475 ( 
.A(n_1318),
.B(n_1355),
.C(n_1351),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1314),
.A2(n_1320),
.B1(n_1408),
.B2(n_1340),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1297),
.B(n_1299),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1333),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1399),
.B(n_1404),
.Y(n_1479)
);

OA21x2_ASAP7_75t_L g1480 ( 
.A1(n_1386),
.A2(n_1389),
.B(n_1398),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1324),
.B(n_1331),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1368),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1399),
.B(n_1404),
.Y(n_1483)
);

AO21x2_ASAP7_75t_L g1484 ( 
.A1(n_1370),
.A2(n_1359),
.B(n_1371),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1298),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1327),
.B(n_1344),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1337),
.B(n_1309),
.Y(n_1487)
);

OA21x2_ASAP7_75t_L g1488 ( 
.A1(n_1273),
.A2(n_1265),
.B(n_1298),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_1393),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1363),
.A2(n_1265),
.B(n_1309),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1366),
.B(n_1286),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1286),
.Y(n_1492)
);

INVx2_ASAP7_75t_SL g1493 ( 
.A(n_1281),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1343),
.A2(n_1265),
.B(n_1363),
.Y(n_1494)
);

CKINVDCx11_ASAP7_75t_R g1495 ( 
.A(n_1411),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1380),
.B(n_1396),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1396),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1394),
.Y(n_1498)
);

NAND2x1p5_ASAP7_75t_L g1499 ( 
.A(n_1369),
.B(n_1396),
.Y(n_1499)
);

A2O1A1Ixp33_ASAP7_75t_L g1500 ( 
.A1(n_1322),
.A2(n_1402),
.B(n_1369),
.C(n_1271),
.Y(n_1500)
);

AOI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1381),
.A2(n_1412),
.B(n_1284),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1278),
.A2(n_1401),
.B1(n_981),
.B2(n_1040),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1306),
.Y(n_1503)
);

AO32x2_ASAP7_75t_L g1504 ( 
.A1(n_1409),
.A2(n_1414),
.A3(n_981),
.B1(n_1295),
.B2(n_1159),
.Y(n_1504)
);

NAND2x1p5_ASAP7_75t_L g1505 ( 
.A(n_1288),
.B(n_1292),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1278),
.A2(n_1401),
.B1(n_981),
.B2(n_1040),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1384),
.B(n_1388),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1278),
.A2(n_1401),
.B1(n_981),
.B2(n_1040),
.Y(n_1508)
);

BUFx2_ASAP7_75t_L g1509 ( 
.A(n_1280),
.Y(n_1509)
);

OAI211xp5_ASAP7_75t_L g1510 ( 
.A1(n_1401),
.A2(n_1238),
.B(n_873),
.C(n_1383),
.Y(n_1510)
);

OAI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1387),
.A2(n_1278),
.B1(n_1341),
.B2(n_1360),
.Y(n_1511)
);

A2O1A1Ixp33_ASAP7_75t_L g1512 ( 
.A1(n_1401),
.A2(n_993),
.B(n_1317),
.C(n_1278),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1288),
.B(n_1292),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1376),
.A2(n_1405),
.B(n_1395),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1411),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1266),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1298),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1384),
.B(n_1388),
.Y(n_1518)
);

OAI22x1_ASAP7_75t_L g1519 ( 
.A1(n_1383),
.A2(n_1407),
.B1(n_1218),
.B2(n_1264),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1376),
.A2(n_1405),
.B(n_1395),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1298),
.Y(n_1521)
);

INVx8_ASAP7_75t_L g1522 ( 
.A(n_1286),
.Y(n_1522)
);

AOI22x1_ASAP7_75t_L g1523 ( 
.A1(n_1413),
.A2(n_1285),
.B1(n_1349),
.B2(n_1329),
.Y(n_1523)
);

CKINVDCx12_ASAP7_75t_R g1524 ( 
.A(n_1397),
.Y(n_1524)
);

AOI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1381),
.A2(n_1412),
.B(n_1284),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1269),
.Y(n_1526)
);

OAI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1401),
.A2(n_993),
.B(n_996),
.Y(n_1527)
);

O2A1O1Ixp33_ASAP7_75t_SL g1528 ( 
.A1(n_1278),
.A2(n_1328),
.B(n_1317),
.C(n_1318),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1384),
.B(n_1388),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_SL g1530 ( 
.A(n_1307),
.B(n_666),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1269),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1392),
.B(n_1303),
.Y(n_1532)
);

INVx1_ASAP7_75t_SL g1533 ( 
.A(n_1374),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1298),
.Y(n_1534)
);

INVx2_ASAP7_75t_SL g1535 ( 
.A(n_1266),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1269),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1384),
.B(n_1388),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1298),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1384),
.B(n_1388),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1392),
.B(n_1303),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1288),
.B(n_1292),
.Y(n_1541)
);

A2O1A1Ixp33_ASAP7_75t_L g1542 ( 
.A1(n_1401),
.A2(n_993),
.B(n_1317),
.C(n_1278),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1384),
.B(n_1388),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1266),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_SL g1545 ( 
.A1(n_1264),
.A2(n_1317),
.B(n_1321),
.Y(n_1545)
);

NOR2xp67_ASAP7_75t_L g1546 ( 
.A(n_1283),
.B(n_963),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1269),
.Y(n_1547)
);

OAI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1376),
.A2(n_1405),
.B(n_1395),
.Y(n_1548)
);

OAI22xp33_ASAP7_75t_SL g1549 ( 
.A1(n_1387),
.A2(n_1341),
.B1(n_1360),
.B2(n_1330),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1376),
.A2(n_1405),
.B(n_1395),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1288),
.B(n_1292),
.Y(n_1551)
);

AOI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1401),
.A2(n_1387),
.B1(n_1188),
.B2(n_970),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1298),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1411),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1298),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1306),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1288),
.B(n_1292),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1384),
.B(n_1388),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1269),
.Y(n_1559)
);

AO31x2_ASAP7_75t_L g1560 ( 
.A1(n_1263),
.A2(n_1284),
.A3(n_1412),
.B(n_1381),
.Y(n_1560)
);

OAI21x1_ASAP7_75t_L g1561 ( 
.A1(n_1376),
.A2(n_1405),
.B(n_1395),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1269),
.Y(n_1562)
);

A2O1A1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1401),
.A2(n_993),
.B(n_1317),
.C(n_1278),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1298),
.Y(n_1564)
);

AOI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1381),
.A2(n_1412),
.B(n_1284),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1384),
.B(n_1388),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1288),
.B(n_1292),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1436),
.B(n_1453),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1512),
.A2(n_1563),
.B(n_1542),
.Y(n_1569)
);

NOR2xp67_ASAP7_75t_L g1570 ( 
.A(n_1498),
.B(n_1475),
.Y(n_1570)
);

HB1xp67_ASAP7_75t_L g1571 ( 
.A(n_1482),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1419),
.A2(n_1510),
.B1(n_1552),
.B2(n_1542),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1532),
.B(n_1540),
.Y(n_1573)
);

NOR2xp67_ASAP7_75t_L g1574 ( 
.A(n_1443),
.B(n_1535),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1528),
.A2(n_1430),
.B(n_1545),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1419),
.A2(n_1502),
.B1(n_1508),
.B2(n_1506),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1450),
.B(n_1427),
.Y(n_1577)
);

OAI31xp33_ASAP7_75t_L g1578 ( 
.A1(n_1511),
.A2(n_1549),
.A3(n_1508),
.B(n_1502),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1463),
.B(n_1487),
.Y(n_1579)
);

OA22x2_ASAP7_75t_L g1580 ( 
.A1(n_1519),
.A2(n_1434),
.B1(n_1438),
.B2(n_1473),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1516),
.Y(n_1581)
);

AOI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1528),
.A2(n_1430),
.B(n_1452),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1447),
.B(n_1466),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1420),
.B(n_1449),
.Y(n_1584)
);

OA21x2_ASAP7_75t_L g1585 ( 
.A1(n_1465),
.A2(n_1467),
.B(n_1458),
.Y(n_1585)
);

O2A1O1Ixp33_ASAP7_75t_L g1586 ( 
.A1(n_1511),
.A2(n_1440),
.B(n_1420),
.C(n_1527),
.Y(n_1586)
);

A2O1A1Ixp33_ASAP7_75t_L g1587 ( 
.A1(n_1506),
.A2(n_1449),
.B(n_1455),
.C(n_1456),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1483),
.B(n_1479),
.Y(n_1588)
);

AOI221x1_ASAP7_75t_SL g1589 ( 
.A1(n_1507),
.A2(n_1537),
.B1(n_1558),
.B2(n_1539),
.C(n_1566),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1455),
.A2(n_1518),
.B1(n_1529),
.B2(n_1543),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1496),
.B(n_1477),
.Y(n_1591)
);

OA21x2_ASAP7_75t_L g1592 ( 
.A1(n_1461),
.A2(n_1432),
.B(n_1446),
.Y(n_1592)
);

BUFx12f_ASAP7_75t_L g1593 ( 
.A(n_1495),
.Y(n_1593)
);

AOI21x1_ASAP7_75t_SL g1594 ( 
.A1(n_1428),
.A2(n_1469),
.B(n_1460),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1464),
.B(n_1490),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1495),
.Y(n_1596)
);

XOR2xp5_ASAP7_75t_L g1597 ( 
.A(n_1515),
.B(n_1554),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1462),
.B(n_1468),
.Y(n_1598)
);

O2A1O1Ixp33_ASAP7_75t_L g1599 ( 
.A1(n_1500),
.A2(n_1441),
.B(n_1444),
.C(n_1451),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1445),
.B(n_1435),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1462),
.B(n_1468),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1434),
.B(n_1478),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1464),
.B(n_1442),
.Y(n_1603)
);

O2A1O1Ixp33_ASAP7_75t_L g1604 ( 
.A1(n_1438),
.A2(n_1533),
.B(n_1424),
.C(n_1476),
.Y(n_1604)
);

O2A1O1Ixp33_ASAP7_75t_L g1605 ( 
.A1(n_1438),
.A2(n_1476),
.B(n_1493),
.C(n_1536),
.Y(n_1605)
);

INVx6_ASAP7_75t_L g1606 ( 
.A(n_1418),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_SL g1607 ( 
.A1(n_1433),
.A2(n_1513),
.B(n_1541),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1524),
.Y(n_1608)
);

AOI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1415),
.A2(n_1530),
.B1(n_1474),
.B2(n_1489),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1464),
.B(n_1471),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_SL g1611 ( 
.A1(n_1513),
.A2(n_1551),
.B(n_1567),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1471),
.B(n_1480),
.Y(n_1612)
);

O2A1O1Ixp33_ASAP7_75t_L g1613 ( 
.A1(n_1526),
.A2(n_1531),
.B(n_1562),
.C(n_1559),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1547),
.B(n_1480),
.Y(n_1614)
);

NOR2xp67_ASAP7_75t_L g1615 ( 
.A(n_1546),
.B(n_1417),
.Y(n_1615)
);

O2A1O1Ixp33_ASAP7_75t_L g1616 ( 
.A1(n_1503),
.A2(n_1556),
.B(n_1509),
.C(n_1431),
.Y(n_1616)
);

BUFx2_ASAP7_75t_L g1617 ( 
.A(n_1516),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1523),
.A2(n_1481),
.B1(n_1486),
.B2(n_1544),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1541),
.B(n_1567),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1418),
.A2(n_1505),
.B1(n_1491),
.B2(n_1470),
.Y(n_1620)
);

AOI21xp5_ASAP7_75t_SL g1621 ( 
.A1(n_1557),
.A2(n_1499),
.B(n_1484),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_1515),
.Y(n_1622)
);

OA21x2_ASAP7_75t_L g1623 ( 
.A1(n_1494),
.A2(n_1561),
.B(n_1514),
.Y(n_1623)
);

AOI21xp5_ASAP7_75t_SL g1624 ( 
.A1(n_1499),
.A2(n_1484),
.B(n_1492),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1522),
.Y(n_1625)
);

A2O1A1Ixp33_ASAP7_75t_L g1626 ( 
.A1(n_1504),
.A2(n_1521),
.B(n_1555),
.C(n_1553),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_1522),
.Y(n_1627)
);

CKINVDCx20_ASAP7_75t_R g1628 ( 
.A(n_1522),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1457),
.B(n_1488),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1497),
.B(n_1504),
.Y(n_1630)
);

OA21x2_ASAP7_75t_L g1631 ( 
.A1(n_1423),
.A2(n_1561),
.B(n_1520),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1457),
.B(n_1488),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1418),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1485),
.A2(n_1564),
.B1(n_1521),
.B2(n_1534),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1457),
.B(n_1517),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1504),
.B(n_1429),
.Y(n_1636)
);

O2A1O1Ixp33_ASAP7_75t_L g1637 ( 
.A1(n_1485),
.A2(n_1534),
.B(n_1553),
.C(n_1538),
.Y(n_1637)
);

AOI221x1_ASAP7_75t_SL g1638 ( 
.A1(n_1504),
.A2(n_1429),
.B1(n_1437),
.B2(n_1426),
.C(n_1560),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1429),
.B(n_1560),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1429),
.B(n_1425),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1439),
.B(n_1422),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1548),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1550),
.Y(n_1643)
);

A2O1A1Ixp33_ASAP7_75t_L g1644 ( 
.A1(n_1552),
.A2(n_1401),
.B(n_1420),
.C(n_1452),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1532),
.B(n_1540),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1459),
.B(n_1482),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_1495),
.Y(n_1647)
);

OA22x2_ASAP7_75t_L g1648 ( 
.A1(n_1552),
.A2(n_1510),
.B1(n_981),
.B2(n_1407),
.Y(n_1648)
);

CKINVDCx6p67_ASAP7_75t_R g1649 ( 
.A(n_1495),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1472),
.Y(n_1650)
);

OA21x2_ASAP7_75t_L g1651 ( 
.A1(n_1465),
.A2(n_1467),
.B(n_1454),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1419),
.A2(n_1510),
.B1(n_1552),
.B2(n_1542),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1532),
.B(n_1540),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1532),
.B(n_1540),
.Y(n_1654)
);

O2A1O1Ixp33_ASAP7_75t_L g1655 ( 
.A1(n_1512),
.A2(n_1278),
.B(n_1563),
.C(n_1542),
.Y(n_1655)
);

A2O1A1Ixp33_ASAP7_75t_L g1656 ( 
.A1(n_1552),
.A2(n_1401),
.B(n_1420),
.C(n_1452),
.Y(n_1656)
);

AND2x4_ASAP7_75t_SL g1657 ( 
.A(n_1466),
.B(n_1305),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1421),
.B(n_1448),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1501),
.A2(n_1565),
.B(n_1525),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1419),
.A2(n_1510),
.B1(n_1552),
.B2(n_1542),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_1495),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1532),
.B(n_1540),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1416),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1419),
.A2(n_1510),
.B1(n_1552),
.B2(n_1542),
.Y(n_1664)
);

O2A1O1Ixp33_ASAP7_75t_L g1665 ( 
.A1(n_1512),
.A2(n_1278),
.B(n_1563),
.C(n_1542),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_SL g1666 ( 
.A1(n_1512),
.A2(n_1563),
.B(n_1542),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_SL g1667 ( 
.A1(n_1512),
.A2(n_1563),
.B(n_1542),
.Y(n_1667)
);

OR2x6_ASAP7_75t_L g1668 ( 
.A(n_1434),
.B(n_1441),
.Y(n_1668)
);

CKINVDCx20_ASAP7_75t_R g1669 ( 
.A(n_1495),
.Y(n_1669)
);

OA21x2_ASAP7_75t_L g1670 ( 
.A1(n_1465),
.A2(n_1467),
.B(n_1454),
.Y(n_1670)
);

AND2x2_ASAP7_75t_SL g1671 ( 
.A(n_1420),
.B(n_1452),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1419),
.A2(n_1510),
.B1(n_1552),
.B2(n_1542),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1419),
.A2(n_1510),
.B1(n_1552),
.B2(n_1542),
.Y(n_1673)
);

O2A1O1Ixp33_ASAP7_75t_L g1674 ( 
.A1(n_1512),
.A2(n_1278),
.B(n_1563),
.C(n_1542),
.Y(n_1674)
);

OR2x6_ASAP7_75t_L g1675 ( 
.A(n_1668),
.B(n_1666),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1614),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1636),
.B(n_1639),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1640),
.B(n_1630),
.Y(n_1678)
);

AOI21xp33_ASAP7_75t_L g1679 ( 
.A1(n_1655),
.A2(n_1674),
.B(n_1665),
.Y(n_1679)
);

BUFx2_ASAP7_75t_L g1680 ( 
.A(n_1635),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1603),
.B(n_1612),
.Y(n_1681)
);

OR2x6_ASAP7_75t_L g1682 ( 
.A(n_1668),
.B(n_1667),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1595),
.B(n_1603),
.Y(n_1683)
);

BUFx6f_ASAP7_75t_L g1684 ( 
.A(n_1635),
.Y(n_1684)
);

BUFx3_ASAP7_75t_L g1685 ( 
.A(n_1617),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1595),
.B(n_1629),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1642),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1612),
.B(n_1629),
.Y(n_1688)
);

OR2x6_ASAP7_75t_L g1689 ( 
.A(n_1668),
.B(n_1575),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1643),
.Y(n_1690)
);

OAI221xp5_ASAP7_75t_L g1691 ( 
.A1(n_1578),
.A2(n_1587),
.B1(n_1576),
.B2(n_1664),
.C(n_1572),
.Y(n_1691)
);

INVx5_ASAP7_75t_L g1692 ( 
.A(n_1641),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1623),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1623),
.Y(n_1694)
);

INVx3_ASAP7_75t_L g1695 ( 
.A(n_1651),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1631),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1631),
.Y(n_1697)
);

OR2x6_ASAP7_75t_L g1698 ( 
.A(n_1659),
.B(n_1582),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1632),
.B(n_1626),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1632),
.B(n_1610),
.Y(n_1700)
);

BUFx2_ASAP7_75t_L g1701 ( 
.A(n_1580),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1634),
.B(n_1670),
.Y(n_1702)
);

OA21x2_ASAP7_75t_L g1703 ( 
.A1(n_1569),
.A2(n_1577),
.B(n_1584),
.Y(n_1703)
);

OAI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1576),
.A2(n_1656),
.B(n_1644),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1670),
.B(n_1591),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1591),
.B(n_1585),
.Y(n_1706)
);

INVx1_ASAP7_75t_SL g1707 ( 
.A(n_1571),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1592),
.Y(n_1708)
);

NOR2x1_ASAP7_75t_L g1709 ( 
.A(n_1624),
.B(n_1621),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1663),
.B(n_1580),
.Y(n_1710)
);

AO21x2_ASAP7_75t_L g1711 ( 
.A1(n_1637),
.A2(n_1577),
.B(n_1584),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1658),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1613),
.Y(n_1713)
);

BUFx2_ASAP7_75t_L g1714 ( 
.A(n_1602),
.Y(n_1714)
);

AO21x2_ASAP7_75t_L g1715 ( 
.A1(n_1658),
.A2(n_1586),
.B(n_1672),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1638),
.Y(n_1716)
);

AO21x2_ASAP7_75t_L g1717 ( 
.A1(n_1572),
.A2(n_1673),
.B(n_1672),
.Y(n_1717)
);

OA21x2_ASAP7_75t_L g1718 ( 
.A1(n_1598),
.A2(n_1601),
.B(n_1664),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1671),
.Y(n_1719)
);

OA21x2_ASAP7_75t_L g1720 ( 
.A1(n_1652),
.A2(n_1673),
.B(n_1660),
.Y(n_1720)
);

OA21x2_ASAP7_75t_L g1721 ( 
.A1(n_1652),
.A2(n_1660),
.B(n_1618),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1568),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1616),
.Y(n_1723)
);

BUFx3_ASAP7_75t_L g1724 ( 
.A(n_1646),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1620),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1573),
.B(n_1645),
.Y(n_1726)
);

OA21x2_ASAP7_75t_L g1727 ( 
.A1(n_1594),
.A2(n_1590),
.B(n_1570),
.Y(n_1727)
);

OA21x2_ASAP7_75t_L g1728 ( 
.A1(n_1590),
.A2(n_1633),
.B(n_1619),
.Y(n_1728)
);

AO21x2_ASAP7_75t_L g1729 ( 
.A1(n_1599),
.A2(n_1605),
.B(n_1604),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1589),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1579),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1687),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1706),
.B(n_1600),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1706),
.B(n_1653),
.Y(n_1734)
);

BUFx3_ASAP7_75t_L g1735 ( 
.A(n_1685),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1683),
.B(n_1654),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1712),
.B(n_1662),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1683),
.B(n_1686),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1706),
.B(n_1650),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1712),
.B(n_1683),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1686),
.B(n_1583),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1712),
.B(n_1648),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1705),
.B(n_1648),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1690),
.Y(n_1744)
);

CKINVDCx14_ASAP7_75t_R g1745 ( 
.A(n_1714),
.Y(n_1745)
);

NOR3xp33_ASAP7_75t_L g1746 ( 
.A(n_1691),
.B(n_1608),
.C(n_1615),
.Y(n_1746)
);

AOI22xp5_ASAP7_75t_SL g1747 ( 
.A1(n_1720),
.A2(n_1669),
.B1(n_1596),
.B2(n_1661),
.Y(n_1747)
);

INVx8_ASAP7_75t_L g1748 ( 
.A(n_1675),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1691),
.A2(n_1593),
.B1(n_1649),
.B2(n_1588),
.Y(n_1749)
);

INVx2_ASAP7_75t_SL g1750 ( 
.A(n_1692),
.Y(n_1750)
);

BUFx2_ASAP7_75t_L g1751 ( 
.A(n_1676),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1704),
.A2(n_1609),
.B1(n_1657),
.B2(n_1581),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1688),
.B(n_1611),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1700),
.B(n_1607),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1688),
.B(n_1574),
.Y(n_1755)
);

INVx3_ASAP7_75t_L g1756 ( 
.A(n_1695),
.Y(n_1756)
);

AOI222xp33_ASAP7_75t_L g1757 ( 
.A1(n_1704),
.A2(n_1647),
.B1(n_1622),
.B2(n_1628),
.C1(n_1627),
.C2(n_1625),
.Y(n_1757)
);

NAND4xp25_ASAP7_75t_L g1758 ( 
.A(n_1679),
.B(n_1597),
.C(n_1606),
.D(n_1713),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1699),
.B(n_1606),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1688),
.B(n_1681),
.Y(n_1760)
);

BUFx3_ASAP7_75t_L g1761 ( 
.A(n_1684),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1699),
.B(n_1678),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1703),
.B(n_1711),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1699),
.B(n_1678),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1676),
.Y(n_1765)
);

INVx3_ASAP7_75t_L g1766 ( 
.A(n_1695),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1678),
.B(n_1677),
.Y(n_1767)
);

AOI222xp33_ASAP7_75t_L g1768 ( 
.A1(n_1730),
.A2(n_1679),
.B1(n_1716),
.B2(n_1717),
.C1(n_1713),
.C2(n_1719),
.Y(n_1768)
);

BUFx2_ASAP7_75t_L g1769 ( 
.A(n_1710),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1703),
.B(n_1711),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1677),
.B(n_1702),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1733),
.B(n_1722),
.Y(n_1772)
);

INVx5_ASAP7_75t_L g1773 ( 
.A(n_1750),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1732),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1732),
.Y(n_1775)
);

BUFx3_ASAP7_75t_L g1776 ( 
.A(n_1735),
.Y(n_1776)
);

OR2x6_ASAP7_75t_L g1777 ( 
.A(n_1748),
.B(n_1675),
.Y(n_1777)
);

AOI31xp33_ASAP7_75t_L g1778 ( 
.A1(n_1747),
.A2(n_1709),
.A3(n_1730),
.B(n_1719),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1765),
.Y(n_1779)
);

HB1xp67_ASAP7_75t_L g1780 ( 
.A(n_1765),
.Y(n_1780)
);

AO21x2_ASAP7_75t_L g1781 ( 
.A1(n_1763),
.A2(n_1708),
.B(n_1693),
.Y(n_1781)
);

BUFx2_ASAP7_75t_L g1782 ( 
.A(n_1751),
.Y(n_1782)
);

NOR2x1_ASAP7_75t_L g1783 ( 
.A(n_1763),
.B(n_1709),
.Y(n_1783)
);

INVxp67_ASAP7_75t_L g1784 ( 
.A(n_1755),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_R g1785 ( 
.A(n_1745),
.B(n_1724),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_R g1786 ( 
.A(n_1749),
.B(n_1724),
.Y(n_1786)
);

OAI31xp33_ASAP7_75t_L g1787 ( 
.A1(n_1746),
.A2(n_1758),
.A3(n_1701),
.B(n_1723),
.Y(n_1787)
);

INVx5_ASAP7_75t_L g1788 ( 
.A(n_1750),
.Y(n_1788)
);

BUFx2_ASAP7_75t_L g1789 ( 
.A(n_1751),
.Y(n_1789)
);

AOI22xp33_ASAP7_75t_SL g1790 ( 
.A1(n_1747),
.A2(n_1717),
.B1(n_1720),
.B2(n_1721),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1746),
.A2(n_1717),
.B1(n_1720),
.B2(n_1721),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1758),
.A2(n_1717),
.B1(n_1720),
.B2(n_1721),
.Y(n_1792)
);

AND2x2_ASAP7_75t_SL g1793 ( 
.A(n_1753),
.B(n_1701),
.Y(n_1793)
);

NOR4xp25_ASAP7_75t_SL g1794 ( 
.A(n_1769),
.B(n_1723),
.C(n_1680),
.D(n_1725),
.Y(n_1794)
);

XNOR2xp5_ASAP7_75t_L g1795 ( 
.A(n_1752),
.B(n_1726),
.Y(n_1795)
);

NOR2x1_ASAP7_75t_SL g1796 ( 
.A(n_1753),
.B(n_1689),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1760),
.B(n_1739),
.Y(n_1797)
);

OAI221xp5_ASAP7_75t_SL g1798 ( 
.A1(n_1768),
.A2(n_1698),
.B1(n_1675),
.B2(n_1682),
.C(n_1719),
.Y(n_1798)
);

NAND2xp33_ASAP7_75t_R g1799 ( 
.A(n_1755),
.B(n_1721),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1768),
.A2(n_1715),
.B1(n_1675),
.B2(n_1682),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_L g1801 ( 
.A(n_1737),
.B(n_1731),
.Y(n_1801)
);

OAI211xp5_ASAP7_75t_L g1802 ( 
.A1(n_1770),
.A2(n_1718),
.B(n_1757),
.C(n_1742),
.Y(n_1802)
);

OAI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1742),
.A2(n_1675),
.B1(n_1682),
.B2(n_1718),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1760),
.B(n_1681),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_SL g1805 ( 
.A1(n_1743),
.A2(n_1729),
.B1(n_1715),
.B2(n_1675),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1762),
.B(n_1714),
.Y(n_1806)
);

BUFx6f_ASAP7_75t_L g1807 ( 
.A(n_1761),
.Y(n_1807)
);

AOI22xp33_ASAP7_75t_L g1808 ( 
.A1(n_1743),
.A2(n_1715),
.B1(n_1682),
.B2(n_1729),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1739),
.B(n_1681),
.Y(n_1809)
);

OA21x2_ASAP7_75t_L g1810 ( 
.A1(n_1744),
.A2(n_1694),
.B(n_1693),
.Y(n_1810)
);

NAND2xp33_ASAP7_75t_R g1811 ( 
.A(n_1759),
.B(n_1728),
.Y(n_1811)
);

NAND4xp75_ASAP7_75t_L g1812 ( 
.A(n_1787),
.B(n_1727),
.C(n_1718),
.D(n_1703),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1774),
.Y(n_1813)
);

HB1xp67_ASAP7_75t_L g1814 ( 
.A(n_1779),
.Y(n_1814)
);

INVxp67_ASAP7_75t_SL g1815 ( 
.A(n_1783),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1774),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1810),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1797),
.B(n_1734),
.Y(n_1818)
);

INVx1_ASAP7_75t_SL g1819 ( 
.A(n_1782),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1775),
.Y(n_1820)
);

INVxp67_ASAP7_75t_SL g1821 ( 
.A(n_1783),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1775),
.Y(n_1822)
);

OAI21x1_ASAP7_75t_L g1823 ( 
.A1(n_1803),
.A2(n_1766),
.B(n_1756),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1801),
.B(n_1707),
.Y(n_1824)
);

BUFx3_ASAP7_75t_L g1825 ( 
.A(n_1776),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1780),
.Y(n_1826)
);

AND2x4_ASAP7_75t_L g1827 ( 
.A(n_1773),
.B(n_1788),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1797),
.B(n_1734),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1781),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1773),
.B(n_1761),
.Y(n_1830)
);

INVx1_ASAP7_75t_SL g1831 ( 
.A(n_1782),
.Y(n_1831)
);

OAI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1805),
.A2(n_1790),
.B(n_1778),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1781),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1781),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1793),
.B(n_1762),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1793),
.B(n_1762),
.Y(n_1836)
);

HB1xp67_ASAP7_75t_L g1837 ( 
.A(n_1789),
.Y(n_1837)
);

INVx1_ASAP7_75t_SL g1838 ( 
.A(n_1789),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1784),
.B(n_1736),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_SL g1840 ( 
.A(n_1785),
.B(n_1754),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1804),
.B(n_1738),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1806),
.B(n_1764),
.Y(n_1842)
);

OA21x2_ASAP7_75t_L g1843 ( 
.A1(n_1802),
.A2(n_1697),
.B(n_1696),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1804),
.B(n_1738),
.Y(n_1844)
);

BUFx3_ASAP7_75t_L g1845 ( 
.A(n_1776),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1806),
.B(n_1764),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1809),
.B(n_1740),
.Y(n_1847)
);

INVxp67_ASAP7_75t_L g1848 ( 
.A(n_1799),
.Y(n_1848)
);

CKINVDCx20_ASAP7_75t_R g1849 ( 
.A(n_1786),
.Y(n_1849)
);

AND2x4_ASAP7_75t_SL g1850 ( 
.A(n_1777),
.B(n_1682),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1807),
.B(n_1764),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1817),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1835),
.B(n_1796),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1848),
.B(n_1743),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1813),
.Y(n_1855)
);

INVxp67_ASAP7_75t_L g1856 ( 
.A(n_1837),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1817),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1841),
.B(n_1772),
.Y(n_1858)
);

INVx1_ASAP7_75t_SL g1859 ( 
.A(n_1819),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1835),
.B(n_1836),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1836),
.B(n_1796),
.Y(n_1861)
);

AND2x4_ASAP7_75t_L g1862 ( 
.A(n_1827),
.B(n_1773),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1813),
.Y(n_1863)
);

INVx2_ASAP7_75t_SL g1864 ( 
.A(n_1827),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1851),
.B(n_1807),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1816),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1817),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1814),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1851),
.B(n_1842),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1832),
.A2(n_1798),
.B(n_1800),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1842),
.B(n_1807),
.Y(n_1871)
);

AOI21xp33_ASAP7_75t_L g1872 ( 
.A1(n_1832),
.A2(n_1811),
.B(n_1757),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1846),
.B(n_1830),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1816),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1846),
.B(n_1807),
.Y(n_1875)
);

INVxp67_ASAP7_75t_SL g1876 ( 
.A(n_1829),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1849),
.B(n_1707),
.Y(n_1877)
);

INVxp67_ASAP7_75t_L g1878 ( 
.A(n_1815),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1830),
.B(n_1807),
.Y(n_1879)
);

INVxp67_ASAP7_75t_L g1880 ( 
.A(n_1821),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1830),
.B(n_1827),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1820),
.Y(n_1882)
);

AND2x4_ASAP7_75t_L g1883 ( 
.A(n_1827),
.B(n_1773),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1820),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_L g1885 ( 
.A(n_1824),
.B(n_1726),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1822),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1830),
.B(n_1771),
.Y(n_1887)
);

INVx1_ASAP7_75t_SL g1888 ( 
.A(n_1819),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1822),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1831),
.B(n_1736),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1825),
.B(n_1771),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1825),
.B(n_1771),
.Y(n_1892)
);

INVx2_ASAP7_75t_SL g1893 ( 
.A(n_1825),
.Y(n_1893)
);

INVx1_ASAP7_75t_SL g1894 ( 
.A(n_1831),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1845),
.B(n_1769),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_SL g1896 ( 
.A(n_1840),
.B(n_1808),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1845),
.B(n_1767),
.Y(n_1897)
);

NOR2xp33_ASAP7_75t_L g1898 ( 
.A(n_1845),
.B(n_1726),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1838),
.B(n_1741),
.Y(n_1899)
);

INVx1_ASAP7_75t_SL g1900 ( 
.A(n_1826),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1823),
.B(n_1767),
.Y(n_1901)
);

INVx2_ASAP7_75t_SL g1902 ( 
.A(n_1881),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1855),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1900),
.B(n_1868),
.Y(n_1904)
);

INVx1_ASAP7_75t_SL g1905 ( 
.A(n_1900),
.Y(n_1905)
);

NAND2x1p5_ASAP7_75t_L g1906 ( 
.A(n_1859),
.B(n_1773),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1854),
.B(n_1844),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1854),
.B(n_1818),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1855),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1860),
.B(n_1823),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1852),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1863),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1863),
.Y(n_1913)
);

NAND3xp33_ASAP7_75t_L g1914 ( 
.A(n_1870),
.B(n_1843),
.C(n_1792),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1866),
.Y(n_1915)
);

AND2x4_ASAP7_75t_L g1916 ( 
.A(n_1864),
.B(n_1850),
.Y(n_1916)
);

HB1xp67_ASAP7_75t_L g1917 ( 
.A(n_1859),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1866),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1874),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1898),
.B(n_1839),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1888),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1874),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1882),
.Y(n_1923)
);

OR2x2_ASAP7_75t_L g1924 ( 
.A(n_1858),
.B(n_1818),
.Y(n_1924)
);

OR2x2_ASAP7_75t_L g1925 ( 
.A(n_1858),
.B(n_1828),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1882),
.Y(n_1926)
);

HB1xp67_ASAP7_75t_L g1927 ( 
.A(n_1888),
.Y(n_1927)
);

AOI21xp5_ASAP7_75t_L g1928 ( 
.A1(n_1872),
.A2(n_1843),
.B(n_1791),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1852),
.Y(n_1929)
);

OAI22xp5_ASAP7_75t_L g1930 ( 
.A1(n_1870),
.A2(n_1812),
.B1(n_1794),
.B2(n_1777),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1860),
.B(n_1850),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1893),
.B(n_1795),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1893),
.B(n_1795),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1894),
.B(n_1828),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1881),
.B(n_1850),
.Y(n_1935)
);

OR2x2_ASAP7_75t_L g1936 ( 
.A(n_1894),
.B(n_1847),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1884),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1884),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1886),
.Y(n_1939)
);

AOI21xp5_ASAP7_75t_L g1940 ( 
.A1(n_1872),
.A2(n_1843),
.B(n_1729),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1886),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1852),
.Y(n_1942)
);

INVx1_ASAP7_75t_SL g1943 ( 
.A(n_1905),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1906),
.Y(n_1944)
);

INVxp67_ASAP7_75t_L g1945 ( 
.A(n_1917),
.Y(n_1945)
);

INVx1_ASAP7_75t_SL g1946 ( 
.A(n_1917),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1906),
.Y(n_1947)
);

OAI221xp5_ASAP7_75t_L g1948 ( 
.A1(n_1914),
.A2(n_1896),
.B1(n_1880),
.B2(n_1878),
.C(n_1856),
.Y(n_1948)
);

INVxp67_ASAP7_75t_L g1949 ( 
.A(n_1921),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1921),
.B(n_1856),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1927),
.B(n_1897),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1927),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_L g1953 ( 
.A(n_1904),
.B(n_1877),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1903),
.Y(n_1954)
);

NOR2xp33_ASAP7_75t_L g1955 ( 
.A(n_1932),
.B(n_1885),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1902),
.Y(n_1956)
);

AOI21xp5_ASAP7_75t_L g1957 ( 
.A1(n_1928),
.A2(n_1880),
.B(n_1878),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1909),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1902),
.Y(n_1959)
);

OAI22xp5_ASAP7_75t_L g1960 ( 
.A1(n_1930),
.A2(n_1812),
.B1(n_1861),
.B2(n_1853),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1935),
.B(n_1879),
.Y(n_1961)
);

NAND2x1_ASAP7_75t_SL g1962 ( 
.A(n_1916),
.B(n_1879),
.Y(n_1962)
);

INVx1_ASAP7_75t_SL g1963 ( 
.A(n_1936),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1933),
.B(n_1897),
.Y(n_1964)
);

NOR2xp67_ASAP7_75t_SL g1965 ( 
.A(n_1940),
.B(n_1864),
.Y(n_1965)
);

NOR2x1p5_ASAP7_75t_L g1966 ( 
.A(n_1934),
.B(n_1936),
.Y(n_1966)
);

CKINVDCx16_ASAP7_75t_R g1967 ( 
.A(n_1931),
.Y(n_1967)
);

OAI21x1_ASAP7_75t_L g1968 ( 
.A1(n_1911),
.A2(n_1867),
.B(n_1857),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1912),
.Y(n_1969)
);

CKINVDCx16_ASAP7_75t_R g1970 ( 
.A(n_1931),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1913),
.Y(n_1971)
);

BUFx2_ASAP7_75t_L g1972 ( 
.A(n_1916),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1935),
.B(n_1873),
.Y(n_1973)
);

OAI211xp5_ASAP7_75t_SL g1974 ( 
.A1(n_1948),
.A2(n_1908),
.B(n_1907),
.C(n_1915),
.Y(n_1974)
);

OAI21xp5_ASAP7_75t_L g1975 ( 
.A1(n_1960),
.A2(n_1916),
.B(n_1843),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1950),
.Y(n_1976)
);

AOI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1967),
.A2(n_1853),
.B1(n_1861),
.B2(n_1865),
.Y(n_1977)
);

NAND2x1p5_ASAP7_75t_L g1978 ( 
.A(n_1943),
.B(n_1862),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1950),
.Y(n_1979)
);

OAI21xp5_ASAP7_75t_SL g1980 ( 
.A1(n_1953),
.A2(n_1910),
.B(n_1883),
.Y(n_1980)
);

OAI22xp33_ASAP7_75t_L g1981 ( 
.A1(n_1970),
.A2(n_1908),
.B1(n_1920),
.B2(n_1924),
.Y(n_1981)
);

OAI21xp33_ASAP7_75t_L g1982 ( 
.A1(n_1962),
.A2(n_1910),
.B(n_1925),
.Y(n_1982)
);

OAI221xp5_ASAP7_75t_L g1983 ( 
.A1(n_1957),
.A2(n_1938),
.B1(n_1937),
.B2(n_1926),
.C(n_1923),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1946),
.B(n_1869),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1952),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1962),
.Y(n_1986)
);

OR2x2_ASAP7_75t_L g1987 ( 
.A(n_1963),
.B(n_1951),
.Y(n_1987)
);

O2A1O1Ixp33_ASAP7_75t_L g1988 ( 
.A1(n_1945),
.A2(n_1919),
.B(n_1922),
.C(n_1918),
.Y(n_1988)
);

NOR2x1_ASAP7_75t_L g1989 ( 
.A(n_1952),
.B(n_1939),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1973),
.B(n_1961),
.Y(n_1990)
);

NAND2xp33_ASAP7_75t_L g1991 ( 
.A(n_1966),
.B(n_1895),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1949),
.Y(n_1992)
);

CKINVDCx16_ASAP7_75t_R g1993 ( 
.A(n_1972),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1972),
.B(n_1862),
.Y(n_1994)
);

AOI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1955),
.A2(n_1941),
.B(n_1883),
.Y(n_1995)
);

OAI22xp5_ASAP7_75t_L g1996 ( 
.A1(n_1993),
.A2(n_1964),
.B1(n_1959),
.B2(n_1956),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1989),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1976),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_L g1999 ( 
.A(n_1992),
.B(n_1961),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1979),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1985),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1990),
.B(n_1973),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1984),
.Y(n_2003)
);

OR2x2_ASAP7_75t_L g2004 ( 
.A(n_1987),
.B(n_1956),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1981),
.B(n_1959),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1978),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1978),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1988),
.B(n_1954),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1994),
.Y(n_2009)
);

NAND3xp33_ASAP7_75t_L g2010 ( 
.A(n_1997),
.B(n_1991),
.C(n_1986),
.Y(n_2010)
);

AOI21xp33_ASAP7_75t_L g2011 ( 
.A1(n_1996),
.A2(n_2005),
.B(n_2006),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_2002),
.B(n_1995),
.Y(n_2012)
);

OAI211xp5_ASAP7_75t_SL g2013 ( 
.A1(n_2008),
.A2(n_2009),
.B(n_2003),
.C(n_1975),
.Y(n_2013)
);

AOI211xp5_ASAP7_75t_L g2014 ( 
.A1(n_1996),
.A2(n_1982),
.B(n_2008),
.C(n_1983),
.Y(n_2014)
);

AOI322xp5_ASAP7_75t_L g2015 ( 
.A1(n_1999),
.A2(n_1977),
.A3(n_1969),
.B1(n_1971),
.B2(n_1958),
.C1(n_1947),
.C2(n_1944),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_2004),
.Y(n_2016)
);

NOR3xp33_ASAP7_75t_L g2017 ( 
.A(n_2007),
.B(n_2000),
.C(n_1998),
.Y(n_2017)
);

NOR2x1_ASAP7_75t_L g2018 ( 
.A(n_2001),
.B(n_1980),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_2002),
.B(n_1980),
.Y(n_2019)
);

OAI22xp33_ASAP7_75t_L g2020 ( 
.A1(n_1997),
.A2(n_1947),
.B1(n_1944),
.B2(n_1788),
.Y(n_2020)
);

OAI22xp5_ASAP7_75t_L g2021 ( 
.A1(n_2005),
.A2(n_1883),
.B1(n_1862),
.B2(n_1890),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_2016),
.Y(n_2022)
);

AOI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_2013),
.A2(n_1974),
.B(n_1969),
.Y(n_2023)
);

AOI221x1_ASAP7_75t_L g2024 ( 
.A1(n_2011),
.A2(n_1971),
.B1(n_1958),
.B2(n_1929),
.C(n_1911),
.Y(n_2024)
);

AOI22xp5_ASAP7_75t_L g2025 ( 
.A1(n_2014),
.A2(n_1965),
.B1(n_1862),
.B2(n_1883),
.Y(n_2025)
);

OAI211xp5_ASAP7_75t_L g2026 ( 
.A1(n_2018),
.A2(n_1965),
.B(n_1942),
.C(n_1929),
.Y(n_2026)
);

AOI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_2012),
.A2(n_1968),
.B(n_1942),
.Y(n_2027)
);

INVx1_ASAP7_75t_SL g2028 ( 
.A(n_2019),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_2022),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_2028),
.B(n_2017),
.Y(n_2030)
);

CKINVDCx14_ASAP7_75t_R g2031 ( 
.A(n_2025),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_2024),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_2023),
.B(n_2015),
.Y(n_2033)
);

NOR2xp33_ASAP7_75t_L g2034 ( 
.A(n_2026),
.B(n_2010),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_2027),
.Y(n_2035)
);

NOR2xp33_ASAP7_75t_L g2036 ( 
.A(n_2028),
.B(n_2021),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_2034),
.B(n_2020),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_2030),
.B(n_2031),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_2029),
.Y(n_2039)
);

AOI211xp5_ASAP7_75t_L g2040 ( 
.A1(n_2033),
.A2(n_1968),
.B(n_1901),
.C(n_1876),
.Y(n_2040)
);

AOI211xp5_ASAP7_75t_L g2041 ( 
.A1(n_2033),
.A2(n_2036),
.B(n_2032),
.C(n_2035),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_2030),
.Y(n_2042)
);

NAND3xp33_ASAP7_75t_L g2043 ( 
.A(n_2041),
.B(n_1876),
.C(n_1867),
.Y(n_2043)
);

NAND3xp33_ASAP7_75t_L g2044 ( 
.A(n_2037),
.B(n_1867),
.C(n_1857),
.Y(n_2044)
);

AOI322xp5_ASAP7_75t_L g2045 ( 
.A1(n_2038),
.A2(n_1857),
.A3(n_1895),
.B1(n_1865),
.B2(n_1901),
.C1(n_1829),
.C2(n_1834),
.Y(n_2045)
);

NOR3xp33_ASAP7_75t_L g2046 ( 
.A(n_2042),
.B(n_1873),
.C(n_1890),
.Y(n_2046)
);

INVxp33_ASAP7_75t_SL g2047 ( 
.A(n_2043),
.Y(n_2047)
);

OAI22xp5_ASAP7_75t_L g2048 ( 
.A1(n_2044),
.A2(n_2040),
.B1(n_2039),
.B2(n_2046),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_2048),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_2047),
.B(n_2045),
.Y(n_2050)
);

AOI222xp33_ASAP7_75t_L g2051 ( 
.A1(n_2050),
.A2(n_1834),
.B1(n_1833),
.B2(n_1829),
.C1(n_1889),
.C2(n_1871),
.Y(n_2051)
);

AO21x2_ASAP7_75t_L g2052 ( 
.A1(n_2049),
.A2(n_1889),
.B(n_1834),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_2052),
.Y(n_2053)
);

OA21x2_ASAP7_75t_L g2054 ( 
.A1(n_2051),
.A2(n_1833),
.B(n_1869),
.Y(n_2054)
);

NAND2xp33_ASAP7_75t_SL g2055 ( 
.A(n_2053),
.B(n_1871),
.Y(n_2055)
);

INVxp67_ASAP7_75t_L g2056 ( 
.A(n_2054),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2055),
.Y(n_2057)
);

OAI21xp5_ASAP7_75t_L g2058 ( 
.A1(n_2057),
.A2(n_2056),
.B(n_2054),
.Y(n_2058)
);

AOI21xp5_ASAP7_75t_L g2059 ( 
.A1(n_2058),
.A2(n_2054),
.B(n_1899),
.Y(n_2059)
);

AOI22xp33_ASAP7_75t_L g2060 ( 
.A1(n_2059),
.A2(n_1833),
.B1(n_1875),
.B2(n_1887),
.Y(n_2060)
);

AOI22xp33_ASAP7_75t_L g2061 ( 
.A1(n_2060),
.A2(n_1875),
.B1(n_1887),
.B2(n_1891),
.Y(n_2061)
);

AOI211xp5_ASAP7_75t_L g2062 ( 
.A1(n_2061),
.A2(n_1899),
.B(n_1891),
.C(n_1892),
.Y(n_2062)
);


endmodule