module real_aes_8465_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_119;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AOI22xp33_ASAP7_75t_L g175 ( .A1(n_0), .A2(n_67), .B1(n_176), .B2(n_180), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_1), .Y(n_105) );
A2O1A1Ixp33_ASAP7_75t_L g269 ( .A1(n_2), .A2(n_229), .B(n_233), .C(n_270), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_3), .A2(n_224), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_4), .B(n_260), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g147 ( .A1(n_5), .A2(n_54), .B1(n_148), .B2(n_154), .Y(n_147) );
INVx1_ASAP7_75t_L g209 ( .A(n_6), .Y(n_209) );
AND2x6_ASAP7_75t_L g229 ( .A(n_6), .B(n_207), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_6), .B(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g240 ( .A(n_7), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_8), .B(n_238), .Y(n_274) );
AO22x2_ASAP7_75t_L g94 ( .A1(n_9), .A2(n_26), .B1(n_95), .B2(n_96), .Y(n_94) );
INVx1_ASAP7_75t_L g222 ( .A(n_10), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_11), .A2(n_241), .B(n_255), .C(n_258), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_12), .B(n_260), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_13), .A2(n_85), .B1(n_184), .B2(n_536), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_13), .Y(n_536) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_14), .A2(n_28), .B1(n_95), .B2(n_99), .Y(n_98) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_15), .B(n_365), .Y(n_364) );
A2O1A1Ixp33_ASAP7_75t_L g283 ( .A1(n_16), .A2(n_284), .B(n_285), .C(n_287), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_17), .B(n_238), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_18), .B(n_238), .Y(n_298) );
CKINVDCx16_ASAP7_75t_R g308 ( .A(n_19), .Y(n_308) );
INVx1_ASAP7_75t_L g296 ( .A(n_20), .Y(n_296) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_21), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_22), .Y(n_267) );
INVx1_ASAP7_75t_L g361 ( .A(n_23), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_24), .A2(n_188), .B1(n_189), .B2(n_192), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_24), .Y(n_188) );
INVx2_ASAP7_75t_L g227 ( .A(n_25), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g277 ( .A(n_27), .Y(n_277) );
OAI221xp5_ASAP7_75t_L g200 ( .A1(n_28), .A2(n_43), .B1(n_53), .B2(n_201), .C(n_202), .Y(n_200) );
INVxp67_ASAP7_75t_L g203 ( .A(n_28), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g321 ( .A1(n_29), .A2(n_284), .B(n_322), .C(n_323), .Y(n_321) );
INVxp67_ASAP7_75t_L g362 ( .A(n_30), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_30), .A2(n_85), .B1(n_184), .B2(n_362), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_31), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g294 ( .A1(n_32), .A2(n_233), .B(n_295), .C(n_301), .Y(n_294) );
CKINVDCx14_ASAP7_75t_R g320 ( .A(n_33), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_34), .B(n_128), .Y(n_127) );
AOI22xp33_ASAP7_75t_L g158 ( .A1(n_35), .A2(n_55), .B1(n_159), .B2(n_163), .Y(n_158) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_36), .A2(n_237), .B(n_239), .C(n_242), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g303 ( .A(n_37), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g168 ( .A1(n_38), .A2(n_73), .B1(n_169), .B2(n_172), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g358 ( .A(n_39), .Y(n_358) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_40), .Y(n_126) );
INVx1_ASAP7_75t_L g282 ( .A(n_41), .Y(n_282) );
CKINVDCx20_ASAP7_75t_R g88 ( .A(n_42), .Y(n_88) );
AO22x2_ASAP7_75t_L g104 ( .A1(n_43), .A2(n_64), .B1(n_95), .B2(n_99), .Y(n_104) );
INVxp67_ASAP7_75t_L g204 ( .A(n_43), .Y(n_204) );
CKINVDCx14_ASAP7_75t_R g231 ( .A(n_44), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_45), .Y(n_133) );
INVx1_ASAP7_75t_L g207 ( .A(n_46), .Y(n_207) );
INVx1_ASAP7_75t_L g221 ( .A(n_47), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g82 ( .A1(n_48), .A2(n_63), .B1(n_83), .B2(n_84), .Y(n_82) );
INVx1_ASAP7_75t_SL g83 ( .A(n_48), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_49), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_50), .B(n_260), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_51), .Y(n_118) );
INVx1_ASAP7_75t_L g311 ( .A(n_52), .Y(n_311) );
AO22x2_ASAP7_75t_L g102 ( .A1(n_53), .A2(n_72), .B1(n_95), .B2(n_96), .Y(n_102) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_56), .A2(n_224), .B(n_230), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g315 ( .A(n_57), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_58), .A2(n_224), .B(n_252), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g355 ( .A1(n_59), .A2(n_356), .B(n_357), .Y(n_355) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_59), .Y(n_534) );
INVx1_ASAP7_75t_L g253 ( .A(n_60), .Y(n_253) );
CKINVDCx16_ASAP7_75t_R g293 ( .A(n_61), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_62), .A2(n_224), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g84 ( .A(n_63), .Y(n_84) );
INVx2_ASAP7_75t_L g219 ( .A(n_65), .Y(n_219) );
INVx1_ASAP7_75t_L g271 ( .A(n_66), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_68), .A2(n_69), .B1(n_190), .B2(n_191), .Y(n_189) );
CKINVDCx14_ASAP7_75t_R g191 ( .A(n_68), .Y(n_191) );
INVx1_ASAP7_75t_L g190 ( .A(n_69), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g309 ( .A1(n_70), .A2(n_233), .B(n_310), .C(n_313), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g193 ( .A1(n_71), .A2(n_76), .B1(n_194), .B2(n_195), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_71), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_74), .B(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g95 ( .A(n_75), .Y(n_95) );
INVx1_ASAP7_75t_L g97 ( .A(n_75), .Y(n_97) );
INVx1_ASAP7_75t_L g195 ( .A(n_76), .Y(n_195) );
INVx2_ASAP7_75t_L g286 ( .A(n_77), .Y(n_286) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_197), .B1(n_210), .B2(n_521), .C(n_524), .Y(n_78) );
XNOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_185), .Y(n_79) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_81), .A2(n_82), .B1(n_85), .B2(n_184), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_83), .B(n_284), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_84), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g184 ( .A(n_85), .Y(n_184) );
AND2x2_ASAP7_75t_L g85 ( .A(n_86), .B(n_145), .Y(n_85) );
NOR3xp33_ASAP7_75t_L g86 ( .A(n_87), .B(n_111), .C(n_132), .Y(n_86) );
OAI22xp5_ASAP7_75t_L g87 ( .A1(n_88), .A2(n_89), .B1(n_105), .B2(n_106), .Y(n_87) );
INVx2_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
OR2x2_ASAP7_75t_L g91 ( .A(n_92), .B(n_100), .Y(n_91) );
INVx2_ASAP7_75t_L g162 ( .A(n_92), .Y(n_162) );
OR2x2_ASAP7_75t_L g92 ( .A(n_93), .B(n_98), .Y(n_92) );
AND2x2_ASAP7_75t_L g110 ( .A(n_93), .B(n_98), .Y(n_110) );
AND2x2_ASAP7_75t_L g153 ( .A(n_93), .B(n_124), .Y(n_153) );
INVx2_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
AND2x2_ASAP7_75t_L g115 ( .A(n_94), .B(n_98), .Y(n_115) );
AND2x2_ASAP7_75t_L g125 ( .A(n_94), .B(n_104), .Y(n_125) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx1_ASAP7_75t_L g99 ( .A(n_97), .Y(n_99) );
INVx2_ASAP7_75t_L g124 ( .A(n_98), .Y(n_124) );
INVx1_ASAP7_75t_L g183 ( .A(n_98), .Y(n_183) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
NAND2x1p5_ASAP7_75t_L g109 ( .A(n_101), .B(n_110), .Y(n_109) );
AND2x4_ASAP7_75t_L g174 ( .A(n_101), .B(n_153), .Y(n_174) );
AND2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_103), .Y(n_101) );
INVx1_ASAP7_75t_L g117 ( .A(n_102), .Y(n_117) );
INVx1_ASAP7_75t_L g123 ( .A(n_102), .Y(n_123) );
INVx1_ASAP7_75t_L g144 ( .A(n_102), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_102), .B(n_104), .Y(n_157) );
AND2x2_ASAP7_75t_L g116 ( .A(n_103), .B(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g152 ( .A(n_104), .B(n_144), .Y(n_152) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x4_ASAP7_75t_L g166 ( .A(n_110), .B(n_116), .Y(n_166) );
AND2x2_ASAP7_75t_L g179 ( .A(n_110), .B(n_152), .Y(n_179) );
OAI221xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_118), .B1(n_119), .B2(n_126), .C(n_127), .Y(n_111) );
INVx2_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x6_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
INVx1_ASAP7_75t_L g141 ( .A(n_115), .Y(n_141) );
AND2x6_ASAP7_75t_L g161 ( .A(n_116), .B(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g171 ( .A(n_116), .B(n_153), .Y(n_171) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx4f_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_125), .Y(n_121) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
INVx1_ASAP7_75t_L g131 ( .A(n_123), .Y(n_131) );
INVx1_ASAP7_75t_L g136 ( .A(n_124), .Y(n_136) );
AND2x4_ASAP7_75t_L g130 ( .A(n_125), .B(n_131), .Y(n_130) );
NAND2x1p5_ASAP7_75t_L g135 ( .A(n_125), .B(n_136), .Y(n_135) );
BUFx4f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OAI22xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_134), .B1(n_137), .B2(n_138), .Y(n_132) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
CKINVDCx16_ASAP7_75t_R g139 ( .A(n_140), .Y(n_139) );
OR2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_146), .B(n_167), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_158), .Y(n_146) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
AND2x4_ASAP7_75t_L g155 ( .A(n_153), .B(n_156), .Y(n_155) );
BUFx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
OR2x6_ASAP7_75t_L g182 ( .A(n_157), .B(n_183), .Y(n_182) );
INVx4_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx11_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_168), .B(n_175), .Y(n_167) );
BUFx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
BUFx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx5_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx8_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
BUFx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx6_ASAP7_75t_SL g181 ( .A(n_182), .Y(n_181) );
OAI22xp5_ASAP7_75t_SL g185 ( .A1(n_186), .A2(n_187), .B1(n_193), .B2(n_196), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_187), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_189), .Y(n_192) );
INVx1_ASAP7_75t_L g196 ( .A(n_193), .Y(n_196) );
CKINVDCx16_ASAP7_75t_R g197 ( .A(n_198), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_199), .Y(n_198) );
AND3x1_ASAP7_75t_SL g199 ( .A(n_200), .B(n_205), .C(n_208), .Y(n_199) );
INVxp67_ASAP7_75t_L g529 ( .A(n_200), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
INVx1_ASAP7_75t_SL g531 ( .A(n_205), .Y(n_531) );
OA21x2_ASAP7_75t_L g532 ( .A1(n_205), .A2(n_225), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g538 ( .A(n_205), .Y(n_538) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_206), .B(n_209), .Y(n_533) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
OR2x2_ASAP7_75t_SL g537 ( .A(n_208), .B(n_538), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
OR2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_451), .Y(n_212) );
NAND5xp2_ASAP7_75t_L g213 ( .A(n_214), .B(n_366), .C(n_398), .D(n_415), .E(n_438), .Y(n_213) );
AOI221xp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_290), .B1(n_326), .B2(n_330), .C(n_334), .Y(n_214) );
INVx1_ASAP7_75t_L g478 ( .A(n_215), .Y(n_478) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_262), .Y(n_215) );
AND3x2_ASAP7_75t_L g453 ( .A(n_216), .B(n_264), .C(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_248), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_217), .B(n_332), .Y(n_331) );
BUFx3_ASAP7_75t_L g341 ( .A(n_217), .Y(n_341) );
AND2x2_ASAP7_75t_L g345 ( .A(n_217), .B(n_278), .Y(n_345) );
INVx2_ASAP7_75t_L g375 ( .A(n_217), .Y(n_375) );
OR2x2_ASAP7_75t_L g386 ( .A(n_217), .B(n_279), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_217), .B(n_263), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_217), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g465 ( .A(n_217), .B(n_279), .Y(n_465) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_223), .B(n_245), .Y(n_217) );
INVx1_ASAP7_75t_L g265 ( .A(n_218), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_L g292 ( .A1(n_218), .A2(n_268), .B(n_293), .C(n_294), .Y(n_292) );
INVx2_ASAP7_75t_L g316 ( .A(n_218), .Y(n_316) );
AND2x2_ASAP7_75t_SL g218 ( .A(n_219), .B(n_220), .Y(n_218) );
AND2x2_ASAP7_75t_L g247 ( .A(n_219), .B(n_220), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
BUFx2_ASAP7_75t_L g356 ( .A(n_224), .Y(n_356) );
AND2x4_ASAP7_75t_L g224 ( .A(n_225), .B(n_229), .Y(n_224) );
NAND2x1p5_ASAP7_75t_L g268 ( .A(n_225), .B(n_229), .Y(n_268) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_228), .Y(n_225) );
INVx1_ASAP7_75t_L g300 ( .A(n_226), .Y(n_300) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g234 ( .A(n_227), .Y(n_234) );
INVx1_ASAP7_75t_L g288 ( .A(n_227), .Y(n_288) );
INVx1_ASAP7_75t_L g235 ( .A(n_228), .Y(n_235) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_228), .Y(n_238) );
INVx3_ASAP7_75t_L g241 ( .A(n_228), .Y(n_241) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_228), .Y(n_257) );
INVx4_ASAP7_75t_SL g244 ( .A(n_229), .Y(n_244) );
BUFx3_ASAP7_75t_L g301 ( .A(n_229), .Y(n_301) );
O2A1O1Ixp33_ASAP7_75t_SL g230 ( .A1(n_231), .A2(n_232), .B(n_236), .C(n_244), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_SL g252 ( .A1(n_232), .A2(n_244), .B(n_253), .C(n_254), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_SL g281 ( .A1(n_232), .A2(n_244), .B(n_282), .C(n_283), .Y(n_281) );
O2A1O1Ixp33_ASAP7_75t_L g319 ( .A1(n_232), .A2(n_244), .B(n_320), .C(n_321), .Y(n_319) );
O2A1O1Ixp33_ASAP7_75t_SL g357 ( .A1(n_232), .A2(n_244), .B(n_358), .C(n_359), .Y(n_357) );
INVx5_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x6_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
BUFx3_ASAP7_75t_L g243 ( .A(n_234), .Y(n_243) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_234), .Y(n_324) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx4_ASAP7_75t_L g284 ( .A(n_238), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
INVx5_ASAP7_75t_L g297 ( .A(n_241), .Y(n_297) );
INVx2_ASAP7_75t_L g275 ( .A(n_242), .Y(n_275) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g258 ( .A(n_243), .Y(n_258) );
INVx1_ASAP7_75t_L g313 ( .A(n_244), .Y(n_313) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_246), .Y(n_250) );
INVx4_ASAP7_75t_L g261 ( .A(n_246), .Y(n_261) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g353 ( .A(n_247), .Y(n_353) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_248), .Y(n_344) );
AND2x2_ASAP7_75t_L g406 ( .A(n_248), .B(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_248), .B(n_263), .Y(n_425) );
INVx1_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g333 ( .A(n_249), .B(n_263), .Y(n_333) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_249), .Y(n_340) );
AND2x2_ASAP7_75t_L g392 ( .A(n_249), .B(n_279), .Y(n_392) );
NAND3xp33_ASAP7_75t_L g417 ( .A(n_249), .B(n_262), .C(n_375), .Y(n_417) );
AND2x2_ASAP7_75t_L g482 ( .A(n_249), .B(n_264), .Y(n_482) );
AND2x2_ASAP7_75t_L g516 ( .A(n_249), .B(n_263), .Y(n_516) );
OA21x2_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_251), .B(n_259), .Y(n_249) );
OA21x2_ASAP7_75t_L g279 ( .A1(n_250), .A2(n_280), .B(n_289), .Y(n_279) );
OA21x2_ASAP7_75t_L g317 ( .A1(n_250), .A2(n_318), .B(n_325), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_256), .B(n_286), .Y(n_285) );
OAI22xp33_ASAP7_75t_L g360 ( .A1(n_256), .A2(n_297), .B1(n_361), .B2(n_362), .Y(n_360) );
INVx4_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g273 ( .A(n_257), .Y(n_273) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_261), .B(n_277), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_261), .B(n_303), .Y(n_302) );
AO21x2_ASAP7_75t_L g306 ( .A1(n_261), .A2(n_307), .B(n_314), .Y(n_306) );
INVxp67_ASAP7_75t_L g342 ( .A(n_262), .Y(n_342) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_278), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_263), .B(n_375), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_263), .B(n_406), .Y(n_414) );
AND2x2_ASAP7_75t_L g464 ( .A(n_263), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g492 ( .A(n_263), .Y(n_492) );
INVx4_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g399 ( .A(n_264), .B(n_392), .Y(n_399) );
BUFx3_ASAP7_75t_L g431 ( .A(n_264), .Y(n_431) );
AO21x2_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_266), .B(n_276), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_268), .B(n_269), .Y(n_266) );
OAI21xp5_ASAP7_75t_L g307 ( .A1(n_268), .A2(n_308), .B(n_309), .Y(n_307) );
O2A1O1Ixp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_272), .B(n_274), .C(n_275), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_L g310 ( .A1(n_272), .A2(n_275), .B(n_311), .C(n_312), .Y(n_310) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g407 ( .A(n_278), .Y(n_407) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_279), .Y(n_376) );
INVx3_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_290), .A2(n_467), .B1(n_469), .B2(n_470), .Y(n_466) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_304), .Y(n_290) );
AND2x2_ASAP7_75t_L g326 ( .A(n_291), .B(n_327), .Y(n_326) );
INVx3_ASAP7_75t_SL g337 ( .A(n_291), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_291), .B(n_370), .Y(n_402) );
OR2x2_ASAP7_75t_L g421 ( .A(n_291), .B(n_305), .Y(n_421) );
AND2x2_ASAP7_75t_L g426 ( .A(n_291), .B(n_378), .Y(n_426) );
AND2x2_ASAP7_75t_L g429 ( .A(n_291), .B(n_371), .Y(n_429) );
AND2x2_ASAP7_75t_L g441 ( .A(n_291), .B(n_317), .Y(n_441) );
AND2x2_ASAP7_75t_L g457 ( .A(n_291), .B(n_306), .Y(n_457) );
AND2x4_ASAP7_75t_L g460 ( .A(n_291), .B(n_328), .Y(n_460) );
OR2x2_ASAP7_75t_L g477 ( .A(n_291), .B(n_413), .Y(n_477) );
OR2x2_ASAP7_75t_L g508 ( .A(n_291), .B(n_350), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_291), .B(n_436), .Y(n_510) );
OR2x6_ASAP7_75t_L g291 ( .A(n_292), .B(n_302), .Y(n_291) );
O2A1O1Ixp33_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_297), .B(n_298), .C(n_299), .Y(n_295) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g359 ( .A(n_300), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g384 ( .A(n_304), .B(n_348), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_304), .B(n_371), .Y(n_503) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_317), .Y(n_304) );
AND2x2_ASAP7_75t_L g336 ( .A(n_305), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g370 ( .A(n_305), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g378 ( .A(n_305), .B(n_350), .Y(n_378) );
AND2x2_ASAP7_75t_L g396 ( .A(n_305), .B(n_328), .Y(n_396) );
OR2x2_ASAP7_75t_L g413 ( .A(n_305), .B(n_371), .Y(n_413) );
INVx2_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
BUFx2_ASAP7_75t_L g329 ( .A(n_306), .Y(n_329) );
AND2x2_ASAP7_75t_L g436 ( .A(n_306), .B(n_317), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx1_ASAP7_75t_L g365 ( .A(n_316), .Y(n_365) );
INVx2_ASAP7_75t_L g328 ( .A(n_317), .Y(n_328) );
INVx1_ASAP7_75t_L g448 ( .A(n_317), .Y(n_448) );
AND2x2_ASAP7_75t_L g498 ( .A(n_317), .B(n_337), .Y(n_498) );
INVx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g347 ( .A(n_327), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g382 ( .A(n_327), .B(n_337), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_327), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
AND2x2_ASAP7_75t_L g369 ( .A(n_328), .B(n_337), .Y(n_369) );
OR2x2_ASAP7_75t_L g485 ( .A(n_329), .B(n_459), .Y(n_485) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_332), .B(n_465), .Y(n_471) );
INVx2_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
OAI32xp33_ASAP7_75t_L g427 ( .A1(n_333), .A2(n_428), .A3(n_430), .B1(n_432), .B2(n_433), .Y(n_427) );
OR2x2_ASAP7_75t_L g444 ( .A(n_333), .B(n_386), .Y(n_444) );
OAI21xp33_ASAP7_75t_SL g469 ( .A1(n_333), .A2(n_343), .B(n_374), .Y(n_469) );
OAI22xp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_338), .B1(n_343), .B2(n_346), .Y(n_334) );
INVxp33_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_336), .B(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_337), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g395 ( .A(n_337), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g495 ( .A(n_337), .B(n_436), .Y(n_495) );
OR2x2_ASAP7_75t_L g519 ( .A(n_337), .B(n_413), .Y(n_519) );
AOI21xp33_ASAP7_75t_L g502 ( .A1(n_338), .A2(n_401), .B(n_503), .Y(n_502) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_342), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g379 ( .A(n_340), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_340), .B(n_345), .Y(n_397) );
AND2x2_ASAP7_75t_L g419 ( .A(n_341), .B(n_392), .Y(n_419) );
INVx1_ASAP7_75t_L g432 ( .A(n_341), .Y(n_432) );
OR2x2_ASAP7_75t_L g437 ( .A(n_341), .B(n_371), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_344), .B(n_386), .Y(n_385) );
OAI22xp33_ASAP7_75t_L g367 ( .A1(n_345), .A2(n_368), .B1(n_373), .B2(n_377), .Y(n_367) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_348), .A2(n_410), .B1(n_417), .B2(n_418), .Y(n_416) );
AND2x2_ASAP7_75t_L g494 ( .A(n_348), .B(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_350), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g513 ( .A(n_350), .B(n_396), .Y(n_513) );
AO21x2_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_354), .B(n_363), .Y(n_350) );
INVx1_ASAP7_75t_L g372 ( .A(n_351), .Y(n_372) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OA21x2_ASAP7_75t_L g371 ( .A1(n_355), .A2(n_364), .B(n_372), .Y(n_371) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_356), .Y(n_523) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_379), .B1(n_380), .B2(n_385), .C(n_387), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_369), .B(n_371), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_369), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g388 ( .A(n_370), .Y(n_388) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_370), .A2(n_476), .B(n_477), .C(n_478), .Y(n_475) );
AND2x2_ASAP7_75t_L g480 ( .A(n_370), .B(n_460), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_SL g518 ( .A1(n_370), .A2(n_459), .B(n_519), .C(n_520), .Y(n_518) );
BUFx3_ASAP7_75t_L g410 ( .A(n_371), .Y(n_410) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_374), .B(n_431), .Y(n_474) );
AOI211xp5_ASAP7_75t_L g493 ( .A1(n_374), .A2(n_494), .B(n_496), .C(n_502), .Y(n_493) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
INVxp67_ASAP7_75t_L g454 ( .A(n_376), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_378), .B(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
AOI211xp5_ASAP7_75t_L g398 ( .A1(n_382), .A2(n_399), .B(n_400), .C(n_408), .Y(n_398) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g483 ( .A(n_386), .Y(n_483) );
OR2x2_ASAP7_75t_L g500 ( .A(n_386), .B(n_430), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B1(n_394), .B2(n_397), .Y(n_387) );
OAI22xp33_ASAP7_75t_L g400 ( .A1(n_389), .A2(n_401), .B1(n_402), .B2(n_403), .Y(n_400) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
OR2x2_ASAP7_75t_L g487 ( .A(n_391), .B(n_431), .Y(n_487) );
INVx1_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g442 ( .A(n_392), .B(n_432), .Y(n_442) );
INVx1_ASAP7_75t_L g450 ( .A(n_393), .Y(n_450) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_396), .B(n_410), .Y(n_458) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_406), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g515 ( .A(n_407), .Y(n_515) );
AOI21xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_411), .B(n_414), .Y(n_408) );
INVx1_ASAP7_75t_L g445 ( .A(n_409), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_410), .B(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_410), .B(n_441), .Y(n_440) );
NAND2x1p5_ASAP7_75t_L g461 ( .A(n_410), .B(n_436), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_410), .B(n_457), .Y(n_468) );
OAI211xp5_ASAP7_75t_L g472 ( .A1(n_410), .A2(n_420), .B(n_460), .C(n_473), .Y(n_472) );
INVx1_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
AOI221xp5_ASAP7_75t_SL g415 ( .A1(n_416), .A2(n_420), .B1(n_422), .B2(n_426), .C(n_427), .Y(n_415) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVxp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_424), .B(n_432), .Y(n_506) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
O2A1O1Ixp33_ASAP7_75t_L g517 ( .A1(n_426), .A2(n_441), .B(n_443), .C(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_429), .B(n_436), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_430), .B(n_483), .Y(n_520) );
CKINVDCx16_ASAP7_75t_R g430 ( .A(n_431), .Y(n_430) );
INVxp33_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .Y(n_434) );
AOI21xp33_ASAP7_75t_SL g446 ( .A1(n_435), .A2(n_447), .B(n_449), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_435), .B(n_508), .Y(n_507) );
INVx2_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_436), .B(n_490), .Y(n_489) );
AOI221xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_442), .B1(n_443), .B2(n_445), .C(n_446), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_442), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g476 ( .A(n_448), .Y(n_476) );
NAND5xp2_ASAP7_75t_L g451 ( .A(n_452), .B(n_479), .C(n_493), .D(n_504), .E(n_517), .Y(n_451) );
AOI211xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_455), .B(n_462), .C(n_475), .Y(n_452) );
INVx2_ASAP7_75t_SL g499 ( .A(n_453), .Y(n_499) );
NAND4xp25_ASAP7_75t_SL g455 ( .A(n_456), .B(n_458), .C(n_459), .D(n_461), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OAI211xp5_ASAP7_75t_SL g462 ( .A1(n_461), .A2(n_463), .B(n_466), .C(n_472), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_464), .Y(n_463) );
AOI221xp5_ASAP7_75t_L g504 ( .A1(n_464), .A2(n_505), .B1(n_507), .B2(n_509), .C(n_511), .Y(n_504) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AOI221xp5_ASAP7_75t_SL g479 ( .A1(n_480), .A2(n_481), .B1(n_484), .B2(n_486), .C(n_488), .Y(n_479) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_487), .A2(n_510), .B1(n_512), .B2(n_514), .Y(n_511) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_499), .B1(n_500), .B2(n_501), .Y(n_496) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_522), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_523), .Y(n_522) );
OAI322xp33_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_526), .A3(n_530), .B1(n_532), .B2(n_534), .C1(n_535), .C2(n_537), .Y(n_524) );
INVx1_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
endmodule