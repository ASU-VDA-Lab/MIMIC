module fake_jpeg_1716_n_131 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_131);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx2_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_53),
.Y(n_58)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_34),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_52),
.B(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_0),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_54),
.Y(n_64)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_54),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_50),
.A2(n_37),
.B1(n_35),
.B2(n_48),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_63),
.B1(n_64),
.B2(n_38),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_40),
.B1(n_45),
.B2(n_42),
.Y(n_63)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_68),
.Y(n_80)
);

AND2x6_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_58),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_37),
.B1(n_35),
.B2(n_48),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_72),
.Y(n_81)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_73),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_61),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_74),
.B(n_76),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_57),
.A2(n_36),
.B1(n_47),
.B2(n_44),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_38),
.B1(n_44),
.B2(n_39),
.Y(n_77)
);

INVxp33_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_61),
.C(n_65),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_86),
.C(n_87),
.Y(n_93)
);

NAND3xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_5),
.C(n_6),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_47),
.Y(n_86)
);

FAx1_ASAP7_75t_SL g87 ( 
.A(n_73),
.B(n_39),
.CI(n_2),
.CON(n_87),
.SN(n_87)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_88),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_36),
.C(n_17),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_15),
.C(n_29),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_1),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_12),
.Y(n_101)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_94),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_66),
.B1(n_3),
.B2(n_4),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_100),
.Y(n_105)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_18),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_9),
.C(n_10),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_16),
.B1(n_32),
.B2(n_30),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_83),
.B(n_22),
.Y(n_110)
);

NAND3xp33_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_101),
.C(n_103),
.Y(n_108)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_83),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_102)
);

NAND2xp33_ASAP7_75t_SL g111 ( 
.A(n_102),
.B(n_104),
.Y(n_111)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_93),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_109),
.Y(n_118)
);

BUFx12f_ASAP7_75t_SL g121 ( 
.A(n_110),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_103),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_87),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_115),
.C(n_96),
.Y(n_117)
);

AO221x1_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.C(n_10),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_11),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_117),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_107),
.A2(n_96),
.B1(n_20),
.B2(n_23),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_119),
.A2(n_121),
.B(n_116),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_124),
.Y(n_126)
);

AOI321xp33_ASAP7_75t_L g124 ( 
.A1(n_118),
.A2(n_109),
.A3(n_120),
.B1(n_121),
.B2(n_105),
.C(n_108),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_105),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_126),
.C(n_106),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_111),
.B(n_26),
.C(n_27),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_19),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_33),
.Y(n_131)
);


endmodule