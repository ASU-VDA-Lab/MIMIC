module fake_netlist_6_1432_n_1666 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1666);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1666;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_124),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_137),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_71),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_66),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_10),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_143),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_78),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_25),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_38),
.Y(n_159)
);

BUFx10_ASAP7_75t_L g160 ( 
.A(n_149),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_45),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_48),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_76),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_47),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_106),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_91),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_27),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_21),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_64),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_77),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_62),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_110),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_68),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_83),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_38),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_107),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_32),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_54),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_10),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_69),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_65),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_141),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_40),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_22),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_36),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_51),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_87),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_23),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_52),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_53),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_130),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_121),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_114),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_24),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_48),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_134),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_82),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_9),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_98),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_22),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_132),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_13),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_104),
.Y(n_207)
);

INVxp33_ASAP7_75t_R g208 ( 
.A(n_92),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_46),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_40),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_30),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_43),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_57),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_14),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_109),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_112),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_0),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_81),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_13),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_105),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_15),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_27),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_14),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_51),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_5),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_75),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_23),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_29),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_113),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_120),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_111),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_63),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_8),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_39),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_73),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_58),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_136),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_31),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_24),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_103),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_12),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_2),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_15),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_8),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_16),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_147),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_99),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_85),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_125),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_56),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_148),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g252 ( 
.A(n_47),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_95),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_45),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_3),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_18),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_1),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_18),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_5),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_145),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_32),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_30),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_6),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_108),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_89),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_11),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_1),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_57),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_56),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_4),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_0),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_84),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_61),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_59),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_7),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_29),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_55),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_88),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_33),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_55),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_52),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_34),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_100),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_43),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_96),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_127),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_17),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_115),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_7),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_9),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_11),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_35),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_102),
.Y(n_293)
);

BUFx10_ASAP7_75t_L g294 ( 
.A(n_35),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_60),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_128),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_33),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_166),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_191),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_166),
.Y(n_300)
);

INVxp33_ASAP7_75t_L g301 ( 
.A(n_182),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_166),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_196),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_203),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_178),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_166),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_205),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_166),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_166),
.B(n_168),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_166),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_198),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_166),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_215),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_222),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_239),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_210),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_265),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_210),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_289),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_210),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_150),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_193),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_210),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_202),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_210),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_150),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_204),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_213),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_152),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_227),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_227),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_296),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_168),
.B(n_220),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_152),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_227),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_156),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_155),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_156),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_L g339 ( 
.A(n_242),
.B(n_2),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_221),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_160),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_223),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_164),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_227),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_164),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_165),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_165),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_220),
.B(n_3),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_175),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_227),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_153),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_175),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_176),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_155),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_290),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_290),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_176),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_290),
.Y(n_358)
);

BUFx10_ASAP7_75t_L g359 ( 
.A(n_173),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_219),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_290),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_173),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_184),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_184),
.Y(n_364)
);

NOR2xp67_ASAP7_75t_L g365 ( 
.A(n_242),
.B(n_4),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_153),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_290),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_159),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_185),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_185),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_235),
.Y(n_371)
);

INVxp33_ASAP7_75t_L g372 ( 
.A(n_171),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_159),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_316),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_316),
.B(n_151),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_318),
.B(n_151),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_366),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_303),
.B(n_172),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_359),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_318),
.Y(n_380)
);

OA21x2_ASAP7_75t_L g381 ( 
.A1(n_362),
.A2(n_186),
.B(n_172),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_320),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_311),
.Y(n_383)
);

AND2x6_ASAP7_75t_L g384 ( 
.A(n_333),
.B(n_173),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_360),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_366),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_359),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_343),
.B(n_179),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_307),
.B(n_313),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_351),
.B(n_217),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_320),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_323),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_366),
.B(n_345),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_323),
.Y(n_394)
);

INVx5_ASAP7_75t_L g395 ( 
.A(n_359),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_325),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_325),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_317),
.A2(n_275),
.B1(n_291),
.B2(n_282),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_330),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_330),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_331),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_331),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_346),
.B(n_186),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_335),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_335),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_332),
.B(n_217),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_359),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_372),
.B(n_244),
.Y(n_408)
);

AND3x1_ASAP7_75t_L g409 ( 
.A(n_348),
.B(n_190),
.C(n_181),
.Y(n_409)
);

AND2x6_ASAP7_75t_L g410 ( 
.A(n_362),
.B(n_173),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_344),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_344),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_347),
.B(n_349),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_350),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_350),
.B(n_207),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_360),
.A2(n_158),
.B1(n_161),
.B2(n_292),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_355),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_355),
.B(n_207),
.Y(n_418)
);

OR2x6_ASAP7_75t_L g419 ( 
.A(n_339),
.B(n_181),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_356),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_341),
.A2(n_258),
.B1(n_214),
.B2(n_282),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_362),
.Y(n_422)
);

INVx5_ASAP7_75t_L g423 ( 
.A(n_341),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_356),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_358),
.Y(n_425)
);

AND2x6_ASAP7_75t_L g426 ( 
.A(n_298),
.B(n_173),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_358),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_321),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_361),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_315),
.B(n_160),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_319),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_357),
.B(n_226),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_361),
.B(n_226),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_322),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_367),
.B(n_230),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_367),
.B(n_230),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_309),
.B(n_154),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_298),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_305),
.A2(n_270),
.B1(n_280),
.B2(n_162),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_300),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_326),
.B(n_329),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_300),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_425),
.Y(n_443)
);

NAND3xp33_ASAP7_75t_L g444 ( 
.A(n_388),
.B(n_327),
.C(n_324),
.Y(n_444)
);

BUFx4f_ASAP7_75t_L g445 ( 
.A(n_437),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_393),
.B(n_363),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_438),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_377),
.B(n_364),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_438),
.Y(n_449)
);

NAND3xp33_ASAP7_75t_L g450 ( 
.A(n_390),
.B(n_340),
.C(n_328),
.Y(n_450)
);

INVx5_ASAP7_75t_L g451 ( 
.A(n_426),
.Y(n_451)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_379),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_377),
.B(n_371),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_425),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_413),
.A2(n_299),
.B1(n_304),
.B2(n_369),
.Y(n_455)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_379),
.Y(n_456)
);

AND3x2_ASAP7_75t_L g457 ( 
.A(n_431),
.B(n_169),
.C(n_157),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g458 ( 
.A(n_385),
.Y(n_458)
);

OR2x2_ASAP7_75t_L g459 ( 
.A(n_408),
.B(n_337),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_442),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_442),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_380),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_378),
.B(n_342),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_437),
.B(n_302),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_440),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_380),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_440),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_L g468 ( 
.A1(n_437),
.A2(n_365),
.B1(n_339),
.B2(n_212),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_400),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_SL g470 ( 
.A(n_403),
.B(n_162),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_379),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_442),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_389),
.B(n_334),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_386),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_374),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_425),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_386),
.B(n_368),
.Y(n_477)
);

OR2x6_ASAP7_75t_L g478 ( 
.A(n_419),
.B(n_244),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_419),
.B(n_368),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_432),
.B(n_302),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_400),
.Y(n_481)
);

NAND3xp33_ASAP7_75t_L g482 ( 
.A(n_390),
.B(n_354),
.C(n_314),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_408),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_423),
.B(n_434),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_384),
.A2(n_212),
.B1(n_256),
.B2(n_259),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_379),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_425),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_405),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_379),
.B(n_306),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_430),
.A2(n_336),
.B1(n_370),
.B2(n_353),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_374),
.Y(n_491)
);

NAND2xp33_ASAP7_75t_L g492 ( 
.A(n_384),
.B(n_180),
.Y(n_492)
);

INVx6_ASAP7_75t_L g493 ( 
.A(n_387),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_441),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_405),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_382),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_419),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_423),
.B(n_338),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_382),
.Y(n_499)
);

NAND3xp33_ASAP7_75t_L g500 ( 
.A(n_406),
.B(n_301),
.C(n_187),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_387),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_423),
.B(n_352),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_412),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_391),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_419),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_423),
.B(n_160),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_419),
.Y(n_507)
);

BUFx10_ASAP7_75t_L g508 ( 
.A(n_384),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_406),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_391),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_383),
.B(n_208),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_387),
.B(n_407),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_428),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_423),
.B(n_235),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_423),
.B(n_237),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_412),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_392),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_392),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_394),
.Y(n_519)
);

OR2x6_ASAP7_75t_L g520 ( 
.A(n_434),
.B(n_259),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_398),
.B(n_225),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_387),
.B(n_306),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_387),
.B(n_308),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_407),
.Y(n_524)
);

OR2x6_ASAP7_75t_L g525 ( 
.A(n_431),
.B(n_261),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_425),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_420),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_422),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_396),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_409),
.A2(n_249),
.B1(n_197),
.B2(n_238),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_422),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_439),
.B(n_237),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_407),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_375),
.B(n_373),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_422),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_375),
.B(n_373),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_396),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_441),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_397),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_397),
.Y(n_540)
);

NAND2xp33_ASAP7_75t_R g541 ( 
.A(n_381),
.B(n_240),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_375),
.B(n_312),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_399),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_420),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_407),
.B(n_308),
.Y(n_545)
);

AND2x6_ASAP7_75t_L g546 ( 
.A(n_407),
.B(n_180),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_416),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_399),
.Y(n_548)
);

INVxp33_ASAP7_75t_L g549 ( 
.A(n_416),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_401),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_439),
.B(n_240),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_381),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_384),
.B(n_401),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_381),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_402),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_402),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_404),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_404),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_375),
.B(n_312),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_411),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_411),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_376),
.Y(n_562)
);

AND2x6_ASAP7_75t_L g563 ( 
.A(n_376),
.B(n_180),
.Y(n_563)
);

NOR2x1p5_ASAP7_75t_L g564 ( 
.A(n_414),
.B(n_170),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_414),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_417),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_417),
.Y(n_567)
);

BUFx6f_ASAP7_75t_SL g568 ( 
.A(n_384),
.Y(n_568)
);

INVx5_ASAP7_75t_L g569 ( 
.A(n_426),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_381),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_384),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_436),
.B(n_310),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_384),
.B(n_310),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_376),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_376),
.B(n_415),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_424),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_415),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_415),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_415),
.A2(n_297),
.B1(n_187),
.B2(n_291),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_428),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_427),
.Y(n_581)
);

BUFx4f_ASAP7_75t_L g582 ( 
.A(n_426),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_427),
.Y(n_583)
);

AND2x6_ASAP7_75t_L g584 ( 
.A(n_418),
.B(n_180),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_418),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_418),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_429),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_418),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_429),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_458),
.B(n_421),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_548),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_548),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_555),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_480),
.B(n_433),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_446),
.B(n_433),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_575),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_445),
.B(n_395),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_513),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_445),
.B(n_509),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_463),
.B(n_444),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_445),
.B(n_395),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_555),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_575),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_509),
.A2(n_231),
.B1(n_278),
.B2(n_251),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_483),
.B(n_395),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_556),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_556),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_447),
.B(n_483),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_447),
.B(n_433),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_449),
.B(n_433),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_585),
.B(n_586),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_450),
.B(n_421),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_585),
.B(n_435),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_562),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_562),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_574),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_557),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_513),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_557),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_586),
.B(n_435),
.Y(n_620)
);

NOR3xp33_ASAP7_75t_L g621 ( 
.A(n_511),
.B(n_269),
.C(n_188),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_542),
.B(n_435),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_459),
.B(n_170),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_574),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_474),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_542),
.B(n_435),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_464),
.B(n_395),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_559),
.B(n_572),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_559),
.B(n_436),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_459),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_572),
.B(n_436),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_477),
.B(n_222),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_578),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_577),
.B(n_436),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_578),
.B(n_395),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_577),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_448),
.B(n_246),
.Y(n_637)
);

INVxp33_ASAP7_75t_L g638 ( 
.A(n_500),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_578),
.B(n_588),
.Y(n_639)
);

NAND2xp33_ASAP7_75t_SL g640 ( 
.A(n_468),
.B(n_180),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_560),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_560),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_564),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_578),
.B(n_395),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_479),
.B(n_426),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_479),
.B(n_426),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_565),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_588),
.B(n_260),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_479),
.B(n_426),
.Y(n_649)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_521),
.B(n_189),
.Y(n_650)
);

NAND2xp33_ASAP7_75t_L g651 ( 
.A(n_485),
.B(n_260),
.Y(n_651)
);

OR2x2_ASAP7_75t_SL g652 ( 
.A(n_521),
.B(n_261),
.Y(n_652)
);

INVx8_ASAP7_75t_L g653 ( 
.A(n_478),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_452),
.B(n_163),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_565),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_452),
.A2(n_247),
.B(n_295),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_477),
.Y(n_657)
);

NOR2xp67_ASAP7_75t_L g658 ( 
.A(n_455),
.B(n_490),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_534),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_534),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_453),
.B(n_246),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_456),
.B(n_167),
.Y(n_662)
);

O2A1O1Ixp33_ASAP7_75t_L g663 ( 
.A1(n_497),
.A2(n_206),
.B(n_211),
.C(n_209),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_588),
.B(n_497),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_534),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_474),
.B(n_174),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_566),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_456),
.B(n_471),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_588),
.B(n_260),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_473),
.B(n_251),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_588),
.Y(n_671)
);

NAND2xp33_ASAP7_75t_L g672 ( 
.A(n_571),
.B(n_260),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_456),
.B(n_177),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_566),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_536),
.Y(n_675)
);

A2O1A1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_549),
.A2(n_224),
.B(n_228),
.C(n_199),
.Y(n_676)
);

OAI22xp5_ASAP7_75t_SL g677 ( 
.A1(n_580),
.A2(n_243),
.B1(n_297),
.B2(n_254),
.Y(n_677)
);

INVxp67_ASAP7_75t_L g678 ( 
.A(n_482),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_505),
.A2(n_253),
.B1(n_264),
.B2(n_293),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_505),
.B(n_260),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_525),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_507),
.B(n_508),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_507),
.B(n_195),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_475),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_475),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_471),
.B(n_200),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_510),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_471),
.B(n_201),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_501),
.B(n_216),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_536),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_536),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_L g692 ( 
.A(n_571),
.B(n_410),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_508),
.B(n_582),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_501),
.B(n_218),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_510),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_520),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_532),
.B(n_253),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_517),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_508),
.B(n_229),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_517),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_533),
.B(n_491),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_533),
.B(n_496),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_499),
.B(n_232),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_518),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_528),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_525),
.B(n_222),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_518),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_504),
.B(n_567),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_582),
.B(n_236),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_519),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_519),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_582),
.B(n_248),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_520),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_478),
.B(n_520),
.Y(n_714)
);

NOR3xp33_ASAP7_75t_L g715 ( 
.A(n_551),
.B(n_470),
.C(n_494),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_529),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_529),
.B(n_272),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_537),
.Y(n_718)
);

NAND3xp33_ASAP7_75t_L g719 ( 
.A(n_470),
.B(n_293),
.C(n_288),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_478),
.A2(n_273),
.B1(n_274),
.B2(n_264),
.Y(n_720)
);

INVx4_ASAP7_75t_L g721 ( 
.A(n_493),
.Y(n_721)
);

INVxp33_ASAP7_75t_L g722 ( 
.A(n_547),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_573),
.B(n_286),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_539),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_540),
.Y(n_725)
);

OR2x6_ASAP7_75t_L g726 ( 
.A(n_478),
.B(n_183),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_520),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_540),
.B(n_273),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_543),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_543),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_550),
.B(n_274),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_550),
.Y(n_732)
);

OAI221xp5_ASAP7_75t_L g733 ( 
.A1(n_530),
.A2(n_284),
.B1(n_241),
.B2(n_234),
.C(n_194),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_L g734 ( 
.A(n_546),
.B(n_410),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_558),
.Y(n_735)
);

NOR3xp33_ASAP7_75t_L g736 ( 
.A(n_538),
.B(n_287),
.C(n_192),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_558),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_541),
.A2(n_283),
.B1(n_288),
.B2(n_285),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_561),
.B(n_576),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_561),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_576),
.Y(n_741)
);

OAI22xp33_ASAP7_75t_L g742 ( 
.A1(n_525),
.A2(n_589),
.B1(n_587),
.B2(n_583),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_581),
.B(n_583),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_581),
.A2(n_268),
.B1(n_245),
.B2(n_250),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_589),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_460),
.B(n_283),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_525),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_528),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_579),
.Y(n_749)
);

INVxp67_ASAP7_75t_L g750 ( 
.A(n_498),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_461),
.B(n_285),
.Y(n_751)
);

AO21x1_ASAP7_75t_L g752 ( 
.A1(n_742),
.A2(n_553),
.B(n_472),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_636),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_600),
.A2(n_484),
.B1(n_502),
.B2(n_506),
.Y(n_754)
);

INVx1_ASAP7_75t_SL g755 ( 
.A(n_630),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_670),
.A2(n_515),
.B1(n_514),
.B2(n_472),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_668),
.A2(n_524),
.B(n_486),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_595),
.B(n_552),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_608),
.B(n_552),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_640),
.A2(n_492),
.B1(n_568),
.B2(n_271),
.Y(n_760)
);

NAND3xp33_ASAP7_75t_L g761 ( 
.A(n_697),
.B(n_457),
.C(n_263),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_684),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_596),
.A2(n_545),
.B1(n_489),
.B2(n_522),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_695),
.B(n_552),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_603),
.A2(n_523),
.B1(n_568),
.B2(n_467),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_639),
.A2(n_486),
.B(n_524),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_722),
.B(n_554),
.Y(n_767)
);

OAI21xp5_ASAP7_75t_L g768 ( 
.A1(n_628),
.A2(n_626),
.B(n_622),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_722),
.B(n_554),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_666),
.Y(n_770)
);

AO21x2_ASAP7_75t_L g771 ( 
.A1(n_599),
.A2(n_512),
.B(n_492),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_639),
.A2(n_570),
.B(n_554),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_684),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_685),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_685),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_700),
.B(n_570),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_687),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_707),
.B(n_570),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_594),
.A2(n_451),
.B(n_569),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_710),
.B(n_465),
.Y(n_780)
);

BUFx2_ASAP7_75t_L g781 ( 
.A(n_714),
.Y(n_781)
);

O2A1O1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_676),
.A2(n_467),
.B(n_465),
.C(n_462),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_711),
.B(n_528),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_724),
.B(n_531),
.Y(n_784)
);

INVx4_ASAP7_75t_L g785 ( 
.A(n_633),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_625),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_725),
.B(n_531),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_623),
.B(n_580),
.Y(n_788)
);

AOI21x1_ASAP7_75t_L g789 ( 
.A1(n_605),
.A2(n_488),
.B(n_481),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_729),
.B(n_531),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_730),
.B(n_535),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_638),
.B(n_535),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_SL g793 ( 
.A(n_590),
.B(n_252),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_737),
.B(n_740),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_698),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_741),
.B(n_443),
.Y(n_796)
);

AOI21x1_ASAP7_75t_L g797 ( 
.A1(n_605),
.A2(n_481),
.B(n_466),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_611),
.A2(n_451),
.B(n_569),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_633),
.B(n_451),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_637),
.B(n_443),
.Y(n_800)
);

OAI22xp5_ASAP7_75t_L g801 ( 
.A1(n_750),
.A2(n_493),
.B1(n_462),
.B2(n_495),
.Y(n_801)
);

OAI21xp5_ASAP7_75t_L g802 ( 
.A1(n_629),
.A2(n_503),
.B(n_469),
.Y(n_802)
);

O2A1O1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_676),
.A2(n_749),
.B(n_733),
.C(n_743),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_661),
.B(n_443),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_704),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_706),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_633),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_704),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_739),
.B(n_454),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_690),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_633),
.B(n_451),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_666),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_634),
.A2(n_569),
.B(n_454),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_716),
.Y(n_814)
);

OAI21xp33_ASAP7_75t_L g815 ( 
.A1(n_612),
.A2(n_255),
.B(n_254),
.Y(n_815)
);

O2A1O1Ixp5_ASAP7_75t_L g816 ( 
.A1(n_709),
.A2(n_487),
.B(n_476),
.C(n_454),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_632),
.B(n_252),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_638),
.B(n_476),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_678),
.B(n_476),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_640),
.A2(n_279),
.B1(n_257),
.B2(n_277),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_613),
.A2(n_620),
.B(n_631),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_693),
.A2(n_569),
.B(n_487),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_721),
.A2(n_526),
.B(n_493),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_650),
.B(n_526),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_721),
.A2(n_516),
.B(n_469),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_716),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_625),
.B(n_252),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_718),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_671),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_732),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_732),
.B(n_503),
.Y(n_831)
);

A2O1A1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_658),
.A2(n_276),
.B(n_233),
.C(n_238),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_671),
.B(n_690),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_651),
.A2(n_584),
.B1(n_563),
.B2(n_544),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_599),
.A2(n_584),
.B1(n_563),
.B2(n_546),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_735),
.B(n_516),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_735),
.B(n_527),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_721),
.A2(n_544),
.B(n_527),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_671),
.B(n_267),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_652),
.B(n_189),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_745),
.B(n_546),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_745),
.B(n_708),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_657),
.B(n_546),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_738),
.B(n_233),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_701),
.A2(n_702),
.B(n_627),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_675),
.A2(n_584),
.B1(n_563),
.B2(n_546),
.Y(n_846)
);

NAND3xp33_ASAP7_75t_L g847 ( 
.A(n_621),
.B(n_267),
.C(n_255),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_690),
.A2(n_584),
.B1(n_563),
.B2(n_546),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_691),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_666),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_691),
.B(n_671),
.Y(n_851)
);

OAI21xp33_ASAP7_75t_L g852 ( 
.A1(n_604),
.A2(n_243),
.B(n_262),
.Y(n_852)
);

AOI21xp33_ASAP7_75t_L g853 ( 
.A1(n_659),
.A2(n_262),
.B(n_263),
.Y(n_853)
);

O2A1O1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_683),
.A2(n_563),
.B(n_584),
.C(n_281),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_627),
.A2(n_584),
.B(n_563),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_681),
.B(n_294),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_691),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_645),
.A2(n_649),
.B(n_646),
.Y(n_858)
);

A2O1A1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_663),
.A2(n_266),
.B(n_270),
.C(n_280),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_705),
.B(n_266),
.Y(n_860)
);

O2A1O1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_683),
.A2(n_281),
.B(n_294),
.C(n_16),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_L g862 ( 
.A1(n_714),
.A2(n_72),
.B1(n_74),
.B2(n_144),
.Y(n_862)
);

INVxp67_ASAP7_75t_L g863 ( 
.A(n_643),
.Y(n_863)
);

NOR2xp67_ASAP7_75t_L g864 ( 
.A(n_719),
.B(n_67),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_651),
.A2(n_294),
.B(n_12),
.C(n_17),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_598),
.B(n_6),
.Y(n_866)
);

NAND2xp33_ASAP7_75t_L g867 ( 
.A(n_653),
.B(n_410),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_614),
.B(n_410),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_727),
.A2(n_19),
.B(n_20),
.C(n_21),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_714),
.A2(n_79),
.B1(n_142),
.B2(n_140),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_615),
.B(n_410),
.Y(n_871)
);

NAND2xp33_ASAP7_75t_L g872 ( 
.A(n_653),
.B(n_410),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_705),
.B(n_138),
.Y(n_873)
);

BUFx8_ASAP7_75t_SL g874 ( 
.A(n_618),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_616),
.B(n_19),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_624),
.B(n_660),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_696),
.B(n_20),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_591),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_665),
.B(n_25),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_664),
.A2(n_70),
.B(n_131),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_591),
.B(n_26),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_592),
.Y(n_882)
);

OR2x2_ASAP7_75t_L g883 ( 
.A(n_728),
.B(n_26),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_705),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_664),
.A2(n_86),
.B(n_129),
.Y(n_885)
);

OAI21xp33_ASAP7_75t_L g886 ( 
.A1(n_744),
.A2(n_28),
.B(n_31),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_592),
.B(n_28),
.Y(n_887)
);

AOI21x1_ASAP7_75t_L g888 ( 
.A1(n_635),
.A2(n_90),
.B(n_123),
.Y(n_888)
);

AOI21x1_ASAP7_75t_L g889 ( 
.A1(n_635),
.A2(n_133),
.B(n_122),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_731),
.B(n_713),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_597),
.A2(n_119),
.B(n_118),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_597),
.A2(n_117),
.B(n_116),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_727),
.Y(n_893)
);

INVx1_ASAP7_75t_SL g894 ( 
.A(n_677),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_680),
.A2(n_34),
.B(n_36),
.C(n_37),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_593),
.B(n_37),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_748),
.B(n_101),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_593),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_602),
.B(n_39),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_748),
.B(n_97),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_602),
.B(n_41),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_606),
.B(n_41),
.Y(n_902)
);

AOI21x1_ASAP7_75t_L g903 ( 
.A1(n_644),
.A2(n_94),
.B(n_93),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_606),
.Y(n_904)
);

INVx11_ASAP7_75t_L g905 ( 
.A(n_715),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_601),
.A2(n_42),
.B(n_44),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_601),
.A2(n_42),
.B(n_44),
.Y(n_907)
);

BUFx4f_ASAP7_75t_L g908 ( 
.A(n_653),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_607),
.B(n_46),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_747),
.B(n_49),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_746),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_609),
.A2(n_49),
.B(n_50),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_607),
.B(n_50),
.Y(n_913)
);

NOR3xp33_ASAP7_75t_L g914 ( 
.A(n_747),
.B(n_53),
.C(n_54),
.Y(n_914)
);

NAND2xp33_ASAP7_75t_L g915 ( 
.A(n_653),
.B(n_682),
.Y(n_915)
);

AOI21x1_ASAP7_75t_L g916 ( 
.A1(n_644),
.A2(n_688),
.B(n_673),
.Y(n_916)
);

INVx1_ASAP7_75t_SL g917 ( 
.A(n_751),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_682),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_617),
.B(n_655),
.Y(n_919)
);

BUFx8_ASAP7_75t_L g920 ( 
.A(n_617),
.Y(n_920)
);

A2O1A1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_720),
.A2(n_655),
.B(n_619),
.C(n_641),
.Y(n_921)
);

INVxp67_ASAP7_75t_L g922 ( 
.A(n_736),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_610),
.A2(n_699),
.B(n_672),
.Y(n_923)
);

BUFx12f_ASAP7_75t_L g924 ( 
.A(n_726),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_641),
.B(n_642),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_699),
.A2(n_672),
.B(n_689),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_654),
.A2(n_694),
.B(n_686),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_662),
.A2(n_709),
.B(n_712),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_712),
.A2(n_692),
.B(n_680),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_692),
.A2(n_723),
.B(n_648),
.Y(n_930)
);

AOI21xp33_ASAP7_75t_L g931 ( 
.A1(n_844),
.A2(n_679),
.B(n_726),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_762),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_773),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_821),
.A2(n_734),
.B(n_648),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_792),
.B(n_647),
.Y(n_935)
);

NAND2x1p5_ASAP7_75t_L g936 ( 
.A(n_908),
.B(n_667),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_774),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_917),
.B(n_726),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_754),
.B(n_703),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_775),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_927),
.A2(n_734),
.B(n_669),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_842),
.A2(n_726),
.B1(n_667),
.B2(n_674),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_777),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_911),
.B(n_717),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_807),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_874),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_770),
.B(n_656),
.Y(n_947)
);

NAND3xp33_ASAP7_75t_SL g948 ( 
.A(n_793),
.B(n_844),
.C(n_815),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_768),
.A2(n_758),
.B(n_772),
.Y(n_949)
);

OAI21xp33_ASAP7_75t_L g950 ( 
.A1(n_886),
.A2(n_912),
.B(n_852),
.Y(n_950)
);

O2A1O1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_832),
.A2(n_803),
.B(n_859),
.C(n_861),
.Y(n_951)
);

CKINVDCx8_ASAP7_75t_R g952 ( 
.A(n_781),
.Y(n_952)
);

NAND2x1_ASAP7_75t_L g953 ( 
.A(n_785),
.B(n_807),
.Y(n_953)
);

OR2x6_ASAP7_75t_L g954 ( 
.A(n_924),
.B(n_786),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_R g955 ( 
.A(n_915),
.B(n_908),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_812),
.B(n_890),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_SL g957 ( 
.A(n_862),
.B(n_870),
.Y(n_957)
);

NOR3xp33_ASAP7_75t_SL g958 ( 
.A(n_847),
.B(n_832),
.C(n_761),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_807),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_SL g960 ( 
.A(n_785),
.B(n_865),
.Y(n_960)
);

AND2x6_ASAP7_75t_L g961 ( 
.A(n_918),
.B(n_884),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_795),
.Y(n_962)
);

INVxp67_ASAP7_75t_L g963 ( 
.A(n_755),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_805),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_756),
.A2(n_849),
.B1(n_810),
.B2(n_851),
.Y(n_965)
);

O2A1O1Ixp5_ASAP7_75t_L g966 ( 
.A1(n_752),
.A2(n_928),
.B(n_926),
.C(n_923),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_893),
.B(n_850),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_767),
.A2(n_769),
.B1(n_913),
.B2(n_824),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_828),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_859),
.A2(n_839),
.B(n_860),
.C(n_875),
.Y(n_970)
);

AOI21xp33_ASAP7_75t_L g971 ( 
.A1(n_890),
.A2(n_806),
.B(n_788),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_830),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_819),
.B(n_818),
.Y(n_973)
);

OAI22x1_ASAP7_75t_L g974 ( 
.A1(n_894),
.A2(n_922),
.B1(n_840),
.B2(n_866),
.Y(n_974)
);

BUFx2_ASAP7_75t_L g975 ( 
.A(n_920),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_810),
.A2(n_849),
.B1(n_765),
.B2(n_794),
.Y(n_976)
);

BUFx4f_ASAP7_75t_L g977 ( 
.A(n_918),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_882),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_807),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_920),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_898),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_819),
.B(n_818),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_839),
.A2(n_860),
.B(n_853),
.C(n_883),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_808),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_913),
.A2(n_865),
.B(n_869),
.C(n_879),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_759),
.B(n_814),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_817),
.B(n_827),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_826),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_905),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_845),
.A2(n_929),
.B(n_778),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_878),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_876),
.B(n_753),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_SL g993 ( 
.A1(n_840),
.A2(n_804),
.B(n_800),
.C(n_802),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_764),
.A2(n_776),
.B(n_858),
.Y(n_994)
);

NAND2x1p5_ASAP7_75t_L g995 ( 
.A(n_829),
.B(n_857),
.Y(n_995)
);

CKINVDCx8_ASAP7_75t_R g996 ( 
.A(n_918),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_863),
.B(n_877),
.Y(n_997)
);

O2A1O1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_869),
.A2(n_921),
.B(n_895),
.C(n_914),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_904),
.Y(n_999)
);

OAI21xp33_ASAP7_75t_L g1000 ( 
.A1(n_820),
.A2(n_910),
.B(n_760),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_856),
.B(n_833),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_780),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_930),
.A2(n_809),
.B(n_757),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_820),
.B(n_919),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_833),
.B(n_783),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_823),
.A2(n_766),
.B(n_779),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_763),
.B(n_784),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_787),
.B(n_791),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_760),
.A2(n_921),
.B1(n_829),
.B2(n_790),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_897),
.A2(n_900),
.B1(n_864),
.B2(n_909),
.Y(n_1010)
);

CKINVDCx14_ASAP7_75t_R g1011 ( 
.A(n_829),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_897),
.A2(n_900),
.B1(n_899),
.B2(n_881),
.Y(n_1012)
);

AOI21x1_ASAP7_75t_L g1013 ( 
.A1(n_916),
.A2(n_789),
.B(n_797),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_831),
.A2(n_836),
.B(n_837),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_829),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_843),
.A2(n_811),
.B(n_799),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_796),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_834),
.A2(n_841),
.B1(n_848),
.B2(n_873),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_887),
.A2(n_902),
.B1(n_896),
.B2(n_901),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_782),
.A2(n_854),
.B(n_907),
.C(n_906),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_801),
.Y(n_1021)
);

BUFx8_ASAP7_75t_L g1022 ( 
.A(n_880),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_925),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_868),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_888),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_867),
.A2(n_872),
.B(n_816),
.C(n_871),
.Y(n_1026)
);

NOR3xp33_ASAP7_75t_L g1027 ( 
.A(n_885),
.B(n_891),
.C(n_892),
.Y(n_1027)
);

INVx5_ASAP7_75t_L g1028 ( 
.A(n_889),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_771),
.B(n_846),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_834),
.B(n_825),
.Y(n_1030)
);

NAND2xp33_ASAP7_75t_SL g1031 ( 
.A(n_903),
.B(n_835),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_855),
.A2(n_813),
.B(n_838),
.C(n_822),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_798),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_773),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_762),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_874),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_917),
.B(n_458),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_762),
.Y(n_1038)
);

BUFx12f_ASAP7_75t_L g1039 ( 
.A(n_924),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_807),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_817),
.B(n_385),
.Y(n_1041)
);

NAND2x1p5_ASAP7_75t_L g1042 ( 
.A(n_908),
.B(n_785),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_803),
.A2(n_600),
.B(n_670),
.C(n_612),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_SL g1044 ( 
.A(n_908),
.B(n_612),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_754),
.A2(n_445),
.B1(n_842),
.B2(n_595),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_781),
.B(n_786),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_754),
.A2(n_445),
.B1(n_842),
.B2(n_595),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_792),
.B(n_600),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_917),
.B(n_458),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_767),
.A2(n_612),
.B1(n_769),
.B2(n_600),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_917),
.B(n_458),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_917),
.B(n_458),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_917),
.B(n_458),
.Y(n_1053)
);

CKINVDCx6p67_ASAP7_75t_R g1054 ( 
.A(n_924),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_917),
.B(n_458),
.Y(n_1055)
);

AOI221xp5_ASAP7_75t_L g1056 ( 
.A1(n_815),
.A2(n_549),
.B1(n_547),
.B2(n_612),
.C(n_844),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_807),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_755),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_754),
.A2(n_445),
.B1(n_842),
.B2(n_595),
.Y(n_1059)
);

BUFx5_ASAP7_75t_L g1060 ( 
.A(n_773),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_917),
.B(n_458),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_762),
.Y(n_1062)
);

NAND2xp33_ASAP7_75t_SL g1063 ( 
.A(n_883),
.B(n_638),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_754),
.A2(n_445),
.B1(n_842),
.B2(n_595),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_991),
.Y(n_1065)
);

INVxp67_ASAP7_75t_L g1066 ( 
.A(n_1052),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_1053),
.B(n_1061),
.Y(n_1067)
);

AOI221x1_ASAP7_75t_L g1068 ( 
.A1(n_1043),
.A2(n_948),
.B1(n_950),
.B2(n_1031),
.C(n_1027),
.Y(n_1068)
);

BUFx10_ASAP7_75t_L g1069 ( 
.A(n_946),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_1048),
.A2(n_1050),
.B(n_1047),
.Y(n_1070)
);

NAND3xp33_ASAP7_75t_L g1071 ( 
.A(n_1056),
.B(n_931),
.C(n_958),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_933),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_1044),
.A2(n_1041),
.B1(n_957),
.B2(n_987),
.Y(n_1073)
);

AO31x2_ASAP7_75t_L g1074 ( 
.A1(n_1045),
.A2(n_1064),
.A3(n_1059),
.B(n_1020),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_971),
.A2(n_983),
.B(n_950),
.C(n_957),
.Y(n_1075)
);

AO31x2_ASAP7_75t_L g1076 ( 
.A1(n_1029),
.A2(n_1009),
.A3(n_1032),
.B(n_1003),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1002),
.B(n_1050),
.Y(n_1077)
);

NOR2x1_ASAP7_75t_R g1078 ( 
.A(n_1036),
.B(n_980),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_939),
.A2(n_994),
.B(n_941),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_1007),
.A2(n_934),
.B(n_1014),
.Y(n_1080)
);

AOI221x1_ASAP7_75t_L g1081 ( 
.A1(n_974),
.A2(n_973),
.B1(n_982),
.B2(n_1063),
.C(n_976),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_1037),
.B(n_1049),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_996),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_989),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_966),
.A2(n_1008),
.B(n_993),
.Y(n_1085)
);

OAI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_968),
.A2(n_970),
.B(n_985),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_945),
.Y(n_1087)
);

BUFx10_ASAP7_75t_L g1088 ( 
.A(n_938),
.Y(n_1088)
);

AO32x2_ASAP7_75t_L g1089 ( 
.A1(n_965),
.A2(n_942),
.A3(n_1018),
.B1(n_951),
.B2(n_998),
.Y(n_1089)
);

OR2x2_ASAP7_75t_L g1090 ( 
.A(n_1051),
.B(n_1055),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1001),
.B(n_992),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_1013),
.A2(n_1016),
.B(n_1026),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_1044),
.B(n_963),
.Y(n_1093)
);

NOR2xp67_ASAP7_75t_L g1094 ( 
.A(n_1058),
.B(n_997),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1030),
.A2(n_1012),
.B(n_1019),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_945),
.Y(n_1096)
);

NAND3xp33_ASAP7_75t_L g1097 ( 
.A(n_956),
.B(n_944),
.C(n_1010),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1012),
.A2(n_986),
.B(n_1010),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_937),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1017),
.B(n_935),
.Y(n_1100)
);

INVx4_ASAP7_75t_L g1101 ( 
.A(n_945),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_1039),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_952),
.B(n_967),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_960),
.A2(n_1021),
.B(n_1000),
.C(n_947),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_968),
.A2(n_977),
.B1(n_1004),
.B2(n_1000),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_940),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1005),
.B(n_967),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_1046),
.B(n_975),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_1046),
.B(n_954),
.Y(n_1109)
);

AOI221x1_ASAP7_75t_L g1110 ( 
.A1(n_1025),
.A2(n_1033),
.B1(n_1024),
.B2(n_1034),
.C(n_962),
.Y(n_1110)
);

AOI31xp67_ASAP7_75t_L g1111 ( 
.A1(n_999),
.A2(n_988),
.A3(n_981),
.B(n_978),
.Y(n_1111)
);

AO31x2_ASAP7_75t_L g1112 ( 
.A1(n_964),
.A2(n_984),
.A3(n_1062),
.B(n_943),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_932),
.A2(n_972),
.B(n_1035),
.C(n_1038),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_969),
.Y(n_1114)
);

AO31x2_ASAP7_75t_L g1115 ( 
.A1(n_1028),
.A2(n_1060),
.A3(n_1022),
.B(n_961),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1011),
.A2(n_1042),
.B1(n_936),
.B2(n_995),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_954),
.B(n_1015),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_SL g1118 ( 
.A1(n_959),
.A2(n_1057),
.B(n_979),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1060),
.B(n_961),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_995),
.A2(n_961),
.B(n_953),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1022),
.A2(n_979),
.B(n_959),
.C(n_1057),
.Y(n_1121)
);

AO31x2_ASAP7_75t_L g1122 ( 
.A1(n_1060),
.A2(n_1040),
.A3(n_1057),
.B(n_954),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1054),
.A2(n_948),
.B1(n_1053),
.B2(n_1052),
.Y(n_1123)
);

INVx8_ASAP7_75t_L g1124 ( 
.A(n_1040),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1060),
.B(n_1040),
.Y(n_1125)
);

OA21x2_ASAP7_75t_L g1126 ( 
.A1(n_966),
.A2(n_949),
.B(n_990),
.Y(n_1126)
);

AOI221xp5_ASAP7_75t_SL g1127 ( 
.A1(n_1056),
.A2(n_844),
.B1(n_815),
.B2(n_832),
.C(n_950),
.Y(n_1127)
);

NOR2x1_ASAP7_75t_L g1128 ( 
.A(n_1052),
.B(n_1053),
.Y(n_1128)
);

AO31x2_ASAP7_75t_L g1129 ( 
.A1(n_1045),
.A2(n_752),
.A3(n_1059),
.B(n_1047),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1048),
.B(n_1002),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1013),
.A2(n_1006),
.B(n_990),
.Y(n_1131)
);

O2A1O1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_948),
.A2(n_1043),
.B(n_670),
.C(n_793),
.Y(n_1132)
);

NAND2xp33_ASAP7_75t_SL g1133 ( 
.A(n_955),
.B(n_989),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_SL g1134 ( 
.A1(n_1043),
.A2(n_993),
.B(n_873),
.C(n_900),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1043),
.A2(n_1048),
.B(n_1050),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_948),
.A2(n_1056),
.B1(n_612),
.B2(n_658),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1043),
.A2(n_1048),
.B(n_1050),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1045),
.A2(n_456),
.B(n_452),
.Y(n_1138)
);

BUFx10_ASAP7_75t_L g1139 ( 
.A(n_1052),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1041),
.B(n_458),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1045),
.A2(n_456),
.B(n_452),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1048),
.B(n_1002),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1013),
.A2(n_1006),
.B(n_990),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_948),
.A2(n_1043),
.B(n_670),
.C(n_793),
.Y(n_1144)
);

BUFx10_ASAP7_75t_L g1145 ( 
.A(n_1052),
.Y(n_1145)
);

AOI31xp67_ASAP7_75t_L g1146 ( 
.A1(n_1012),
.A2(n_1010),
.A3(n_939),
.B(n_968),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1013),
.A2(n_1006),
.B(n_990),
.Y(n_1147)
);

OA21x2_ASAP7_75t_L g1148 ( 
.A1(n_966),
.A2(n_949),
.B(n_990),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1048),
.B(n_1002),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1023),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1048),
.B(n_1002),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1048),
.B(n_1002),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_948),
.A2(n_1056),
.B1(n_612),
.B2(n_658),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1045),
.A2(n_456),
.B(n_452),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_948),
.A2(n_1052),
.B1(n_1061),
.B2(n_1053),
.Y(n_1155)
);

AO31x2_ASAP7_75t_L g1156 ( 
.A1(n_1045),
.A2(n_752),
.A3(n_1059),
.B(n_1047),
.Y(n_1156)
);

BUFx2_ASAP7_75t_SL g1157 ( 
.A(n_996),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_1045),
.A2(n_752),
.A3(n_1059),
.B(n_1047),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1048),
.B(n_1002),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1013),
.A2(n_1006),
.B(n_990),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1045),
.A2(n_456),
.B(n_452),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1046),
.B(n_781),
.Y(n_1162)
);

BUFx3_ASAP7_75t_L g1163 ( 
.A(n_1058),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1052),
.B(n_1053),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1043),
.A2(n_1048),
.B(n_1050),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1045),
.A2(n_456),
.B(n_452),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1041),
.B(n_458),
.Y(n_1167)
);

OR2x2_ASAP7_75t_L g1168 ( 
.A(n_1037),
.B(n_458),
.Y(n_1168)
);

AOI22x1_ASAP7_75t_L g1169 ( 
.A1(n_1021),
.A2(n_928),
.B1(n_1002),
.B2(n_1003),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1052),
.B(n_458),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_SL g1171 ( 
.A1(n_985),
.A2(n_752),
.B(n_970),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1041),
.B(n_458),
.Y(n_1172)
);

AOI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1013),
.A2(n_939),
.B(n_1045),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_991),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1052),
.B(n_458),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1048),
.B(n_1002),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1013),
.A2(n_1006),
.B(n_990),
.Y(n_1177)
);

BUFx10_ASAP7_75t_L g1178 ( 
.A(n_1052),
.Y(n_1178)
);

OR2x6_ASAP7_75t_L g1179 ( 
.A(n_980),
.B(n_653),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_1045),
.A2(n_752),
.A3(n_1059),
.B(n_1047),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_991),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1048),
.B(n_1002),
.Y(n_1182)
);

A2O1A1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_1043),
.A2(n_600),
.B(n_950),
.C(n_983),
.Y(n_1183)
);

BUFx8_ASAP7_75t_SL g1184 ( 
.A(n_946),
.Y(n_1184)
);

AO21x1_ASAP7_75t_L g1185 ( 
.A1(n_957),
.A2(n_985),
.B(n_1048),
.Y(n_1185)
);

NAND3xp33_ASAP7_75t_L g1186 ( 
.A(n_1056),
.B(n_670),
.C(n_793),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_991),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1052),
.B(n_458),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1013),
.A2(n_1006),
.B(n_990),
.Y(n_1189)
);

INVx1_ASAP7_75t_SL g1190 ( 
.A(n_1058),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1013),
.A2(n_1006),
.B(n_990),
.Y(n_1191)
);

AO31x2_ASAP7_75t_L g1192 ( 
.A1(n_1045),
.A2(n_752),
.A3(n_1059),
.B(n_1047),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1043),
.A2(n_600),
.B(n_950),
.C(n_983),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_933),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_SL g1195 ( 
.A1(n_1056),
.A2(n_385),
.B(n_549),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_948),
.A2(n_1052),
.B1(n_1061),
.B2(n_1053),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1045),
.A2(n_456),
.B(n_452),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1043),
.A2(n_600),
.B(n_950),
.C(n_983),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1023),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1045),
.A2(n_456),
.B(n_452),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_948),
.A2(n_1056),
.B1(n_612),
.B2(n_658),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1045),
.A2(n_456),
.B(n_452),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_SL g1203 ( 
.A1(n_1186),
.A2(n_1071),
.B1(n_1067),
.B2(n_1170),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1136),
.A2(n_1201),
.B1(n_1153),
.B2(n_1185),
.Y(n_1204)
);

OAI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1155),
.A2(n_1196),
.B1(n_1195),
.B2(n_1073),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1140),
.B(n_1167),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1072),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1099),
.Y(n_1208)
);

INVxp67_ASAP7_75t_SL g1209 ( 
.A(n_1094),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1190),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1135),
.A2(n_1137),
.B1(n_1165),
.B2(n_1086),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1184),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1070),
.A2(n_1105),
.B1(n_1077),
.B2(n_1095),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1066),
.A2(n_1128),
.B1(n_1188),
.B2(n_1175),
.Y(n_1214)
);

INVx4_ASAP7_75t_L g1215 ( 
.A(n_1124),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1106),
.Y(n_1216)
);

INVx1_ASAP7_75t_SL g1217 ( 
.A(n_1172),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1091),
.A2(n_1164),
.B1(n_1171),
.B2(n_1182),
.Y(n_1218)
);

INVx5_ASAP7_75t_L g1219 ( 
.A(n_1124),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_1084),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1123),
.A2(n_1127),
.B1(n_1093),
.B2(n_1082),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_SL g1222 ( 
.A1(n_1139),
.A2(n_1178),
.B1(n_1145),
.B2(n_1088),
.Y(n_1222)
);

BUFx10_ASAP7_75t_L g1223 ( 
.A(n_1103),
.Y(n_1223)
);

INVx4_ASAP7_75t_SL g1224 ( 
.A(n_1115),
.Y(n_1224)
);

OAI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1130),
.A2(n_1159),
.B1(n_1152),
.B2(n_1151),
.Y(n_1225)
);

INVx2_ASAP7_75t_SL g1226 ( 
.A(n_1163),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1142),
.A2(n_1149),
.B1(n_1176),
.B2(n_1107),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1098),
.A2(n_1097),
.B1(n_1100),
.B2(n_1169),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1090),
.A2(n_1139),
.B1(n_1145),
.B2(n_1178),
.Y(n_1229)
);

CKINVDCx16_ASAP7_75t_R g1230 ( 
.A(n_1069),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1194),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1069),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1065),
.A2(n_1181),
.B1(n_1187),
.B2(n_1174),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1114),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1168),
.B(n_1075),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1150),
.A2(n_1199),
.B1(n_1088),
.B2(n_1085),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1109),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_1087),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1199),
.A2(n_1109),
.B1(n_1083),
.B2(n_1162),
.Y(n_1239)
);

BUFx8_ASAP7_75t_SL g1240 ( 
.A(n_1102),
.Y(n_1240)
);

BUFx8_ASAP7_75t_L g1241 ( 
.A(n_1117),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1183),
.B(n_1193),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_SL g1243 ( 
.A1(n_1157),
.A2(n_1108),
.B1(n_1132),
.B2(n_1144),
.Y(n_1243)
);

BUFx4f_ASAP7_75t_SL g1244 ( 
.A(n_1162),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_SL g1245 ( 
.A1(n_1116),
.A2(n_1179),
.B1(n_1198),
.B2(n_1146),
.Y(n_1245)
);

CKINVDCx16_ASAP7_75t_R g1246 ( 
.A(n_1133),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1112),
.Y(n_1247)
);

INVx6_ASAP7_75t_L g1248 ( 
.A(n_1101),
.Y(n_1248)
);

INVx6_ASAP7_75t_L g1249 ( 
.A(n_1101),
.Y(n_1249)
);

CKINVDCx11_ASAP7_75t_R g1250 ( 
.A(n_1096),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1113),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1122),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1122),
.Y(n_1253)
);

AO22x1_ASAP7_75t_L g1254 ( 
.A1(n_1120),
.A2(n_1119),
.B1(n_1096),
.B2(n_1125),
.Y(n_1254)
);

INVx6_ASAP7_75t_L g1255 ( 
.A(n_1118),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1080),
.A2(n_1079),
.B1(n_1148),
.B2(n_1126),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1122),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1092),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_1078),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1076),
.Y(n_1260)
);

OAI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1068),
.A2(n_1081),
.B1(n_1110),
.B2(n_1173),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1104),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1148),
.A2(n_1089),
.B1(n_1202),
.B2(n_1141),
.Y(n_1263)
);

BUFx10_ASAP7_75t_L g1264 ( 
.A(n_1121),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_SL g1265 ( 
.A1(n_1089),
.A2(n_1134),
.B1(n_1074),
.B2(n_1200),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1089),
.Y(n_1266)
);

CKINVDCx14_ASAP7_75t_R g1267 ( 
.A(n_1129),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1129),
.Y(n_1268)
);

INVx4_ASAP7_75t_L g1269 ( 
.A(n_1131),
.Y(n_1269)
);

CKINVDCx11_ASAP7_75t_R g1270 ( 
.A(n_1129),
.Y(n_1270)
);

BUFx8_ASAP7_75t_L g1271 ( 
.A(n_1156),
.Y(n_1271)
);

AOI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1138),
.A2(n_1166),
.B1(n_1197),
.B2(n_1161),
.Y(n_1272)
);

CKINVDCx6p67_ASAP7_75t_R g1273 ( 
.A(n_1156),
.Y(n_1273)
);

CKINVDCx11_ASAP7_75t_R g1274 ( 
.A(n_1158),
.Y(n_1274)
);

INVxp67_ASAP7_75t_L g1275 ( 
.A(n_1143),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1154),
.A2(n_1177),
.B1(n_1147),
.B2(n_1191),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1158),
.A2(n_1180),
.B1(n_1192),
.B2(n_1160),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_SL g1278 ( 
.A1(n_1180),
.A2(n_1192),
.B(n_1189),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1192),
.A2(n_1071),
.B1(n_948),
.B2(n_1186),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1067),
.B(n_1091),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_1184),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1124),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1111),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1071),
.A2(n_948),
.B1(n_1186),
.B2(n_1056),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1071),
.A2(n_948),
.B1(n_1186),
.B2(n_1056),
.Y(n_1285)
);

CKINVDCx11_ASAP7_75t_R g1286 ( 
.A(n_1069),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1072),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1071),
.A2(n_948),
.B1(n_1186),
.B2(n_1056),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1072),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1071),
.A2(n_948),
.B1(n_1186),
.B2(n_1056),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_SL g1291 ( 
.A1(n_1067),
.A2(n_612),
.B1(n_1196),
.B2(n_1155),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_SL g1292 ( 
.A1(n_1195),
.A2(n_948),
.B(n_1056),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1071),
.A2(n_948),
.B1(n_1186),
.B2(n_1056),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1111),
.Y(n_1294)
);

INVx1_ASAP7_75t_SL g1295 ( 
.A(n_1190),
.Y(n_1295)
);

INVx1_ASAP7_75t_SL g1296 ( 
.A(n_1190),
.Y(n_1296)
);

BUFx12f_ASAP7_75t_L g1297 ( 
.A(n_1102),
.Y(n_1297)
);

INVx6_ASAP7_75t_L g1298 ( 
.A(n_1124),
.Y(n_1298)
);

OAI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1155),
.A2(n_793),
.B1(n_1196),
.B2(n_1186),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1072),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_1184),
.Y(n_1301)
);

CKINVDCx6p67_ASAP7_75t_R g1302 ( 
.A(n_1157),
.Y(n_1302)
);

INVx5_ASAP7_75t_L g1303 ( 
.A(n_1124),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_1163),
.Y(n_1304)
);

BUFx12f_ASAP7_75t_L g1305 ( 
.A(n_1102),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1071),
.A2(n_948),
.B1(n_1186),
.B2(n_1056),
.Y(n_1306)
);

BUFx2_ASAP7_75t_R g1307 ( 
.A(n_1184),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1067),
.B(n_1091),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1247),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1267),
.B(n_1266),
.Y(n_1310)
);

AND2x4_ASAP7_75t_L g1311 ( 
.A(n_1224),
.B(n_1253),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1264),
.Y(n_1312)
);

OA21x2_ASAP7_75t_L g1313 ( 
.A1(n_1278),
.A2(n_1294),
.B(n_1283),
.Y(n_1313)
);

INVx1_ASAP7_75t_SL g1314 ( 
.A(n_1210),
.Y(n_1314)
);

INVxp67_ASAP7_75t_SL g1315 ( 
.A(n_1260),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1211),
.A2(n_1242),
.B(n_1256),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1291),
.A2(n_1299),
.B1(n_1205),
.B2(n_1203),
.Y(n_1317)
);

AO21x2_ASAP7_75t_L g1318 ( 
.A1(n_1261),
.A2(n_1272),
.B(n_1277),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1264),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1252),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1257),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1256),
.A2(n_1228),
.B(n_1213),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1266),
.B(n_1268),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1213),
.B(n_1279),
.Y(n_1324)
);

INVx4_ASAP7_75t_L g1325 ( 
.A(n_1255),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1276),
.A2(n_1263),
.B(n_1258),
.Y(n_1326)
);

INVxp67_ASAP7_75t_L g1327 ( 
.A(n_1207),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1273),
.B(n_1270),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1262),
.B(n_1225),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1279),
.B(n_1270),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1271),
.Y(n_1331)
);

BUFx2_ASAP7_75t_L g1332 ( 
.A(n_1271),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_1241),
.Y(n_1333)
);

NOR2x1_ASAP7_75t_R g1334 ( 
.A(n_1286),
.B(n_1212),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1241),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1234),
.Y(n_1336)
);

OA21x2_ASAP7_75t_L g1337 ( 
.A1(n_1263),
.A2(n_1276),
.B(n_1228),
.Y(n_1337)
);

INVxp67_ASAP7_75t_L g1338 ( 
.A(n_1208),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_1301),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1227),
.B(n_1280),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1216),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1295),
.Y(n_1342)
);

AOI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1254),
.A2(n_1235),
.B(n_1251),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1224),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1269),
.Y(n_1345)
);

INVxp33_ASAP7_75t_L g1346 ( 
.A(n_1206),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1275),
.Y(n_1347)
);

AO21x1_ASAP7_75t_L g1348 ( 
.A1(n_1292),
.A2(n_1221),
.B(n_1231),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1224),
.Y(n_1349)
);

INVxp67_ASAP7_75t_L g1350 ( 
.A(n_1287),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1289),
.Y(n_1351)
);

INVx1_ASAP7_75t_SL g1352 ( 
.A(n_1296),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1218),
.B(n_1236),
.Y(n_1353)
);

INVx2_ASAP7_75t_SL g1354 ( 
.A(n_1255),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1300),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1274),
.Y(n_1356)
);

CKINVDCx16_ASAP7_75t_R g1357 ( 
.A(n_1230),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1265),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1236),
.B(n_1218),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1245),
.Y(n_1360)
);

OA21x2_ASAP7_75t_L g1361 ( 
.A1(n_1284),
.A2(n_1288),
.B(n_1306),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1284),
.B(n_1306),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1233),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1233),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1237),
.B(n_1239),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_1209),
.Y(n_1366)
);

AOI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1214),
.A2(n_1308),
.B(n_1293),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1285),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1239),
.A2(n_1288),
.B(n_1285),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1290),
.A2(n_1293),
.B(n_1204),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1317),
.A2(n_1290),
.B1(n_1204),
.B2(n_1243),
.Y(n_1371)
);

A2O1A1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1370),
.A2(n_1229),
.B(n_1222),
.C(n_1304),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_1312),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1310),
.B(n_1217),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1346),
.B(n_1223),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1340),
.B(n_1223),
.Y(n_1376)
);

O2A1O1Ixp33_ASAP7_75t_SL g1377 ( 
.A1(n_1368),
.A2(n_1226),
.B(n_1307),
.C(n_1286),
.Y(n_1377)
);

OAI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1370),
.A2(n_1232),
.B(n_1219),
.Y(n_1378)
);

NAND4xp25_ASAP7_75t_L g1379 ( 
.A(n_1340),
.B(n_1215),
.C(n_1282),
.D(n_1302),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1366),
.Y(n_1380)
);

AOI221xp5_ASAP7_75t_L g1381 ( 
.A1(n_1362),
.A2(n_1246),
.B1(n_1259),
.B2(n_1220),
.C(n_1238),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1366),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1318),
.B(n_1323),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1369),
.A2(n_1219),
.B(n_1303),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1342),
.B(n_1244),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1322),
.A2(n_1303),
.B(n_1248),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1318),
.B(n_1303),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1314),
.B(n_1362),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1369),
.A2(n_1281),
.B(n_1244),
.Y(n_1389)
);

AOI221xp5_ASAP7_75t_L g1390 ( 
.A1(n_1368),
.A2(n_1250),
.B1(n_1305),
.B2(n_1297),
.C(n_1240),
.Y(n_1390)
);

BUFx4f_ASAP7_75t_SL g1391 ( 
.A(n_1339),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1342),
.B(n_1297),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1355),
.Y(n_1393)
);

OA21x2_ASAP7_75t_L g1394 ( 
.A1(n_1326),
.A2(n_1250),
.B(n_1248),
.Y(n_1394)
);

OA21x2_ASAP7_75t_L g1395 ( 
.A1(n_1326),
.A2(n_1249),
.B(n_1298),
.Y(n_1395)
);

AO32x2_ASAP7_75t_L g1396 ( 
.A1(n_1354),
.A2(n_1298),
.A3(n_1355),
.B1(n_1325),
.B2(n_1348),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_SL g1397 ( 
.A1(n_1343),
.A2(n_1329),
.B(n_1367),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1352),
.B(n_1357),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_SL g1399 ( 
.A1(n_1361),
.A2(n_1357),
.B1(n_1356),
.B2(n_1360),
.Y(n_1399)
);

CKINVDCx11_ASAP7_75t_R g1400 ( 
.A(n_1333),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_1351),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1314),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1316),
.A2(n_1329),
.B(n_1318),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1361),
.B(n_1324),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1318),
.B(n_1347),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_SL g1406 ( 
.A1(n_1361),
.A2(n_1335),
.B1(n_1333),
.B2(n_1331),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1361),
.B(n_1324),
.Y(n_1407)
);

OA21x2_ASAP7_75t_L g1408 ( 
.A1(n_1309),
.A2(n_1315),
.B(n_1321),
.Y(n_1408)
);

AOI221xp5_ASAP7_75t_L g1409 ( 
.A1(n_1360),
.A2(n_1359),
.B1(n_1358),
.B2(n_1330),
.C(n_1364),
.Y(n_1409)
);

OR2x6_ASAP7_75t_L g1410 ( 
.A(n_1311),
.B(n_1344),
.Y(n_1410)
);

AOI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1361),
.A2(n_1330),
.B1(n_1359),
.B2(n_1365),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1320),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1412),
.Y(n_1413)
);

CKINVDCx20_ASAP7_75t_R g1414 ( 
.A(n_1391),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1383),
.B(n_1313),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1371),
.A2(n_1359),
.B1(n_1353),
.B2(n_1358),
.Y(n_1416)
);

INVxp67_ASAP7_75t_L g1417 ( 
.A(n_1380),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1408),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1405),
.B(n_1313),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1405),
.B(n_1313),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1404),
.B(n_1327),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1386),
.B(n_1367),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1383),
.B(n_1313),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1371),
.A2(n_1319),
.B1(n_1312),
.B2(n_1364),
.Y(n_1424)
);

AOI21xp33_ASAP7_75t_L g1425 ( 
.A1(n_1397),
.A2(n_1363),
.B(n_1337),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1410),
.B(n_1345),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1408),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1408),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1396),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1407),
.B(n_1327),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1376),
.B(n_1312),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1393),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1395),
.B(n_1337),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1401),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1403),
.B(n_1338),
.Y(n_1435)
);

INVx3_ASAP7_75t_R g1436 ( 
.A(n_1387),
.Y(n_1436)
);

INVx1_ASAP7_75t_SL g1437 ( 
.A(n_1434),
.Y(n_1437)
);

OAI33xp33_ASAP7_75t_L g1438 ( 
.A1(n_1435),
.A2(n_1399),
.A3(n_1388),
.B1(n_1406),
.B2(n_1350),
.B3(n_1341),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1413),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1419),
.B(n_1420),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1415),
.B(n_1382),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1419),
.B(n_1396),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1418),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1419),
.B(n_1396),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1421),
.B(n_1402),
.Y(n_1445)
);

NAND3xp33_ASAP7_75t_L g1446 ( 
.A(n_1416),
.B(n_1409),
.C(n_1372),
.Y(n_1446)
);

AOI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1416),
.A2(n_1424),
.B1(n_1399),
.B2(n_1411),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1413),
.Y(n_1448)
);

AOI33xp33_ASAP7_75t_L g1449 ( 
.A1(n_1424),
.A2(n_1411),
.A3(n_1352),
.B1(n_1390),
.B2(n_1374),
.B3(n_1377),
.Y(n_1449)
);

CKINVDCx20_ASAP7_75t_R g1450 ( 
.A(n_1414),
.Y(n_1450)
);

NOR2x1_ASAP7_75t_SL g1451 ( 
.A(n_1422),
.B(n_1410),
.Y(n_1451)
);

OR2x6_ASAP7_75t_L g1452 ( 
.A(n_1435),
.B(n_1384),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1420),
.B(n_1396),
.Y(n_1453)
);

OAI33xp33_ASAP7_75t_L g1454 ( 
.A1(n_1421),
.A2(n_1341),
.A3(n_1350),
.B1(n_1336),
.B2(n_1387),
.B3(n_1379),
.Y(n_1454)
);

OAI31xp33_ASAP7_75t_L g1455 ( 
.A1(n_1425),
.A2(n_1319),
.A3(n_1328),
.B(n_1331),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1420),
.B(n_1396),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1431),
.B(n_1319),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1423),
.B(n_1429),
.Y(n_1458)
);

AND4x1_ASAP7_75t_SL g1459 ( 
.A(n_1428),
.B(n_1381),
.C(n_1344),
.D(n_1349),
.Y(n_1459)
);

NOR2x1_ASAP7_75t_SL g1460 ( 
.A(n_1415),
.B(n_1410),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1434),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1426),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1415),
.B(n_1401),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1427),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1423),
.B(n_1394),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1439),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1439),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1442),
.B(n_1429),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1442),
.B(n_1429),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1445),
.B(n_1432),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1448),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1448),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1461),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1445),
.B(n_1432),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1441),
.B(n_1430),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1460),
.B(n_1462),
.Y(n_1476)
);

CKINVDCx16_ASAP7_75t_R g1477 ( 
.A(n_1450),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1441),
.B(n_1417),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1452),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1437),
.B(n_1417),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1443),
.Y(n_1481)
);

NOR4xp25_ASAP7_75t_SL g1482 ( 
.A(n_1451),
.B(n_1332),
.C(n_1436),
.D(n_1427),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1450),
.B(n_1414),
.Y(n_1483)
);

INVxp67_ASAP7_75t_L g1484 ( 
.A(n_1461),
.Y(n_1484)
);

INVx3_ASAP7_75t_L g1485 ( 
.A(n_1462),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1443),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1444),
.B(n_1433),
.Y(n_1487)
);

INVxp67_ASAP7_75t_L g1488 ( 
.A(n_1454),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1462),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1464),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1463),
.B(n_1427),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1468),
.B(n_1453),
.Y(n_1492)
);

NAND2x1p5_ASAP7_75t_L g1493 ( 
.A(n_1476),
.B(n_1394),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1466),
.Y(n_1494)
);

NAND2x1p5_ASAP7_75t_L g1495 ( 
.A(n_1476),
.B(n_1394),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1466),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1481),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1481),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1473),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1481),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1488),
.A2(n_1446),
.B1(n_1447),
.B2(n_1438),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1488),
.B(n_1484),
.Y(n_1502)
);

NOR4xp25_ASAP7_75t_L g1503 ( 
.A(n_1484),
.B(n_1446),
.C(n_1449),
.D(n_1398),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1476),
.Y(n_1504)
);

AOI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1477),
.A2(n_1447),
.B1(n_1438),
.B2(n_1454),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1467),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1486),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1468),
.B(n_1456),
.Y(n_1508)
);

INVxp33_ASAP7_75t_L g1509 ( 
.A(n_1483),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1467),
.Y(n_1510)
);

OAI21xp33_ASAP7_75t_L g1511 ( 
.A1(n_1470),
.A2(n_1449),
.B(n_1452),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1486),
.Y(n_1512)
);

NOR2x1p5_ASAP7_75t_L g1513 ( 
.A(n_1485),
.B(n_1333),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1471),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1471),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1473),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1468),
.B(n_1456),
.Y(n_1517)
);

OR2x6_ASAP7_75t_L g1518 ( 
.A(n_1479),
.B(n_1452),
.Y(n_1518)
);

NOR3xp33_ASAP7_75t_L g1519 ( 
.A(n_1477),
.B(n_1459),
.C(n_1392),
.Y(n_1519)
);

BUFx2_ASAP7_75t_SL g1520 ( 
.A(n_1476),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1469),
.B(n_1456),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1486),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1469),
.B(n_1460),
.Y(n_1523)
);

NAND2x1_ASAP7_75t_SL g1524 ( 
.A(n_1476),
.B(n_1465),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1470),
.B(n_1458),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1474),
.B(n_1458),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1491),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1472),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1469),
.B(n_1458),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1474),
.B(n_1440),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1472),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1475),
.B(n_1440),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1513),
.B(n_1479),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1501),
.B(n_1503),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1516),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1513),
.B(n_1451),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_1502),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1516),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1527),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1520),
.B(n_1485),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1494),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1503),
.B(n_1505),
.Y(n_1542)
);

INVx1_ASAP7_75t_SL g1543 ( 
.A(n_1509),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1494),
.Y(n_1544)
);

NAND4xp25_ASAP7_75t_L g1545 ( 
.A(n_1502),
.B(n_1455),
.C(n_1378),
.D(n_1335),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1525),
.B(n_1526),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1496),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1496),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1527),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1506),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1505),
.A2(n_1482),
.B1(n_1452),
.B2(n_1332),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1506),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1520),
.B(n_1485),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1510),
.Y(n_1554)
);

AOI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1511),
.A2(n_1452),
.B(n_1482),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1510),
.Y(n_1556)
);

NAND2x1p5_ASAP7_75t_L g1557 ( 
.A(n_1504),
.B(n_1373),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1511),
.B(n_1400),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1529),
.B(n_1485),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_L g1560 ( 
.A(n_1519),
.B(n_1334),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1514),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1519),
.B(n_1478),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1527),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1497),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1497),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1499),
.B(n_1478),
.Y(n_1566)
);

OAI21x1_ASAP7_75t_L g1567 ( 
.A1(n_1524),
.A2(n_1489),
.B(n_1485),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1543),
.B(n_1530),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1537),
.B(n_1530),
.Y(n_1569)
);

INVxp33_ASAP7_75t_L g1570 ( 
.A(n_1558),
.Y(n_1570)
);

AOI211xp5_ASAP7_75t_L g1571 ( 
.A1(n_1542),
.A2(n_1455),
.B(n_1523),
.C(n_1389),
.Y(n_1571)
);

NAND3xp33_ASAP7_75t_L g1572 ( 
.A(n_1534),
.B(n_1518),
.C(n_1452),
.Y(n_1572)
);

OAI211xp5_ASAP7_75t_L g1573 ( 
.A1(n_1555),
.A2(n_1524),
.B(n_1523),
.C(n_1504),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1541),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1541),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1562),
.B(n_1529),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1544),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1544),
.Y(n_1578)
);

OAI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1551),
.A2(n_1518),
.B(n_1452),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1547),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1547),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1548),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1560),
.B(n_1334),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1566),
.A2(n_1518),
.B1(n_1523),
.B2(n_1525),
.Y(n_1584)
);

OAI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1545),
.A2(n_1518),
.B1(n_1459),
.B2(n_1526),
.Y(n_1585)
);

INVxp67_ASAP7_75t_SL g1586 ( 
.A(n_1535),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1536),
.B(n_1529),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1548),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1545),
.A2(n_1518),
.B(n_1480),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1535),
.A2(n_1518),
.B(n_1480),
.Y(n_1590)
);

AOI211xp5_ASAP7_75t_L g1591 ( 
.A1(n_1536),
.A2(n_1504),
.B(n_1425),
.C(n_1431),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1540),
.Y(n_1592)
);

AND2x2_ASAP7_75t_SL g1593 ( 
.A(n_1583),
.B(n_1533),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1586),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1576),
.B(n_1538),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1587),
.B(n_1533),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1592),
.B(n_1538),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1568),
.B(n_1546),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1592),
.B(n_1546),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1587),
.B(n_1559),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1574),
.Y(n_1601)
);

AOI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1570),
.A2(n_1567),
.B(n_1553),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1570),
.A2(n_1567),
.B(n_1553),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1575),
.Y(n_1604)
);

OAI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1572),
.A2(n_1540),
.B(n_1550),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1583),
.B(n_1335),
.Y(n_1606)
);

AOI322xp5_ASAP7_75t_L g1607 ( 
.A1(n_1585),
.A2(n_1569),
.A3(n_1517),
.B1(n_1492),
.B2(n_1521),
.C1(n_1508),
.C2(n_1487),
.Y(n_1607)
);

AOI211xp5_ASAP7_75t_L g1608 ( 
.A1(n_1585),
.A2(n_1550),
.B(n_1552),
.C(n_1554),
.Y(n_1608)
);

AOI222xp33_ASAP7_75t_L g1609 ( 
.A1(n_1579),
.A2(n_1552),
.B1(n_1554),
.B2(n_1556),
.C1(n_1561),
.C2(n_1492),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1584),
.B(n_1532),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1577),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1594),
.B(n_1571),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1597),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1601),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1596),
.B(n_1559),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1593),
.B(n_1589),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1600),
.B(n_1590),
.Y(n_1617)
);

XNOR2xp5_ASAP7_75t_L g1618 ( 
.A(n_1608),
.B(n_1573),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1605),
.A2(n_1588),
.B1(n_1582),
.B2(n_1581),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1606),
.B(n_1578),
.Y(n_1620)
);

NAND2xp33_ASAP7_75t_SL g1621 ( 
.A(n_1598),
.B(n_1580),
.Y(n_1621)
);

AOI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1605),
.A2(n_1591),
.B(n_1561),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1618),
.B(n_1595),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1615),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1616),
.B(n_1595),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1614),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1620),
.B(n_1599),
.Y(n_1627)
);

NOR3xp33_ASAP7_75t_L g1628 ( 
.A(n_1612),
.B(n_1611),
.C(n_1604),
.Y(n_1628)
);

INVxp67_ASAP7_75t_L g1629 ( 
.A(n_1621),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1613),
.Y(n_1630)
);

OAI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1622),
.A2(n_1603),
.B(n_1602),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1620),
.Y(n_1632)
);

AOI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1631),
.A2(n_1619),
.B(n_1617),
.Y(n_1633)
);

NAND2xp33_ASAP7_75t_L g1634 ( 
.A(n_1625),
.B(n_1619),
.Y(n_1634)
);

OAI211xp5_ASAP7_75t_L g1635 ( 
.A1(n_1629),
.A2(n_1607),
.B(n_1609),
.C(n_1610),
.Y(n_1635)
);

OAI211xp5_ASAP7_75t_SL g1636 ( 
.A1(n_1623),
.A2(n_1609),
.B(n_1539),
.C(n_1549),
.Y(n_1636)
);

AOI221xp5_ASAP7_75t_L g1637 ( 
.A1(n_1629),
.A2(n_1556),
.B1(n_1563),
.B2(n_1539),
.C(n_1549),
.Y(n_1637)
);

AOI222xp33_ASAP7_75t_L g1638 ( 
.A1(n_1632),
.A2(n_1549),
.B1(n_1539),
.B2(n_1563),
.C1(n_1504),
.C2(n_1565),
.Y(n_1638)
);

NAND4xp25_ASAP7_75t_L g1639 ( 
.A(n_1633),
.B(n_1624),
.C(n_1628),
.D(n_1627),
.Y(n_1639)
);

NAND4xp75_ASAP7_75t_L g1640 ( 
.A(n_1637),
.B(n_1630),
.C(n_1626),
.D(n_1563),
.Y(n_1640)
);

OAI21xp33_ASAP7_75t_L g1641 ( 
.A1(n_1635),
.A2(n_1565),
.B(n_1564),
.Y(n_1641)
);

AOI211xp5_ASAP7_75t_L g1642 ( 
.A1(n_1634),
.A2(n_1565),
.B(n_1564),
.C(n_1385),
.Y(n_1642)
);

AOI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1636),
.A2(n_1564),
.B1(n_1495),
.B2(n_1493),
.Y(n_1643)
);

AOI221xp5_ASAP7_75t_L g1644 ( 
.A1(n_1638),
.A2(n_1557),
.B1(n_1498),
.B2(n_1500),
.C(n_1497),
.Y(n_1644)
);

AOI222xp33_ASAP7_75t_L g1645 ( 
.A1(n_1634),
.A2(n_1490),
.B1(n_1492),
.B2(n_1508),
.C1(n_1521),
.C2(n_1517),
.Y(n_1645)
);

AOI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1645),
.A2(n_1557),
.B1(n_1493),
.B2(n_1495),
.Y(n_1646)
);

NOR2xp67_ASAP7_75t_L g1647 ( 
.A(n_1639),
.B(n_1514),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1641),
.B(n_1515),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1640),
.Y(n_1649)
);

XNOR2xp5_ASAP7_75t_L g1650 ( 
.A(n_1642),
.B(n_1557),
.Y(n_1650)
);

NAND4xp25_ASAP7_75t_L g1651 ( 
.A(n_1647),
.B(n_1643),
.C(n_1644),
.D(n_1375),
.Y(n_1651)
);

NOR3xp33_ASAP7_75t_L g1652 ( 
.A(n_1649),
.B(n_1459),
.C(n_1457),
.Y(n_1652)
);

NOR3xp33_ASAP7_75t_L g1653 ( 
.A(n_1648),
.B(n_1650),
.C(n_1646),
.Y(n_1653)
);

XNOR2x1_ASAP7_75t_L g1654 ( 
.A(n_1653),
.B(n_1493),
.Y(n_1654)
);

AOI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1654),
.A2(n_1651),
.B1(n_1652),
.B2(n_1512),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1655),
.A2(n_1498),
.B1(n_1507),
.B2(n_1512),
.Y(n_1656)
);

XNOR2xp5_ASAP7_75t_L g1657 ( 
.A(n_1655),
.B(n_1493),
.Y(n_1657)
);

NAND3xp33_ASAP7_75t_L g1658 ( 
.A(n_1657),
.B(n_1500),
.C(n_1498),
.Y(n_1658)
);

AOI22x1_ASAP7_75t_L g1659 ( 
.A1(n_1656),
.A2(n_1507),
.B1(n_1512),
.B2(n_1522),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1659),
.A2(n_1500),
.B1(n_1507),
.B2(n_1522),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1658),
.A2(n_1522),
.B1(n_1515),
.B2(n_1531),
.Y(n_1661)
);

OAI22xp5_ASAP7_75t_SL g1662 ( 
.A1(n_1660),
.A2(n_1495),
.B1(n_1528),
.B2(n_1531),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1662),
.B(n_1661),
.Y(n_1663)
);

BUFx4_ASAP7_75t_R g1664 ( 
.A(n_1663),
.Y(n_1664)
);

AOI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1664),
.A2(n_1528),
.B1(n_1490),
.B2(n_1489),
.C(n_1532),
.Y(n_1665)
);

AOI211xp5_ASAP7_75t_L g1666 ( 
.A1(n_1665),
.A2(n_1457),
.B(n_1373),
.C(n_1517),
.Y(n_1666)
);


endmodule