module fake_netlist_5_1478_n_1956 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1956);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1956;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_604;
wire n_368;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_968;
wire n_912;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_108),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_29),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_65),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_44),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_120),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_107),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_31),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_33),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_81),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_38),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_139),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_176),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_2),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_43),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_104),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_154),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_88),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_150),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_63),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_70),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_192),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_158),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_89),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_43),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_168),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_86),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_27),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_105),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_92),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_82),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_170),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_5),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_44),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_119),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_145),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_67),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_11),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_130),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_69),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_78),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_166),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_28),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_162),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_103),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_171),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_47),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_156),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_99),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_51),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_73),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_72),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_93),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_134),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_102),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_132),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_76),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_32),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_84),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_109),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_33),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_17),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_185),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_14),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_2),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_153),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_151),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_125),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_143),
.Y(n_264)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_138),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_49),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_110),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_135),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_144),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_121),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_51),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_28),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_172),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_21),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_163),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_95),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_52),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_189),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_24),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_4),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_101),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_50),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_83),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_57),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_40),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_53),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_39),
.Y(n_287)
);

INVx2_ASAP7_75t_SL g288 ( 
.A(n_173),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_142),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_169),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_57),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_165),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_129),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_112),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_16),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_5),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_48),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_148),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_98),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_37),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_175),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_32),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_13),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_113),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_45),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_75),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_118),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_123),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_56),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_116),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_180),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_9),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_133),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_37),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_27),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_179),
.Y(n_316)
);

BUFx10_ASAP7_75t_L g317 ( 
.A(n_96),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_14),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_62),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_87),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_167),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_61),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_10),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_111),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_186),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_97),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_114),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_48),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_190),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_1),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_26),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_71),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_91),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_60),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_9),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_94),
.Y(n_336)
);

INVxp33_ASAP7_75t_L g337 ( 
.A(n_19),
.Y(n_337)
);

BUFx10_ASAP7_75t_L g338 ( 
.A(n_140),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_174),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_115),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_152),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_21),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_124),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_45),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_58),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_20),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_10),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_22),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_188),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_187),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_39),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_137),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_41),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_63),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_13),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_54),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_183),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_100),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_30),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_177),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_60),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_79),
.Y(n_362)
);

BUFx5_ASAP7_75t_L g363 ( 
.A(n_55),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_126),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_191),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_127),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_20),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_74),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_4),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_38),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_8),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_122),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_53),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_0),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_160),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_68),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_117),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_22),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_146),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_131),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_46),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_61),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_106),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_6),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_181),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_363),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_241),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_198),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_322),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_363),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_267),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_273),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_363),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_236),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_363),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_255),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_237),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_363),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_226),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_346),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_307),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_363),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_329),
.Y(n_403)
);

BUFx10_ASAP7_75t_L g404 ( 
.A(n_280),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_363),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_240),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_226),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_319),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_319),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_339),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_319),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_243),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_319),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_305),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_319),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_384),
.Y(n_416)
);

INVxp33_ASAP7_75t_SL g417 ( 
.A(n_202),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_384),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_384),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_305),
.Y(n_420)
);

INVxp33_ASAP7_75t_SL g421 ( 
.A(n_202),
.Y(n_421)
);

INVxp33_ASAP7_75t_SL g422 ( 
.A(n_204),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_345),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_349),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_231),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_294),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_321),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_244),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_323),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_246),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_323),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_254),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_263),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_384),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_204),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_384),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_276),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_268),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_270),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_201),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_278),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_265),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_374),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_374),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_378),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_378),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_228),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_207),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_229),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_276),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_281),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_276),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_233),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_259),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_283),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_299),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_271),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_272),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_291),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_297),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_314),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g462 ( 
.A(n_308),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_306),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_315),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_328),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_311),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_313),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_316),
.Y(n_468)
);

INVxp33_ASAP7_75t_L g469 ( 
.A(n_337),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_344),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_347),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_354),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_326),
.Y(n_473)
);

INVxp33_ASAP7_75t_SL g474 ( 
.A(n_207),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_359),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_308),
.Y(n_476)
);

INVxp33_ASAP7_75t_SL g477 ( 
.A(n_209),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_369),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_373),
.Y(n_479)
);

CKINVDCx14_ASAP7_75t_R g480 ( 
.A(n_317),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_209),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_386),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_425),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_408),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_408),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_409),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_390),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_481),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_409),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_399),
.B(n_239),
.Y(n_490)
);

AND2x2_ASAP7_75t_SL g491 ( 
.A(n_437),
.B(n_211),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_462),
.B(n_436),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_407),
.B(n_325),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_411),
.B(n_239),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_411),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_413),
.Y(n_496)
);

AND2x6_ASAP7_75t_L g497 ( 
.A(n_390),
.B(n_205),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_469),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_388),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_394),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_442),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_397),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_393),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_442),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_393),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_400),
.A2(n_282),
.B1(n_361),
.B2(n_257),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_448),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_413),
.B(n_250),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_417),
.B(n_250),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_395),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_395),
.Y(n_511)
);

CKINVDCx16_ASAP7_75t_R g512 ( 
.A(n_423),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_406),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_412),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_414),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_387),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_398),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_398),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_402),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_402),
.Y(n_520)
);

NOR2x1_ASAP7_75t_L g521 ( 
.A(n_415),
.B(n_325),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_450),
.B(n_317),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_405),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_428),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_405),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_415),
.Y(n_526)
);

AND3x2_ASAP7_75t_L g527 ( 
.A(n_435),
.B(n_330),
.C(n_215),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_416),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_416),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_418),
.B(n_288),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_418),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_419),
.B(n_362),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_419),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_426),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_434),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_434),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_449),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_443),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_443),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_449),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_453),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_407),
.B(n_288),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_453),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_457),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_444),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_457),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_458),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_430),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_389),
.A2(n_334),
.B1(n_382),
.B2(n_381),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_458),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_414),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_444),
.Y(n_552)
);

INVx6_ASAP7_75t_L g553 ( 
.A(n_476),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_459),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_391),
.B(n_214),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_459),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_445),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_445),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_460),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_392),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_509),
.B(n_432),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_487),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_516),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_505),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_498),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_487),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_526),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_526),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_509),
.B(n_433),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_499),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_498),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_526),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_487),
.Y(n_573)
);

BUFx4f_ASAP7_75t_L g574 ( 
.A(n_505),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_533),
.Y(n_575)
);

AND3x2_ASAP7_75t_L g576 ( 
.A(n_507),
.B(n_215),
.C(n_211),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_553),
.B(n_438),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_553),
.Y(n_578)
);

INVxp33_ASAP7_75t_SL g579 ( 
.A(n_555),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_553),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_491),
.B(n_452),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_533),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_533),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_503),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_505),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_505),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_501),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_553),
.B(n_439),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_501),
.Y(n_589)
);

AO21x2_ASAP7_75t_L g590 ( 
.A1(n_490),
.A2(n_197),
.B(n_195),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_553),
.B(n_441),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_503),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_553),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_506),
.B(n_401),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_491),
.B(n_455),
.Y(n_595)
);

BUFx10_ASAP7_75t_L g596 ( 
.A(n_500),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_491),
.B(n_456),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_503),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_493),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_511),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_511),
.Y(n_601)
);

INVxp67_ASAP7_75t_SL g602 ( 
.A(n_492),
.Y(n_602)
);

CKINVDCx6p67_ASAP7_75t_R g603 ( 
.A(n_512),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_532),
.B(n_362),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_511),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_501),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_501),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_520),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_501),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_504),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_502),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_505),
.Y(n_612)
);

OR2x6_ASAP7_75t_L g613 ( 
.A(n_542),
.B(n_227),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_513),
.B(n_463),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_549),
.A2(n_396),
.B1(n_488),
.B2(n_506),
.Y(n_615)
);

INVx5_ASAP7_75t_L g616 ( 
.A(n_497),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_505),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_532),
.B(n_466),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_520),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_514),
.B(n_467),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_532),
.B(n_480),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_493),
.B(n_476),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_504),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_SL g624 ( 
.A(n_512),
.B(n_427),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_520),
.Y(n_625)
);

OAI22xp33_ASAP7_75t_SL g626 ( 
.A1(n_490),
.A2(n_422),
.B1(n_474),
.B2(n_421),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_504),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_525),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_493),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_555),
.Y(n_630)
);

BUFx6f_ASAP7_75t_SL g631 ( 
.A(n_532),
.Y(n_631)
);

CKINVDCx16_ASAP7_75t_R g632 ( 
.A(n_560),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_524),
.B(n_477),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_525),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_505),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_517),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_504),
.Y(n_637)
);

INVx5_ASAP7_75t_L g638 ( 
.A(n_497),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_525),
.Y(n_639)
);

NOR2x1p5_ASAP7_75t_L g640 ( 
.A(n_548),
.B(n_214),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_517),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_532),
.B(n_327),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_510),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_517),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_510),
.B(n_333),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_483),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_510),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_510),
.Y(n_648)
);

OR2x2_ASAP7_75t_L g649 ( 
.A(n_515),
.B(n_435),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_482),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_518),
.A2(n_279),
.B1(n_227),
.B2(n_379),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_518),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_518),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_482),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_517),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_518),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_504),
.Y(n_657)
);

AND3x2_ASAP7_75t_L g658 ( 
.A(n_507),
.B(n_376),
.C(n_340),
.Y(n_658)
);

BUFx6f_ASAP7_75t_SL g659 ( 
.A(n_537),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_492),
.B(n_429),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_542),
.B(n_537),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_540),
.B(n_541),
.Y(n_662)
);

AOI21x1_ASAP7_75t_L g663 ( 
.A1(n_494),
.A2(n_376),
.B(n_340),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_488),
.B(n_451),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_523),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_515),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_549),
.A2(n_277),
.B1(n_253),
.B2(n_219),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_522),
.B(n_468),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_482),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_SL g670 ( 
.A1(n_551),
.A2(n_424),
.B1(n_403),
.B2(n_410),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_484),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_523),
.Y(n_672)
);

BUFx10_ASAP7_75t_L g673 ( 
.A(n_551),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_523),
.Y(n_674)
);

OAI22xp33_ASAP7_75t_L g675 ( 
.A1(n_522),
.A2(n_256),
.B1(n_287),
.B2(n_286),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_527),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_540),
.B(n_473),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_541),
.B(n_431),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_484),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_485),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_523),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_517),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_517),
.B(n_336),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_485),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_536),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_543),
.B(n_404),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_536),
.Y(n_687)
);

INVxp33_ASAP7_75t_L g688 ( 
.A(n_483),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_536),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_486),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_486),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_536),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_527),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_543),
.B(n_404),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_544),
.B(n_404),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_544),
.B(n_420),
.Y(n_696)
);

OAI21xp33_ASAP7_75t_SL g697 ( 
.A1(n_546),
.A2(n_279),
.B(n_547),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_517),
.B(n_519),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_489),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_519),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_519),
.B(n_350),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_534),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_546),
.B(n_317),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_489),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_495),
.Y(n_705)
);

AND2x2_ASAP7_75t_SL g706 ( 
.A(n_519),
.B(n_379),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_495),
.Y(n_707)
);

AO22x2_ASAP7_75t_L g708 ( 
.A1(n_494),
.A2(n_247),
.B1(n_199),
.B2(n_203),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_496),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_496),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_547),
.B(n_420),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_519),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_587),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_602),
.B(n_519),
.Y(n_714)
);

HB1xp67_ASAP7_75t_L g715 ( 
.A(n_571),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_662),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_587),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_571),
.B(n_193),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_662),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_587),
.Y(n_720)
);

OAI22xp5_ASAP7_75t_L g721 ( 
.A1(n_599),
.A2(n_298),
.B1(n_221),
.B2(n_220),
.Y(n_721)
);

NOR3xp33_ASAP7_75t_L g722 ( 
.A(n_626),
.B(n_454),
.C(n_447),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_661),
.B(n_519),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_678),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_569),
.B(n_193),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_589),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_565),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_599),
.B(n_528),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_561),
.B(n_200),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_696),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_629),
.B(n_529),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_589),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_570),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_678),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_629),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_706),
.B(n_529),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_589),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_595),
.A2(n_264),
.B1(n_208),
.B2(n_217),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_597),
.B(n_200),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_684),
.Y(n_740)
);

BUFx5_ASAP7_75t_L g741 ( 
.A(n_672),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_706),
.B(n_531),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_684),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_649),
.B(n_666),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_673),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_675),
.B(n_206),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_706),
.B(n_531),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_695),
.B(n_622),
.Y(n_748)
);

NAND2xp33_ASAP7_75t_L g749 ( 
.A(n_618),
.B(n_265),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_SL g750 ( 
.A(n_611),
.B(n_596),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_581),
.B(n_206),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_606),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_660),
.B(n_690),
.Y(n_753)
);

INVx4_ASAP7_75t_L g754 ( 
.A(n_631),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_606),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_691),
.B(n_539),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_622),
.B(n_626),
.Y(n_757)
);

NOR3xp33_ASAP7_75t_L g758 ( 
.A(n_677),
.B(n_475),
.C(n_234),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_649),
.B(n_534),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_642),
.B(n_676),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_606),
.Y(n_761)
);

NOR2x1p5_ASAP7_75t_L g762 ( 
.A(n_603),
.B(n_219),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_676),
.B(n_210),
.Y(n_763)
);

INVx6_ASAP7_75t_L g764 ( 
.A(n_673),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_691),
.B(n_704),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_SL g766 ( 
.A1(n_594),
.A2(n_223),
.B1(n_367),
.B2(n_370),
.Y(n_766)
);

NAND2xp33_ASAP7_75t_SL g767 ( 
.A(n_659),
.B(n_223),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_704),
.B(n_539),
.Y(n_768)
);

NOR3xp33_ASAP7_75t_L g769 ( 
.A(n_697),
.B(n_235),
.C(n_232),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_671),
.Y(n_770)
);

INVxp67_ASAP7_75t_SL g771 ( 
.A(n_598),
.Y(n_771)
);

OAI221xp5_ASAP7_75t_L g772 ( 
.A1(n_697),
.A2(n_651),
.B1(n_615),
.B2(n_667),
.C(n_711),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_620),
.B(n_210),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_693),
.B(n_212),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_672),
.B(n_539),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_673),
.Y(n_776)
);

NOR2x1p5_ASAP7_75t_L g777 ( 
.A(n_603),
.B(n_367),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_604),
.B(n_550),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_607),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_607),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_609),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_621),
.B(n_212),
.Y(n_782)
);

NAND3xp33_ASAP7_75t_L g783 ( 
.A(n_668),
.B(n_196),
.C(n_194),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_693),
.B(n_213),
.Y(n_784)
);

NOR3xp33_ASAP7_75t_L g785 ( 
.A(n_664),
.B(n_251),
.C(n_248),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_674),
.B(n_558),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_SL g787 ( 
.A(n_596),
.B(n_338),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_643),
.A2(n_252),
.B(n_324),
.C(n_332),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_614),
.B(n_686),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_671),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_673),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_694),
.B(n_213),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_679),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_679),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_680),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_680),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_699),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_604),
.B(n_550),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_699),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_596),
.B(n_216),
.Y(n_800)
);

OAI221xp5_ASAP7_75t_L g801 ( 
.A1(n_615),
.A2(n_559),
.B1(n_556),
.B2(n_554),
.C(n_530),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_666),
.B(n_559),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_681),
.B(n_558),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_604),
.A2(n_352),
.B1(n_521),
.B2(n_222),
.Y(n_804)
);

OAI22xp33_ASAP7_75t_L g805 ( 
.A1(n_667),
.A2(n_370),
.B1(n_371),
.B2(n_381),
.Y(n_805)
);

NOR2xp67_ASAP7_75t_L g806 ( 
.A(n_702),
.B(n_554),
.Y(n_806)
);

OR2x6_ASAP7_75t_L g807 ( 
.A(n_670),
.B(n_440),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_646),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_596),
.B(n_216),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_643),
.B(n_552),
.Y(n_810)
);

A2O1A1Ixp33_ASAP7_75t_SL g811 ( 
.A1(n_647),
.A2(n_365),
.B(n_377),
.C(n_375),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_647),
.B(n_552),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_630),
.B(n_556),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_648),
.B(n_552),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_604),
.B(n_460),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_648),
.B(n_552),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_652),
.B(n_508),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_633),
.B(n_218),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_610),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_652),
.B(n_653),
.Y(n_820)
);

NAND3xp33_ASAP7_75t_L g821 ( 
.A(n_703),
.B(n_242),
.C(n_238),
.Y(n_821)
);

NAND2xp33_ASAP7_75t_L g822 ( 
.A(n_577),
.B(n_265),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_613),
.A2(n_262),
.B1(n_275),
.B2(n_289),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_653),
.B(n_508),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_656),
.B(n_530),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_640),
.B(n_461),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_665),
.B(n_205),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_588),
.B(n_591),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_656),
.B(n_521),
.Y(n_829)
);

NAND2xp33_ASAP7_75t_L g830 ( 
.A(n_645),
.B(n_265),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_659),
.B(n_218),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_665),
.B(n_535),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_590),
.A2(n_205),
.B1(n_320),
.B2(n_269),
.Y(n_833)
);

OAI22xp33_ASAP7_75t_L g834 ( 
.A1(n_613),
.A2(n_371),
.B1(n_382),
.B2(n_335),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_624),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_576),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_705),
.B(n_222),
.Y(n_837)
);

INVx8_ASAP7_75t_L g838 ( 
.A(n_659),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_665),
.B(n_224),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_590),
.B(n_535),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_590),
.B(n_535),
.Y(n_841)
);

O2A1O1Ixp5_ASAP7_75t_L g842 ( 
.A1(n_683),
.A2(n_301),
.B(n_304),
.C(n_310),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_705),
.Y(n_843)
);

AO22x2_ASAP7_75t_L g844 ( 
.A1(n_708),
.A2(n_290),
.B1(n_292),
.B2(n_341),
.Y(n_844)
);

INVx5_ASAP7_75t_L g845 ( 
.A(n_617),
.Y(n_845)
);

BUFx5_ASAP7_75t_L g846 ( 
.A(n_700),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_707),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_708),
.A2(n_205),
.B1(n_269),
.B2(n_249),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_707),
.B(n_224),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_L g850 ( 
.A(n_578),
.B(n_265),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_613),
.A2(n_230),
.B1(n_225),
.B2(n_293),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_670),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_623),
.Y(n_853)
);

BUFx4f_ASAP7_75t_L g854 ( 
.A(n_613),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_613),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_709),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_709),
.B(n_225),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_710),
.B(n_230),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_640),
.B(n_461),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_623),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_710),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_701),
.B(n_293),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_564),
.B(n_535),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_564),
.B(n_535),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_708),
.A2(n_205),
.B1(n_269),
.B2(n_261),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_564),
.B(n_535),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_564),
.B(n_535),
.Y(n_867)
);

OA21x2_ASAP7_75t_L g868 ( 
.A1(n_685),
.A2(n_357),
.B(n_364),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_585),
.B(n_497),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_700),
.Y(n_870)
);

INVxp67_ASAP7_75t_L g871 ( 
.A(n_708),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_729),
.B(n_562),
.Y(n_872)
);

NOR2x1_ASAP7_75t_L g873 ( 
.A(n_754),
.B(n_563),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_770),
.Y(n_874)
);

OAI21xp5_ASAP7_75t_L g875 ( 
.A1(n_723),
.A2(n_698),
.B(n_574),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_715),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_790),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_715),
.B(n_688),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_729),
.B(n_562),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_793),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_725),
.B(n_566),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_794),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_753),
.B(n_616),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_730),
.B(n_594),
.Y(n_884)
);

AND2x4_ASAP7_75t_SL g885 ( 
.A(n_754),
.B(n_338),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_795),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_725),
.B(n_566),
.Y(n_887)
);

HB1xp67_ASAP7_75t_L g888 ( 
.A(n_744),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_796),
.Y(n_889)
);

INVxp67_ASAP7_75t_L g890 ( 
.A(n_760),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_714),
.A2(n_574),
.B(n_578),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_733),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_730),
.B(n_760),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_802),
.B(n_632),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_740),
.B(n_573),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_727),
.B(n_632),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_870),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_797),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_799),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_789),
.A2(n_631),
.B1(n_580),
.B2(n_593),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_843),
.Y(n_901)
);

NOR2xp67_ASAP7_75t_L g902 ( 
.A(n_727),
.B(n_663),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_743),
.B(n_584),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_772),
.B(n_585),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_870),
.Y(n_905)
);

NOR2xp67_ASAP7_75t_L g906 ( 
.A(n_783),
.B(n_663),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_735),
.B(n_592),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_765),
.B(n_592),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_808),
.Y(n_909)
);

BUFx4f_ASAP7_75t_L g910 ( 
.A(n_838),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_813),
.Y(n_911)
);

INVxp67_ASAP7_75t_L g912 ( 
.A(n_826),
.Y(n_912)
);

OR2x6_ASAP7_75t_L g913 ( 
.A(n_838),
.B(n_464),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_847),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_716),
.B(n_658),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_848),
.A2(n_631),
.B1(n_654),
.B2(n_669),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_719),
.B(n_600),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_838),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_856),
.Y(n_919)
);

NAND3xp33_ASAP7_75t_L g920 ( 
.A(n_739),
.B(n_260),
.C(n_245),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_SL g921 ( 
.A(n_750),
.B(n_579),
.Y(n_921)
);

AO22x1_ASAP7_75t_L g922 ( 
.A1(n_739),
.A2(n_342),
.B1(n_356),
.B2(n_331),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_862),
.B(n_600),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_833),
.A2(n_593),
.B1(n_580),
.B2(n_574),
.Y(n_924)
);

BUFx4f_ASAP7_75t_SL g925 ( 
.A(n_759),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_861),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_815),
.B(n_464),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_836),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_778),
.Y(n_929)
);

INVx2_ASAP7_75t_SL g930 ( 
.A(n_859),
.Y(n_930)
);

CKINVDCx11_ASAP7_75t_R g931 ( 
.A(n_807),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_724),
.B(n_465),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_778),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_848),
.A2(n_669),
.B1(n_650),
.B2(n_654),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_741),
.B(n_854),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_801),
.B(n_585),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_865),
.A2(n_650),
.B1(n_605),
.B2(n_608),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_862),
.B(n_605),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_865),
.A2(n_625),
.B1(n_608),
.B2(n_619),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_713),
.Y(n_940)
);

INVxp67_ASAP7_75t_L g941 ( 
.A(n_748),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_815),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_798),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_764),
.Y(n_944)
);

INVxp67_ASAP7_75t_L g945 ( 
.A(n_763),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_717),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_741),
.B(n_616),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_828),
.A2(n_636),
.B(n_635),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_R g949 ( 
.A(n_767),
.B(n_358),
.Y(n_949)
);

INVxp67_ASAP7_75t_L g950 ( 
.A(n_763),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_720),
.Y(n_951)
);

NOR3xp33_ASAP7_75t_SL g952 ( 
.A(n_805),
.B(n_274),
.C(n_266),
.Y(n_952)
);

OR2x6_ASAP7_75t_L g953 ( 
.A(n_764),
.B(n_465),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_833),
.A2(n_687),
.B1(n_685),
.B2(n_692),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_798),
.B(n_470),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_726),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_820),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_870),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_771),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_732),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_855),
.Y(n_961)
);

AND2x6_ASAP7_75t_L g962 ( 
.A(n_840),
.B(n_685),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_835),
.B(n_585),
.Y(n_963)
);

INVx5_ASAP7_75t_L g964 ( 
.A(n_870),
.Y(n_964)
);

INVx5_ASAP7_75t_L g965 ( 
.A(n_845),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_771),
.Y(n_966)
);

INVx4_ASAP7_75t_L g967 ( 
.A(n_764),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_835),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_R g969 ( 
.A(n_745),
.B(n_358),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_734),
.B(n_470),
.Y(n_970)
);

OR2x2_ASAP7_75t_L g971 ( 
.A(n_718),
.B(n_471),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_728),
.B(n_731),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_736),
.A2(n_692),
.B1(n_689),
.B2(n_687),
.Y(n_973)
);

NOR2x2_ASAP7_75t_L g974 ( 
.A(n_807),
.B(n_338),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_756),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_774),
.B(n_586),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_737),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_817),
.B(n_619),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_806),
.B(n_471),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_776),
.B(n_472),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_824),
.B(n_625),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_825),
.B(n_586),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_768),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_774),
.B(n_784),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_752),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_810),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_845),
.A2(n_635),
.B(n_636),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_858),
.B(n_586),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_784),
.B(n_472),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_812),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_814),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_858),
.B(n_586),
.Y(n_992)
);

NAND2xp33_ASAP7_75t_L g993 ( 
.A(n_846),
.B(n_616),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_755),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_741),
.B(n_616),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_757),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_741),
.B(n_638),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_871),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_751),
.A2(n_712),
.B1(n_700),
.B2(n_612),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_844),
.A2(n_265),
.B1(n_598),
.B2(n_601),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_839),
.B(n_612),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_761),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_845),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_791),
.B(n_478),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_839),
.B(n_751),
.Y(n_1005)
);

INVx5_ASAP7_75t_L g1006 ( 
.A(n_845),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_741),
.B(n_638),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_816),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_741),
.B(n_612),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_807),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_871),
.Y(n_1011)
);

INVx1_ASAP7_75t_SL g1012 ( 
.A(n_766),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_775),
.Y(n_1013)
);

BUFx12f_ASAP7_75t_L g1014 ( 
.A(n_762),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_854),
.B(n_638),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_844),
.A2(n_265),
.B1(n_601),
.B2(n_628),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_742),
.B(n_612),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_844),
.A2(n_628),
.B1(n_634),
.B2(n_639),
.Y(n_1018)
);

AOI22x1_ASAP7_75t_L g1019 ( 
.A1(n_779),
.A2(n_692),
.B1(n_689),
.B2(n_687),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_747),
.B(n_641),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_R g1021 ( 
.A(n_787),
.B(n_360),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_780),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_786),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_R g1024 ( 
.A(n_749),
.B(n_360),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_829),
.B(n_641),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_832),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_834),
.B(n_638),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_846),
.B(n_638),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_841),
.A2(n_635),
.B(n_636),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_792),
.B(n_641),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_781),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_792),
.B(n_641),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_803),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_773),
.B(n_655),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_831),
.Y(n_1035)
);

NOR3xp33_ASAP7_75t_L g1036 ( 
.A(n_805),
.B(n_385),
.C(n_368),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_868),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_819),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_846),
.B(n_655),
.Y(n_1039)
);

INVx4_ASAP7_75t_L g1040 ( 
.A(n_846),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_834),
.B(n_638),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_853),
.Y(n_1042)
);

INVx2_ASAP7_75t_SL g1043 ( 
.A(n_777),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_860),
.Y(n_1044)
);

AND2x6_ASAP7_75t_SL g1045 ( 
.A(n_831),
.B(n_478),
.Y(n_1045)
);

INVx1_ASAP7_75t_SL g1046 ( 
.A(n_818),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_821),
.B(n_479),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_746),
.B(n_655),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_868),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_800),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_904),
.A2(n_842),
.B(n_869),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_897),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_998),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_984),
.B(n_738),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_878),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_984),
.A2(n_852),
.B1(n_851),
.B2(n_804),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_888),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_888),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_897),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_945),
.B(n_852),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_R g1061 ( 
.A(n_892),
.B(n_822),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_1005),
.A2(n_945),
.B(n_950),
.C(n_893),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_916),
.A2(n_785),
.B1(n_758),
.B2(n_721),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_1040),
.A2(n_635),
.B(n_636),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_998),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1011),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_950),
.A2(n_782),
.B(n_785),
.C(n_722),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_890),
.B(n_809),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_1036),
.A2(n_758),
.B1(n_823),
.B2(n_769),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_965),
.A2(n_712),
.B(n_867),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_972),
.B(n_769),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_957),
.B(n_890),
.Y(n_1072)
);

NOR3xp33_ASAP7_75t_SL g1073 ( 
.A(n_968),
.B(n_285),
.C(n_295),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1011),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_918),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_965),
.A2(n_712),
.B(n_866),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_996),
.A2(n_722),
.B(n_837),
.C(n_857),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_965),
.A2(n_864),
.B(n_863),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_884),
.A2(n_849),
.B1(n_830),
.B2(n_850),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_904),
.A2(n_827),
.B(n_343),
.C(n_366),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_930),
.B(n_846),
.Y(n_1081)
);

NOR2xp67_ASAP7_75t_L g1082 ( 
.A(n_911),
.B(n_827),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_1006),
.A2(n_617),
.B(n_644),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_884),
.B(n_655),
.Y(n_1084)
);

OAI221xp5_ASAP7_75t_L g1085 ( 
.A1(n_1036),
.A2(n_318),
.B1(n_355),
.B2(n_353),
.C(n_351),
.Y(n_1085)
);

INVx8_ASAP7_75t_L g1086 ( 
.A(n_953),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_1035),
.B(n_682),
.Y(n_1087)
);

AO32x2_ASAP7_75t_L g1088 ( 
.A1(n_954),
.A2(n_811),
.A3(n_868),
.B1(n_788),
.B2(n_846),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_941),
.A2(n_249),
.B1(n_320),
.B2(n_261),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_928),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_874),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_909),
.Y(n_1092)
);

CKINVDCx16_ASAP7_75t_R g1093 ( 
.A(n_921),
.Y(n_1093)
);

INVxp67_ASAP7_75t_L g1094 ( 
.A(n_894),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1006),
.A2(n_617),
.B(n_644),
.Y(n_1095)
);

AND2x6_ASAP7_75t_L g1096 ( 
.A(n_975),
.B(n_682),
.Y(n_1096)
);

O2A1O1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_912),
.A2(n_634),
.B(n_639),
.C(n_583),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_876),
.B(n_368),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1006),
.A2(n_1029),
.B(n_1001),
.Y(n_1099)
);

INVx1_ASAP7_75t_SL g1100 ( 
.A(n_925),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_989),
.B(n_682),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_941),
.B(n_682),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1006),
.A2(n_644),
.B(n_617),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_959),
.B(n_567),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_897),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_944),
.B(n_446),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_875),
.A2(n_1039),
.B(n_924),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1017),
.A2(n_1020),
.B(n_1009),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_925),
.Y(n_1109)
);

AND2x6_ASAP7_75t_SL g1110 ( 
.A(n_913),
.B(n_446),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_897),
.Y(n_1111)
);

INVx5_ASAP7_75t_L g1112 ( 
.A(n_1003),
.Y(n_1112)
);

AOI21x1_ASAP7_75t_L g1113 ( 
.A1(n_906),
.A2(n_567),
.B(n_568),
.Y(n_1113)
);

AND3x1_ASAP7_75t_SL g1114 ( 
.A(n_974),
.B(n_284),
.C(n_296),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_880),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_891),
.A2(n_644),
.B(n_617),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_908),
.A2(n_644),
.B(n_657),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_942),
.B(n_538),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_905),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_982),
.A2(n_657),
.B(n_637),
.Y(n_1120)
);

OAI221xp5_ASAP7_75t_L g1121 ( 
.A1(n_1012),
.A2(n_348),
.B1(n_300),
.B2(n_302),
.C(n_303),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_905),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_979),
.B(n_372),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_882),
.Y(n_1124)
);

CKINVDCx14_ASAP7_75t_R g1125 ( 
.A(n_1021),
.Y(n_1125)
);

XOR2xp5_ASAP7_75t_L g1126 ( 
.A(n_873),
.B(n_372),
.Y(n_1126)
);

INVxp67_ASAP7_75t_SL g1127 ( 
.A(n_966),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_935),
.A2(n_627),
.B(n_583),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_915),
.Y(n_1129)
);

INVx3_ASAP7_75t_SL g1130 ( 
.A(n_1043),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1028),
.A2(n_627),
.B(n_582),
.Y(n_1131)
);

OAI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_936),
.A2(n_572),
.B(n_568),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_905),
.Y(n_1133)
);

OAI221xp5_ASAP7_75t_L g1134 ( 
.A1(n_952),
.A2(n_309),
.B1(n_312),
.B2(n_383),
.C(n_380),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_916),
.A2(n_380),
.B1(n_383),
.B2(n_385),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_SL g1136 ( 
.A1(n_936),
.A2(n_575),
.B(n_557),
.C(n_545),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_932),
.B(n_927),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_920),
.A2(n_497),
.B1(n_557),
.B2(n_538),
.Y(n_1138)
);

AO32x1_ASAP7_75t_L g1139 ( 
.A1(n_1049),
.A2(n_557),
.A3(n_545),
.B1(n_538),
.B2(n_6),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_927),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_983),
.B(n_545),
.Y(n_1141)
);

XNOR2xp5_ASAP7_75t_L g1142 ( 
.A(n_896),
.B(n_178),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_872),
.B(n_497),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_879),
.B(n_1013),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_886),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_961),
.B(n_1046),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_961),
.B(n_0),
.Y(n_1147)
);

INVx3_ASAP7_75t_SL g1148 ( 
.A(n_913),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_955),
.B(n_1),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_1050),
.B(n_3),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_SL g1151 ( 
.A(n_967),
.B(n_910),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_929),
.B(n_933),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_973),
.A2(n_497),
.B(n_320),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_948),
.A2(n_320),
.B(n_269),
.Y(n_1154)
);

INVx1_ASAP7_75t_SL g1155 ( 
.A(n_980),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1022),
.Y(n_1156)
);

O2A1O1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_952),
.A2(n_971),
.B(n_881),
.C(n_887),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_1004),
.B(n_3),
.Y(n_1158)
);

INVxp67_ASAP7_75t_L g1159 ( 
.A(n_1047),
.Y(n_1159)
);

INVx4_ASAP7_75t_L g1160 ( 
.A(n_964),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_964),
.A2(n_261),
.B(n_258),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1038),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_943),
.B(n_261),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_976),
.A2(n_261),
.B(n_258),
.C(n_249),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_976),
.A2(n_258),
.B(n_249),
.C(n_11),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_955),
.B(n_7),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_1014),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_964),
.A2(n_258),
.B(n_249),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_SL g1169 ( 
.A(n_967),
.B(n_258),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_939),
.A2(n_7),
.B1(n_8),
.B2(n_12),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_964),
.A2(n_497),
.B(n_164),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_970),
.B(n_157),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_922),
.B(n_12),
.Y(n_1173)
);

OAI21xp33_ASAP7_75t_L g1174 ( 
.A1(n_1021),
.A2(n_15),
.B(n_16),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_988),
.A2(n_992),
.B(n_981),
.Y(n_1175)
);

NOR2x1_ASAP7_75t_SL g1176 ( 
.A(n_1003),
.B(n_155),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_1010),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1023),
.B(n_497),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_963),
.A2(n_970),
.B1(n_1047),
.B2(n_1048),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_963),
.B(n_15),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_978),
.A2(n_149),
.B(n_147),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_917),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_1182)
);

A2O1A1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_1048),
.A2(n_18),
.B(n_23),
.C(n_24),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_889),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_986),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_905),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_953),
.B(n_141),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1045),
.B(n_30),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_940),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_923),
.A2(n_136),
.B(n_128),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_958),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1033),
.A2(n_90),
.B(n_85),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_953),
.B(n_34),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_958),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_913),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_949),
.Y(n_1196)
);

AND2x6_ASAP7_75t_L g1197 ( 
.A(n_990),
.B(n_80),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_898),
.Y(n_1198)
);

AOI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1113),
.A2(n_1032),
.B(n_1030),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1144),
.B(n_991),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_1052),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1175),
.A2(n_938),
.B(n_1015),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1115),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1137),
.B(n_1094),
.Y(n_1204)
);

INVxp67_ASAP7_75t_SL g1205 ( 
.A(n_1057),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1107),
.A2(n_902),
.B(n_1025),
.Y(n_1206)
);

INVx3_ASAP7_75t_SL g1207 ( 
.A(n_1092),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1116),
.A2(n_1019),
.B(n_987),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1124),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1051),
.A2(n_1008),
.B(n_962),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1072),
.B(n_1026),
.Y(n_1211)
);

OA21x2_ASAP7_75t_L g1212 ( 
.A1(n_1051),
.A2(n_895),
.B(n_903),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1060),
.B(n_885),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1099),
.A2(n_1003),
.B(n_883),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1054),
.A2(n_939),
.B1(n_937),
.B2(n_934),
.Y(n_1215)
);

NAND2x1_ASAP7_75t_L g1216 ( 
.A(n_1160),
.B(n_877),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1140),
.B(n_1159),
.Y(n_1217)
);

NOR4xp25_ASAP7_75t_L g1218 ( 
.A(n_1174),
.B(n_1000),
.C(n_1016),
.D(n_1041),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1108),
.A2(n_883),
.B(n_947),
.Y(n_1219)
);

NAND3x1_ASAP7_75t_L g1220 ( 
.A(n_1188),
.B(n_931),
.C(n_910),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1056),
.A2(n_937),
.B1(n_934),
.B2(n_1016),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1169),
.A2(n_1071),
.B(n_1064),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_1075),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1169),
.A2(n_997),
.B(n_947),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1062),
.B(n_907),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1145),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1101),
.A2(n_997),
.B(n_995),
.Y(n_1227)
);

AO31x2_ASAP7_75t_L g1228 ( 
.A1(n_1164),
.A2(n_1034),
.A3(n_901),
.B(n_914),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1084),
.B(n_1026),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1068),
.B(n_1026),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1132),
.A2(n_1157),
.B(n_1120),
.Y(n_1231)
);

AOI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1056),
.A2(n_900),
.B1(n_919),
.B2(n_926),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1129),
.B(n_899),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1184),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1090),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1078),
.A2(n_1018),
.B(n_1044),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1155),
.B(n_949),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1131),
.A2(n_1018),
.B(n_1042),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1117),
.A2(n_995),
.B(n_1007),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1155),
.B(n_1179),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_SL g1241 ( 
.A(n_1093),
.B(n_962),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1160),
.A2(n_1007),
.B(n_1037),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1080),
.A2(n_962),
.B(n_999),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_1055),
.B(n_985),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1127),
.A2(n_1037),
.B(n_1027),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1170),
.A2(n_1000),
.B1(n_1037),
.B2(n_977),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1143),
.A2(n_1037),
.B(n_1031),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1146),
.B(n_1058),
.Y(n_1248)
);

AO21x1_ASAP7_75t_L g1249 ( 
.A1(n_1180),
.A2(n_946),
.B(n_1002),
.Y(n_1249)
);

OR2x6_ASAP7_75t_L g1250 ( 
.A(n_1086),
.B(n_960),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1070),
.A2(n_956),
.B(n_994),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1149),
.B(n_969),
.Y(n_1252)
);

NOR3xp33_ASAP7_75t_SL g1253 ( 
.A(n_1085),
.B(n_969),
.C(n_1024),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1141),
.A2(n_951),
.B(n_962),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1141),
.B(n_962),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1102),
.B(n_1198),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1079),
.A2(n_1024),
.B(n_77),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1076),
.A2(n_66),
.B(n_35),
.Y(n_1258)
);

INVx1_ASAP7_75t_SL g1259 ( 
.A(n_1100),
.Y(n_1259)
);

AO31x2_ASAP7_75t_L g1260 ( 
.A1(n_1165),
.A2(n_34),
.A3(n_35),
.B(n_36),
.Y(n_1260)
);

INVx4_ASAP7_75t_L g1261 ( 
.A(n_1112),
.Y(n_1261)
);

OA21x2_ASAP7_75t_L g1262 ( 
.A1(n_1154),
.A2(n_36),
.B(n_40),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1087),
.B(n_41),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1053),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1065),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1083),
.A2(n_42),
.B(n_46),
.Y(n_1266)
);

OA21x2_ASAP7_75t_L g1267 ( 
.A1(n_1153),
.A2(n_42),
.B(n_47),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1177),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1166),
.B(n_49),
.Y(n_1269)
);

AO21x2_ASAP7_75t_L g1270 ( 
.A1(n_1136),
.A2(n_50),
.B(n_52),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1153),
.A2(n_54),
.B(n_55),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1066),
.Y(n_1272)
);

AOI221x1_ASAP7_75t_L g1273 ( 
.A1(n_1063),
.A2(n_1170),
.B1(n_1183),
.B2(n_1192),
.C(n_1173),
.Y(n_1273)
);

AOI221xp5_ASAP7_75t_SL g1274 ( 
.A1(n_1063),
.A2(n_1069),
.B1(n_1185),
.B2(n_1182),
.C(n_1067),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1100),
.B(n_56),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1077),
.A2(n_58),
.B(n_59),
.Y(n_1276)
);

NOR4xp25_ASAP7_75t_L g1277 ( 
.A(n_1134),
.B(n_59),
.C(n_62),
.D(n_64),
.Y(n_1277)
);

O2A1O1Ixp5_ASAP7_75t_SL g1278 ( 
.A1(n_1192),
.A2(n_64),
.B(n_1163),
.C(n_1123),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1172),
.B(n_1187),
.Y(n_1279)
);

INVx3_ASAP7_75t_SL g1280 ( 
.A(n_1130),
.Y(n_1280)
);

INVx5_ASAP7_75t_L g1281 ( 
.A(n_1112),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1095),
.A2(n_1103),
.B(n_1097),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1074),
.B(n_1118),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1189),
.Y(n_1284)
);

AOI211x1_ASAP7_75t_L g1285 ( 
.A1(n_1121),
.A2(n_1152),
.B(n_1193),
.C(n_1135),
.Y(n_1285)
);

O2A1O1Ixp5_ASAP7_75t_L g1286 ( 
.A1(n_1081),
.A2(n_1190),
.B(n_1181),
.C(n_1135),
.Y(n_1286)
);

NAND2xp33_ASAP7_75t_SL g1287 ( 
.A(n_1061),
.B(n_1148),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1151),
.A2(n_1104),
.B(n_1178),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1118),
.B(n_1187),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1191),
.A2(n_1194),
.B(n_1161),
.Y(n_1290)
);

INVxp67_ASAP7_75t_SL g1291 ( 
.A(n_1052),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1191),
.A2(n_1194),
.B(n_1168),
.Y(n_1292)
);

O2A1O1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1150),
.A2(n_1158),
.B(n_1098),
.C(n_1147),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1156),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1172),
.B(n_1082),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1151),
.B(n_1196),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1162),
.Y(n_1297)
);

INVx1_ASAP7_75t_SL g1298 ( 
.A(n_1106),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1059),
.A2(n_1186),
.B(n_1133),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_1109),
.Y(n_1300)
);

A2O1A1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1089),
.A2(n_1073),
.B(n_1086),
.C(n_1138),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1171),
.A2(n_1096),
.B(n_1197),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1059),
.B(n_1186),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_SL g1304 ( 
.A1(n_1176),
.A2(n_1052),
.B(n_1122),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_SL g1305 ( 
.A1(n_1105),
.A2(n_1122),
.B(n_1119),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1086),
.A2(n_1142),
.B1(n_1112),
.B2(n_1105),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1139),
.A2(n_1133),
.B(n_1105),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1195),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1088),
.A2(n_1096),
.B(n_1139),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1125),
.B(n_1126),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1096),
.B(n_1119),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_1110),
.Y(n_1312)
);

NAND3xp33_ASAP7_75t_SL g1313 ( 
.A(n_1114),
.B(n_1197),
.C(n_1167),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1111),
.B(n_1119),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1111),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1111),
.A2(n_1122),
.B1(n_1139),
.B2(n_1096),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_SL g1317 ( 
.A1(n_1197),
.A2(n_1040),
.B(n_1005),
.Y(n_1317)
);

O2A1O1Ixp33_ASAP7_75t_SL g1318 ( 
.A1(n_1197),
.A2(n_1005),
.B(n_1054),
.C(n_1165),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1088),
.B(n_1144),
.Y(n_1319)
);

AO31x2_ASAP7_75t_L g1320 ( 
.A1(n_1088),
.A2(n_1107),
.A3(n_1164),
.B(n_1175),
.Y(n_1320)
);

NOR2xp67_ASAP7_75t_L g1321 ( 
.A(n_1092),
.B(n_571),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1144),
.B(n_984),
.Y(n_1322)
);

AOI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1060),
.A2(n_884),
.B1(n_668),
.B2(n_729),
.Y(n_1323)
);

INVx2_ASAP7_75t_SL g1324 ( 
.A(n_1090),
.Y(n_1324)
);

OAI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1107),
.A2(n_904),
.B(n_1051),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1113),
.A2(n_1116),
.B(n_1128),
.Y(n_1326)
);

INVx5_ASAP7_75t_L g1327 ( 
.A(n_1160),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1060),
.B(n_387),
.Y(n_1328)
);

AO21x2_ASAP7_75t_L g1329 ( 
.A1(n_1107),
.A2(n_1099),
.B(n_1136),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1107),
.A2(n_904),
.B(n_1051),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1094),
.B(n_571),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1144),
.B(n_984),
.Y(n_1332)
);

NAND2x1p5_ASAP7_75t_L g1333 ( 
.A(n_1112),
.B(n_1160),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1175),
.A2(n_1040),
.B(n_993),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1091),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1090),
.Y(n_1336)
);

AO31x2_ASAP7_75t_L g1337 ( 
.A1(n_1107),
.A2(n_1164),
.A3(n_1175),
.B(n_1099),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1057),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1113),
.A2(n_1116),
.B(n_1128),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1057),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1175),
.A2(n_1040),
.B(n_993),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1175),
.A2(n_1040),
.B(n_993),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1113),
.A2(n_1116),
.B(n_1128),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1113),
.A2(n_1116),
.B(n_1128),
.Y(n_1344)
);

NAND2xp33_ASAP7_75t_R g1345 ( 
.A(n_1092),
.B(n_570),
.Y(n_1345)
);

AO31x2_ASAP7_75t_L g1346 ( 
.A1(n_1107),
.A2(n_1164),
.A3(n_1175),
.B(n_1099),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1175),
.A2(n_1040),
.B(n_993),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1144),
.B(n_984),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1052),
.Y(n_1349)
);

NOR2xp67_ASAP7_75t_L g1350 ( 
.A(n_1092),
.B(n_571),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_1092),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1091),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1054),
.A2(n_984),
.B(n_729),
.C(n_1005),
.Y(n_1353)
);

INVx2_ASAP7_75t_SL g1354 ( 
.A(n_1090),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1208),
.A2(n_1339),
.B(n_1326),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1343),
.A2(n_1344),
.B(n_1254),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1348),
.B(n_1322),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1203),
.Y(n_1358)
);

AO21x2_ASAP7_75t_L g1359 ( 
.A1(n_1231),
.A2(n_1330),
.B(n_1325),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1209),
.Y(n_1360)
);

OR2x6_ASAP7_75t_L g1361 ( 
.A(n_1279),
.B(n_1317),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1322),
.B(n_1332),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1214),
.A2(n_1341),
.B(n_1334),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1342),
.A2(n_1347),
.B(n_1282),
.Y(n_1364)
);

AOI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1199),
.A2(n_1222),
.B(n_1225),
.Y(n_1365)
);

OA21x2_ASAP7_75t_L g1366 ( 
.A1(n_1231),
.A2(n_1309),
.B(n_1325),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1204),
.B(n_1252),
.Y(n_1367)
);

BUFx2_ASAP7_75t_SL g1368 ( 
.A(n_1235),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1226),
.Y(n_1369)
);

A2O1A1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1276),
.A2(n_1271),
.B(n_1353),
.C(n_1323),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1219),
.A2(n_1239),
.B(n_1202),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1234),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1251),
.A2(n_1247),
.B(n_1236),
.Y(n_1373)
);

OAI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1273),
.A2(n_1274),
.B(n_1293),
.Y(n_1374)
);

OAI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1274),
.A2(n_1276),
.B(n_1225),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1332),
.A2(n_1328),
.B1(n_1213),
.B2(n_1200),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1335),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1352),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1200),
.A2(n_1289),
.B1(n_1240),
.B2(n_1230),
.Y(n_1379)
);

O2A1O1Ixp5_ASAP7_75t_L g1380 ( 
.A1(n_1271),
.A2(n_1257),
.B(n_1286),
.C(n_1243),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1269),
.B(n_1237),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1206),
.A2(n_1302),
.B(n_1290),
.Y(n_1382)
);

INVx8_ASAP7_75t_L g1383 ( 
.A(n_1281),
.Y(n_1383)
);

AOI221xp5_ASAP7_75t_L g1384 ( 
.A1(n_1277),
.A2(n_1318),
.B1(n_1221),
.B2(n_1285),
.C(n_1218),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1264),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1265),
.Y(n_1386)
);

OAI211xp5_ASAP7_75t_L g1387 ( 
.A1(n_1263),
.A2(n_1275),
.B(n_1232),
.C(n_1248),
.Y(n_1387)
);

INVxp67_ASAP7_75t_L g1388 ( 
.A(n_1338),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1278),
.A2(n_1288),
.B(n_1229),
.Y(n_1389)
);

NAND2x1p5_ASAP7_75t_L g1390 ( 
.A(n_1281),
.B(n_1327),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_SL g1391 ( 
.A1(n_1256),
.A2(n_1307),
.B(n_1302),
.Y(n_1391)
);

BUFx10_ASAP7_75t_L g1392 ( 
.A(n_1351),
.Y(n_1392)
);

CKINVDCx8_ASAP7_75t_R g1393 ( 
.A(n_1223),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1272),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1250),
.B(n_1314),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1238),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1211),
.B(n_1298),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1284),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1206),
.A2(n_1292),
.B(n_1227),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1340),
.B(n_1298),
.Y(n_1400)
);

CKINVDCx14_ASAP7_75t_R g1401 ( 
.A(n_1287),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1221),
.A2(n_1241),
.B1(n_1306),
.B2(n_1312),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1297),
.Y(n_1403)
);

INVx1_ASAP7_75t_SL g1404 ( 
.A(n_1259),
.Y(n_1404)
);

OA21x2_ASAP7_75t_L g1405 ( 
.A1(n_1210),
.A2(n_1243),
.B(n_1319),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1245),
.A2(n_1266),
.B(n_1242),
.Y(n_1406)
);

CKINVDCx6p67_ASAP7_75t_R g1407 ( 
.A(n_1280),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1215),
.A2(n_1267),
.B1(n_1313),
.B2(n_1295),
.Y(n_1408)
);

O2A1O1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1296),
.A2(n_1301),
.B(n_1306),
.C(n_1253),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1255),
.A2(n_1224),
.B(n_1316),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1256),
.B(n_1331),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1250),
.B(n_1294),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1215),
.A2(n_1267),
.B1(n_1270),
.B2(n_1308),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1255),
.A2(n_1316),
.B(n_1258),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1283),
.B(n_1217),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1299),
.A2(n_1246),
.B(n_1212),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1246),
.A2(n_1212),
.B(n_1319),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1311),
.A2(n_1262),
.B(n_1216),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_1281),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1345),
.A2(n_1321),
.B1(n_1350),
.B2(n_1241),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1228),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1244),
.A2(n_1233),
.B(n_1217),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1311),
.A2(n_1262),
.B(n_1304),
.Y(n_1423)
);

BUFx12f_ASAP7_75t_L g1424 ( 
.A(n_1324),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1228),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1233),
.A2(n_1303),
.B(n_1291),
.Y(n_1426)
);

BUFx6f_ASAP7_75t_L g1427 ( 
.A(n_1281),
.Y(n_1427)
);

OA21x2_ASAP7_75t_L g1428 ( 
.A1(n_1303),
.A2(n_1320),
.B(n_1329),
.Y(n_1428)
);

AO21x2_ASAP7_75t_L g1429 ( 
.A1(n_1329),
.A2(n_1270),
.B(n_1346),
.Y(n_1429)
);

AO21x2_ASAP7_75t_L g1430 ( 
.A1(n_1337),
.A2(n_1346),
.B(n_1228),
.Y(n_1430)
);

O2A1O1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1250),
.A2(n_1268),
.B(n_1310),
.C(n_1354),
.Y(n_1431)
);

A2O1A1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1260),
.A2(n_1327),
.B(n_1320),
.C(n_1315),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1320),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1336),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1333),
.A2(n_1305),
.B(n_1346),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1337),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1207),
.B(n_1300),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_1261),
.B(n_1201),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1201),
.B(n_1349),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1349),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1220),
.A2(n_1323),
.B1(n_1348),
.B2(n_984),
.Y(n_1441)
);

AND2x6_ASAP7_75t_L g1442 ( 
.A(n_1232),
.B(n_1187),
.Y(n_1442)
);

NAND2x1p5_ASAP7_75t_L g1443 ( 
.A(n_1281),
.B(n_1327),
.Y(n_1443)
);

OA21x2_ASAP7_75t_L g1444 ( 
.A1(n_1231),
.A2(n_1309),
.B(n_1325),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1208),
.A2(n_1339),
.B(n_1326),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1208),
.A2(n_1339),
.B(n_1326),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1348),
.B(n_1322),
.Y(n_1447)
);

OAI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1323),
.A2(n_729),
.B(n_984),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_SL g1449 ( 
.A(n_1351),
.B(n_733),
.Y(n_1449)
);

CKINVDCx16_ASAP7_75t_R g1450 ( 
.A(n_1345),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1204),
.B(n_1137),
.Y(n_1451)
);

NOR2xp67_ASAP7_75t_L g1452 ( 
.A(n_1351),
.B(n_571),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1208),
.A2(n_1339),
.B(n_1326),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1204),
.B(n_1137),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_SL g1455 ( 
.A1(n_1276),
.A2(n_1271),
.B(n_1256),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1208),
.A2(n_1339),
.B(n_1326),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1208),
.A2(n_1339),
.B(n_1326),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1345),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1205),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1208),
.A2(n_1339),
.B(n_1326),
.Y(n_1460)
);

OA21x2_ASAP7_75t_L g1461 ( 
.A1(n_1231),
.A2(n_1309),
.B(n_1325),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_1351),
.Y(n_1462)
);

AO31x2_ASAP7_75t_L g1463 ( 
.A1(n_1249),
.A2(n_1273),
.A3(n_1316),
.B(n_1319),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1348),
.B(n_1322),
.Y(n_1464)
);

OAI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1323),
.A2(n_729),
.B(n_984),
.Y(n_1465)
);

AO21x2_ASAP7_75t_L g1466 ( 
.A1(n_1231),
.A2(n_1330),
.B(n_1325),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1205),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1348),
.B(n_1322),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1203),
.Y(n_1469)
);

AO21x2_ASAP7_75t_L g1470 ( 
.A1(n_1231),
.A2(n_1330),
.B(n_1325),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1276),
.A2(n_984),
.B1(n_1323),
.B2(n_1036),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1208),
.A2(n_1339),
.B(n_1326),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1208),
.A2(n_1339),
.B(n_1326),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1203),
.Y(n_1474)
);

AO31x2_ASAP7_75t_L g1475 ( 
.A1(n_1249),
.A2(n_1273),
.A3(n_1316),
.B(n_1319),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1208),
.A2(n_1339),
.B(n_1326),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1208),
.A2(n_1339),
.B(n_1326),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1203),
.Y(n_1478)
);

INVxp67_ASAP7_75t_L g1479 ( 
.A(n_1338),
.Y(n_1479)
);

INVx3_ASAP7_75t_L g1480 ( 
.A(n_1281),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_SL g1481 ( 
.A1(n_1276),
.A2(n_1271),
.B(n_1256),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1204),
.B(n_1137),
.Y(n_1482)
);

AO21x2_ASAP7_75t_L g1483 ( 
.A1(n_1231),
.A2(n_1330),
.B(n_1325),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1203),
.Y(n_1484)
);

OR2x6_ASAP7_75t_L g1485 ( 
.A(n_1279),
.B(n_1317),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1323),
.A2(n_1348),
.B1(n_984),
.B2(n_1332),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1203),
.Y(n_1487)
);

INVx2_ASAP7_75t_SL g1488 ( 
.A(n_1235),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1203),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_SL g1490 ( 
.A1(n_1276),
.A2(n_1271),
.B(n_1256),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1250),
.B(n_1279),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1276),
.A2(n_984),
.B1(n_1323),
.B2(n_1036),
.Y(n_1492)
);

BUFx12f_ASAP7_75t_L g1493 ( 
.A(n_1351),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1203),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1348),
.B(n_1322),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1235),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1203),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1205),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1208),
.A2(n_1339),
.B(n_1326),
.Y(n_1499)
);

O2A1O1Ixp5_ASAP7_75t_L g1500 ( 
.A1(n_1448),
.A2(n_1465),
.B(n_1380),
.C(n_1370),
.Y(n_1500)
);

NOR2xp67_ASAP7_75t_L g1501 ( 
.A(n_1420),
.B(n_1452),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1376),
.B(n_1362),
.Y(n_1502)
);

O2A1O1Ixp33_ASAP7_75t_L g1503 ( 
.A1(n_1370),
.A2(n_1441),
.B(n_1492),
.C(n_1471),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1357),
.B(n_1447),
.Y(n_1504)
);

OA21x2_ASAP7_75t_L g1505 ( 
.A1(n_1371),
.A2(n_1417),
.B(n_1389),
.Y(n_1505)
);

CKINVDCx6p67_ASAP7_75t_R g1506 ( 
.A(n_1462),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1451),
.B(n_1454),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1482),
.B(n_1381),
.Y(n_1508)
);

AOI21x1_ASAP7_75t_SL g1509 ( 
.A1(n_1425),
.A2(n_1491),
.B(n_1468),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1367),
.B(n_1415),
.Y(n_1510)
);

AOI21xp5_ASAP7_75t_SL g1511 ( 
.A1(n_1458),
.A2(n_1486),
.B(n_1409),
.Y(n_1511)
);

O2A1O1Ixp5_ASAP7_75t_L g1512 ( 
.A1(n_1375),
.A2(n_1374),
.B(n_1387),
.C(n_1365),
.Y(n_1512)
);

AOI21xp5_ASAP7_75t_SL g1513 ( 
.A1(n_1458),
.A2(n_1443),
.B(n_1390),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1415),
.B(n_1422),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1471),
.A2(n_1492),
.B1(n_1402),
.B2(n_1401),
.Y(n_1515)
);

OA21x2_ASAP7_75t_L g1516 ( 
.A1(n_1371),
.A2(n_1417),
.B(n_1355),
.Y(n_1516)
);

INVx2_ASAP7_75t_SL g1517 ( 
.A(n_1496),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1397),
.B(n_1411),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1442),
.A2(n_1450),
.B1(n_1491),
.B2(n_1449),
.Y(n_1519)
);

AOI211xp5_ASAP7_75t_L g1520 ( 
.A1(n_1431),
.A2(n_1384),
.B(n_1379),
.C(n_1495),
.Y(n_1520)
);

O2A1O1Ixp33_ASAP7_75t_L g1521 ( 
.A1(n_1455),
.A2(n_1490),
.B(n_1481),
.C(n_1464),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_SL g1522 ( 
.A1(n_1390),
.A2(n_1443),
.B(n_1427),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1395),
.B(n_1404),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1369),
.Y(n_1524)
);

A2O1A1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1408),
.A2(n_1413),
.B(n_1442),
.C(n_1432),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1395),
.B(n_1400),
.Y(n_1526)
);

AOI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1442),
.A2(n_1401),
.B1(n_1437),
.B2(n_1395),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1359),
.A2(n_1466),
.B(n_1483),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1359),
.A2(n_1466),
.B(n_1483),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1360),
.B(n_1489),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1360),
.B(n_1489),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1426),
.B(n_1358),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_SL g1533 ( 
.A1(n_1419),
.A2(n_1427),
.B(n_1361),
.Y(n_1533)
);

AOI21xp5_ASAP7_75t_SL g1534 ( 
.A1(n_1419),
.A2(n_1427),
.B(n_1361),
.Y(n_1534)
);

O2A1O1Ixp33_ASAP7_75t_L g1535 ( 
.A1(n_1388),
.A2(n_1479),
.B(n_1459),
.C(n_1498),
.Y(n_1535)
);

O2A1O1Ixp5_ASAP7_75t_L g1536 ( 
.A1(n_1436),
.A2(n_1421),
.B(n_1432),
.C(n_1433),
.Y(n_1536)
);

OA21x2_ASAP7_75t_L g1537 ( 
.A1(n_1355),
.A2(n_1460),
.B(n_1477),
.Y(n_1537)
);

NOR2x1_ASAP7_75t_SL g1538 ( 
.A(n_1361),
.B(n_1485),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1470),
.A2(n_1363),
.B(n_1485),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1469),
.B(n_1474),
.Y(n_1540)
);

OA22x2_ASAP7_75t_L g1541 ( 
.A1(n_1412),
.A2(n_1467),
.B1(n_1498),
.B2(n_1386),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1372),
.B(n_1377),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1378),
.Y(n_1543)
);

OA21x2_ASAP7_75t_L g1544 ( 
.A1(n_1445),
.A2(n_1499),
.B(n_1477),
.Y(n_1544)
);

O2A1O1Ixp5_ASAP7_75t_L g1545 ( 
.A1(n_1436),
.A2(n_1433),
.B(n_1396),
.C(n_1394),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1478),
.B(n_1484),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1487),
.B(n_1494),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1497),
.B(n_1398),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1408),
.A2(n_1437),
.B1(n_1413),
.B2(n_1434),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1496),
.A2(n_1385),
.B1(n_1368),
.B2(n_1488),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1403),
.B(n_1405),
.Y(n_1551)
);

INVx1_ASAP7_75t_SL g1552 ( 
.A(n_1462),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1440),
.B(n_1439),
.Y(n_1553)
);

OA21x2_ASAP7_75t_L g1554 ( 
.A1(n_1445),
.A2(n_1499),
.B(n_1476),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1438),
.B(n_1442),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1405),
.B(n_1463),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1405),
.B(n_1463),
.Y(n_1557)
);

A2O1A1Ixp33_ASAP7_75t_L g1558 ( 
.A1(n_1414),
.A2(n_1435),
.B(n_1410),
.C(n_1382),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1438),
.B(n_1393),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1392),
.B(n_1480),
.Y(n_1560)
);

O2A1O1Ixp5_ASAP7_75t_L g1561 ( 
.A1(n_1391),
.A2(n_1429),
.B(n_1430),
.C(n_1463),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1428),
.Y(n_1562)
);

NAND2xp33_ASAP7_75t_SL g1563 ( 
.A(n_1383),
.B(n_1430),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1392),
.B(n_1475),
.Y(n_1564)
);

AOI21x1_ASAP7_75t_SL g1565 ( 
.A1(n_1383),
.A2(n_1423),
.B(n_1463),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1475),
.B(n_1461),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1475),
.B(n_1461),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1475),
.B(n_1444),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1364),
.A2(n_1399),
.B(n_1435),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1366),
.B(n_1444),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1423),
.B(n_1418),
.Y(n_1571)
);

OAI211xp5_ASAP7_75t_L g1572 ( 
.A1(n_1366),
.A2(n_1382),
.B(n_1418),
.C(n_1416),
.Y(n_1572)
);

O2A1O1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1424),
.A2(n_1407),
.B(n_1406),
.C(n_1493),
.Y(n_1573)
);

OA21x2_ASAP7_75t_L g1574 ( 
.A1(n_1446),
.A2(n_1456),
.B(n_1476),
.Y(n_1574)
);

CKINVDCx20_ASAP7_75t_R g1575 ( 
.A(n_1493),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1424),
.Y(n_1576)
);

OA21x2_ASAP7_75t_L g1577 ( 
.A1(n_1446),
.A2(n_1457),
.B(n_1472),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1373),
.B(n_1356),
.Y(n_1578)
);

CKINVDCx8_ASAP7_75t_R g1579 ( 
.A(n_1453),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1453),
.B(n_1456),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1457),
.B(n_1473),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1473),
.B(n_1460),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1472),
.B(n_1451),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1471),
.A2(n_1323),
.B1(n_1492),
.B2(n_1035),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1376),
.B(n_1362),
.Y(n_1585)
);

O2A1O1Ixp33_ASAP7_75t_L g1586 ( 
.A1(n_1448),
.A2(n_1465),
.B(n_1353),
.C(n_1370),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1451),
.B(n_1454),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1448),
.A2(n_1465),
.B(n_1005),
.Y(n_1588)
);

INVx4_ASAP7_75t_SL g1589 ( 
.A(n_1442),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1471),
.A2(n_1323),
.B1(n_1492),
.B2(n_1035),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1451),
.B(n_1454),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1491),
.B(n_1395),
.Y(n_1592)
);

AOI221x1_ASAP7_75t_SL g1593 ( 
.A1(n_1441),
.A2(n_805),
.B1(n_675),
.B2(n_1188),
.C(n_509),
.Y(n_1593)
);

O2A1O1Ixp5_ASAP7_75t_L g1594 ( 
.A1(n_1448),
.A2(n_1465),
.B(n_1380),
.C(n_1370),
.Y(n_1594)
);

O2A1O1Ixp5_ASAP7_75t_L g1595 ( 
.A1(n_1448),
.A2(n_1465),
.B(n_1380),
.C(n_1370),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_SL g1596 ( 
.A1(n_1450),
.A2(n_1323),
.B1(n_1458),
.B2(n_1471),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1376),
.B(n_1362),
.Y(n_1597)
);

OA21x2_ASAP7_75t_L g1598 ( 
.A1(n_1380),
.A2(n_1371),
.B(n_1417),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1400),
.B(n_1459),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1451),
.B(n_1454),
.Y(n_1600)
);

INVx1_ASAP7_75t_SL g1601 ( 
.A(n_1404),
.Y(n_1601)
);

AND2x6_ASAP7_75t_L g1602 ( 
.A(n_1491),
.B(n_1419),
.Y(n_1602)
);

AOI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1471),
.A2(n_1323),
.B1(n_668),
.B2(n_1035),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1451),
.B(n_1454),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1451),
.B(n_1454),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1471),
.A2(n_1323),
.B1(n_1492),
.B2(n_1035),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1451),
.B(n_1454),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_SL g1608 ( 
.A(n_1449),
.B(n_733),
.Y(n_1608)
);

O2A1O1Ixp33_ASAP7_75t_L g1609 ( 
.A1(n_1448),
.A2(n_1465),
.B(n_1353),
.C(n_1370),
.Y(n_1609)
);

INVx3_ASAP7_75t_SL g1610 ( 
.A(n_1458),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1451),
.B(n_1454),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1376),
.B(n_1362),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1451),
.B(n_1454),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1551),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1570),
.B(n_1583),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1584),
.A2(n_1606),
.B1(n_1590),
.B2(n_1603),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1506),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1567),
.B(n_1568),
.Y(n_1618)
);

INVx4_ASAP7_75t_L g1619 ( 
.A(n_1589),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1502),
.B(n_1585),
.Y(n_1620)
);

INVx2_ASAP7_75t_SL g1621 ( 
.A(n_1541),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1556),
.B(n_1557),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1571),
.B(n_1589),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1596),
.A2(n_1515),
.B1(n_1588),
.B2(n_1597),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1571),
.Y(n_1625)
);

OAI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1500),
.A2(n_1595),
.B(n_1594),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1566),
.B(n_1528),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1529),
.B(n_1564),
.Y(n_1628)
);

AOI211xp5_ASAP7_75t_L g1629 ( 
.A1(n_1503),
.A2(n_1511),
.B(n_1586),
.C(n_1609),
.Y(n_1629)
);

AO21x2_ASAP7_75t_L g1630 ( 
.A1(n_1569),
.A2(n_1525),
.B(n_1572),
.Y(n_1630)
);

INVx3_ASAP7_75t_L g1631 ( 
.A(n_1579),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1505),
.B(n_1598),
.Y(n_1632)
);

AOI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1593),
.A2(n_1500),
.B1(n_1595),
.B2(n_1594),
.C(n_1612),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1562),
.B(n_1598),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1545),
.Y(n_1635)
);

AO21x2_ASAP7_75t_L g1636 ( 
.A1(n_1525),
.A2(n_1558),
.B(n_1539),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1536),
.Y(n_1637)
);

OA21x2_ASAP7_75t_L g1638 ( 
.A1(n_1561),
.A2(n_1512),
.B(n_1558),
.Y(n_1638)
);

NOR2x1_ASAP7_75t_SL g1639 ( 
.A(n_1549),
.B(n_1555),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1524),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1541),
.B(n_1516),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1518),
.B(n_1599),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1516),
.Y(n_1643)
);

BUFx3_ASAP7_75t_L g1644 ( 
.A(n_1602),
.Y(n_1644)
);

BUFx12f_ASAP7_75t_L g1645 ( 
.A(n_1576),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1520),
.B(n_1532),
.Y(n_1646)
);

AO21x2_ASAP7_75t_L g1647 ( 
.A1(n_1578),
.A2(n_1581),
.B(n_1582),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1543),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1589),
.B(n_1538),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1580),
.B(n_1592),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1542),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1516),
.B(n_1514),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1537),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_SL g1654 ( 
.A(n_1512),
.B(n_1521),
.Y(n_1654)
);

AO22x1_ASAP7_75t_L g1655 ( 
.A1(n_1602),
.A2(n_1610),
.B1(n_1560),
.B2(n_1550),
.Y(n_1655)
);

OR2x6_ASAP7_75t_L g1656 ( 
.A(n_1513),
.B(n_1534),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1530),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1544),
.B(n_1574),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1544),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1510),
.B(n_1531),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1548),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1546),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1554),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1554),
.B(n_1574),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1504),
.B(n_1535),
.Y(n_1665)
);

OA21x2_ASAP7_75t_L g1666 ( 
.A1(n_1547),
.A2(n_1519),
.B(n_1527),
.Y(n_1666)
);

INVxp67_ASAP7_75t_L g1667 ( 
.A(n_1614),
.Y(n_1667)
);

INVx4_ASAP7_75t_L g1668 ( 
.A(n_1619),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1640),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1627),
.B(n_1577),
.Y(n_1670)
);

AOI221xp5_ASAP7_75t_L g1671 ( 
.A1(n_1633),
.A2(n_1601),
.B1(n_1508),
.B2(n_1507),
.C(n_1611),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1620),
.B(n_1614),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1640),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1620),
.B(n_1540),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1615),
.B(n_1526),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1615),
.B(n_1592),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1648),
.Y(n_1677)
);

CKINVDCx20_ASAP7_75t_R g1678 ( 
.A(n_1617),
.Y(n_1678)
);

AOI211xp5_ASAP7_75t_L g1679 ( 
.A1(n_1629),
.A2(n_1501),
.B(n_1573),
.C(n_1608),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1615),
.B(n_1523),
.Y(n_1680)
);

OA21x2_ASAP7_75t_L g1681 ( 
.A1(n_1626),
.A2(n_1565),
.B(n_1509),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1616),
.A2(n_1624),
.B1(n_1633),
.B2(n_1646),
.Y(n_1682)
);

NAND2x1p5_ASAP7_75t_L g1683 ( 
.A(n_1654),
.B(n_1509),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1627),
.B(n_1652),
.Y(n_1684)
);

OAI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1646),
.A2(n_1610),
.B1(n_1575),
.B2(n_1559),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1652),
.B(n_1587),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1623),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1652),
.B(n_1563),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1647),
.B(n_1613),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1647),
.B(n_1604),
.Y(n_1690)
);

BUFx3_ASAP7_75t_L g1691 ( 
.A(n_1631),
.Y(n_1691)
);

NAND2x1_ASAP7_75t_L g1692 ( 
.A(n_1619),
.B(n_1533),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1616),
.A2(n_1600),
.B1(n_1591),
.B2(n_1607),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1625),
.B(n_1602),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1647),
.B(n_1605),
.Y(n_1695)
);

BUFx3_ASAP7_75t_L g1696 ( 
.A(n_1631),
.Y(n_1696)
);

OAI21xp5_ASAP7_75t_SL g1697 ( 
.A1(n_1624),
.A2(n_1552),
.B(n_1517),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1653),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1647),
.B(n_1553),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1679),
.A2(n_1654),
.B(n_1629),
.Y(n_1700)
);

AOI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1679),
.A2(n_1656),
.B(n_1639),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1698),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_1672),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_1678),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1669),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1698),
.Y(n_1706)
);

OAI21xp33_ASAP7_75t_SL g1707 ( 
.A1(n_1672),
.A2(n_1656),
.B(n_1621),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1669),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1686),
.B(n_1676),
.Y(n_1709)
);

AOI222xp33_ASAP7_75t_L g1710 ( 
.A1(n_1682),
.A2(n_1639),
.B1(n_1665),
.B2(n_1621),
.C1(n_1642),
.C2(n_1637),
.Y(n_1710)
);

OAI221xp5_ASAP7_75t_L g1711 ( 
.A1(n_1682),
.A2(n_1665),
.B1(n_1621),
.B2(n_1656),
.C(n_1642),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_L g1712 ( 
.A(n_1685),
.B(n_1674),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1673),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1673),
.Y(n_1714)
);

OAI221xp5_ASAP7_75t_L g1715 ( 
.A1(n_1697),
.A2(n_1656),
.B1(n_1631),
.B2(n_1662),
.C(n_1666),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1677),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1671),
.A2(n_1666),
.B1(n_1636),
.B2(n_1656),
.Y(n_1717)
);

INVx3_ASAP7_75t_L g1718 ( 
.A(n_1687),
.Y(n_1718)
);

BUFx10_ASAP7_75t_L g1719 ( 
.A(n_1694),
.Y(n_1719)
);

AOI211xp5_ASAP7_75t_L g1720 ( 
.A1(n_1685),
.A2(n_1655),
.B(n_1662),
.C(n_1628),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1671),
.A2(n_1666),
.B1(n_1636),
.B2(n_1656),
.Y(n_1721)
);

BUFx10_ASAP7_75t_L g1722 ( 
.A(n_1694),
.Y(n_1722)
);

INVx3_ASAP7_75t_L g1723 ( 
.A(n_1687),
.Y(n_1723)
);

OAI21x1_ASAP7_75t_L g1724 ( 
.A1(n_1683),
.A2(n_1635),
.B(n_1643),
.Y(n_1724)
);

AND2x4_ASAP7_75t_SL g1725 ( 
.A(n_1668),
.B(n_1619),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1684),
.B(n_1622),
.Y(n_1726)
);

NAND4xp25_ASAP7_75t_L g1727 ( 
.A(n_1693),
.B(n_1628),
.C(n_1651),
.D(n_1641),
.Y(n_1727)
);

NAND4xp25_ASAP7_75t_SL g1728 ( 
.A(n_1693),
.B(n_1575),
.C(n_1678),
.D(n_1674),
.Y(n_1728)
);

AOI221xp5_ASAP7_75t_L g1729 ( 
.A1(n_1697),
.A2(n_1651),
.B1(n_1661),
.B2(n_1628),
.C(n_1641),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1680),
.Y(n_1730)
);

AOI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1692),
.A2(n_1666),
.B1(n_1649),
.B2(n_1619),
.Y(n_1731)
);

NAND2xp33_ASAP7_75t_R g1732 ( 
.A(n_1681),
.B(n_1631),
.Y(n_1732)
);

AOI221xp5_ASAP7_75t_L g1733 ( 
.A1(n_1689),
.A2(n_1661),
.B1(n_1641),
.B2(n_1657),
.C(n_1660),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1686),
.B(n_1650),
.Y(n_1734)
);

OAI21xp33_ASAP7_75t_L g1735 ( 
.A1(n_1683),
.A2(n_1622),
.B(n_1618),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_R g1736 ( 
.A(n_1668),
.B(n_1645),
.Y(n_1736)
);

INVxp67_ASAP7_75t_L g1737 ( 
.A(n_1680),
.Y(n_1737)
);

AOI221xp5_ASAP7_75t_L g1738 ( 
.A1(n_1689),
.A2(n_1657),
.B1(n_1660),
.B2(n_1636),
.C(n_1622),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_SL g1739 ( 
.A(n_1683),
.B(n_1649),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1686),
.B(n_1650),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1683),
.B(n_1676),
.Y(n_1741)
);

OAI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1692),
.A2(n_1619),
.B1(n_1644),
.B2(n_1631),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1681),
.A2(n_1636),
.B1(n_1630),
.B2(n_1645),
.Y(n_1743)
);

OAI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1692),
.A2(n_1691),
.B1(n_1696),
.B2(n_1688),
.C(n_1667),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1705),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1708),
.Y(n_1746)
);

INVxp67_ASAP7_75t_SL g1747 ( 
.A(n_1732),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1709),
.B(n_1689),
.Y(n_1748)
);

INVx4_ASAP7_75t_L g1749 ( 
.A(n_1725),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1724),
.Y(n_1750)
);

INVxp67_ASAP7_75t_L g1751 ( 
.A(n_1732),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1713),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1702),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1734),
.B(n_1690),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1700),
.B(n_1675),
.Y(n_1755)
);

INVxp67_ASAP7_75t_SL g1756 ( 
.A(n_1706),
.Y(n_1756)
);

INVxp67_ASAP7_75t_SL g1757 ( 
.A(n_1706),
.Y(n_1757)
);

NOR3xp33_ASAP7_75t_L g1758 ( 
.A(n_1728),
.B(n_1655),
.C(n_1668),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1714),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1716),
.Y(n_1760)
);

INVx2_ASAP7_75t_SL g1761 ( 
.A(n_1719),
.Y(n_1761)
);

AND4x1_ASAP7_75t_L g1762 ( 
.A(n_1720),
.B(n_1522),
.C(n_1645),
.D(n_1695),
.Y(n_1762)
);

AOI21x1_ASAP7_75t_L g1763 ( 
.A1(n_1739),
.A2(n_1663),
.B(n_1664),
.Y(n_1763)
);

INVxp67_ASAP7_75t_SL g1764 ( 
.A(n_1743),
.Y(n_1764)
);

BUFx8_ASAP7_75t_L g1765 ( 
.A(n_1736),
.Y(n_1765)
);

INVx4_ASAP7_75t_SL g1766 ( 
.A(n_1740),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1726),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1718),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1723),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1703),
.Y(n_1770)
);

INVx4_ASAP7_75t_L g1771 ( 
.A(n_1725),
.Y(n_1771)
);

OA21x2_ASAP7_75t_L g1772 ( 
.A1(n_1738),
.A2(n_1632),
.B(n_1659),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1737),
.Y(n_1773)
);

OAI21x1_ASAP7_75t_L g1774 ( 
.A1(n_1731),
.A2(n_1658),
.B(n_1634),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1755),
.B(n_1712),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1766),
.B(n_1719),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1745),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1745),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1752),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1767),
.B(n_1684),
.Y(n_1780)
);

NAND4xp25_ASAP7_75t_L g1781 ( 
.A(n_1758),
.B(n_1701),
.C(n_1710),
.D(n_1717),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_1765),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1753),
.Y(n_1783)
);

OAI211xp5_ASAP7_75t_L g1784 ( 
.A1(n_1764),
.A2(n_1717),
.B(n_1721),
.C(n_1712),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1752),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1766),
.B(n_1722),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1766),
.B(n_1722),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1766),
.B(n_1690),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1758),
.A2(n_1711),
.B1(n_1721),
.B2(n_1727),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1766),
.B(n_1690),
.Y(n_1790)
);

NAND2xp33_ASAP7_75t_R g1791 ( 
.A(n_1755),
.B(n_1736),
.Y(n_1791)
);

BUFx3_ASAP7_75t_L g1792 ( 
.A(n_1765),
.Y(n_1792)
);

AOI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1758),
.A2(n_1735),
.B1(n_1707),
.B2(n_1715),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1746),
.Y(n_1794)
);

INVx3_ASAP7_75t_L g1795 ( 
.A(n_1763),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1766),
.B(n_1695),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1767),
.B(n_1684),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1746),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1746),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1759),
.Y(n_1800)
);

AND2x4_ASAP7_75t_L g1801 ( 
.A(n_1766),
.B(n_1694),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1759),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1766),
.B(n_1695),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1759),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1753),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1766),
.B(n_1741),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1770),
.B(n_1741),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1767),
.B(n_1730),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1770),
.B(n_1699),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1773),
.B(n_1670),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1760),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1748),
.B(n_1747),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1748),
.B(n_1747),
.Y(n_1813)
);

NAND4xp75_ASAP7_75t_L g1814 ( 
.A(n_1772),
.B(n_1729),
.C(n_1681),
.D(n_1638),
.Y(n_1814)
);

INVx1_ASAP7_75t_SL g1815 ( 
.A(n_1761),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1760),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1760),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1764),
.B(n_1699),
.Y(n_1818)
);

INVxp67_ASAP7_75t_SL g1819 ( 
.A(n_1791),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1801),
.B(n_1747),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1794),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1794),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1801),
.B(n_1751),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1798),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1801),
.B(n_1751),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1798),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1799),
.Y(n_1827)
);

INVxp67_ASAP7_75t_L g1828 ( 
.A(n_1807),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1812),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1799),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1808),
.B(n_1773),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1800),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1800),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1802),
.Y(n_1834)
);

A2O1A1Ixp33_ASAP7_75t_L g1835 ( 
.A1(n_1781),
.A2(n_1764),
.B(n_1751),
.C(n_1762),
.Y(n_1835)
);

A2O1A1Ixp33_ASAP7_75t_L g1836 ( 
.A1(n_1784),
.A2(n_1762),
.B(n_1774),
.C(n_1704),
.Y(n_1836)
);

NOR3x1_ASAP7_75t_L g1837 ( 
.A(n_1775),
.B(n_1744),
.C(n_1761),
.Y(n_1837)
);

O2A1O1Ixp33_ASAP7_75t_SL g1838 ( 
.A1(n_1815),
.A2(n_1761),
.B(n_1762),
.C(n_1742),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1801),
.B(n_1761),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1802),
.Y(n_1840)
);

AOI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1789),
.A2(n_1765),
.B1(n_1742),
.B2(n_1636),
.Y(n_1841)
);

INVx1_ASAP7_75t_SL g1842 ( 
.A(n_1782),
.Y(n_1842)
);

NAND2x1_ASAP7_75t_SL g1843 ( 
.A(n_1793),
.B(n_1763),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1804),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1804),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1809),
.B(n_1773),
.Y(n_1846)
);

HB1xp67_ASAP7_75t_L g1847 ( 
.A(n_1812),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1818),
.B(n_1813),
.Y(n_1848)
);

OAI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1814),
.A2(n_1771),
.B1(n_1749),
.B2(n_1772),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1806),
.B(n_1749),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1777),
.Y(n_1851)
);

INVx2_ASAP7_75t_SL g1852 ( 
.A(n_1776),
.Y(n_1852)
);

NAND3xp33_ASAP7_75t_L g1853 ( 
.A(n_1777),
.B(n_1765),
.C(n_1772),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1778),
.Y(n_1854)
);

NAND2x1_ASAP7_75t_L g1855 ( 
.A(n_1776),
.B(n_1749),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_SL g1856 ( 
.A1(n_1819),
.A2(n_1792),
.B1(n_1782),
.B2(n_1813),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1823),
.B(n_1806),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1828),
.B(n_1778),
.Y(n_1858)
);

OAI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1835),
.A2(n_1814),
.B1(n_1792),
.B2(n_1749),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1847),
.Y(n_1860)
);

INVx1_ASAP7_75t_SL g1861 ( 
.A(n_1842),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_L g1862 ( 
.A1(n_1841),
.A2(n_1853),
.B1(n_1850),
.B2(n_1849),
.Y(n_1862)
);

AOI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1835),
.A2(n_1765),
.B1(n_1772),
.B2(n_1630),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1829),
.B(n_1779),
.Y(n_1864)
);

OAI221xp5_ASAP7_75t_L g1865 ( 
.A1(n_1836),
.A2(n_1779),
.B1(n_1785),
.B2(n_1795),
.C(n_1772),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1829),
.B(n_1837),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1823),
.B(n_1786),
.Y(n_1867)
);

INVxp67_ASAP7_75t_SL g1868 ( 
.A(n_1843),
.Y(n_1868)
);

HB1xp67_ASAP7_75t_L g1869 ( 
.A(n_1831),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1848),
.B(n_1785),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1850),
.A2(n_1825),
.B1(n_1852),
.B2(n_1820),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1846),
.B(n_1780),
.Y(n_1872)
);

INVx1_ASAP7_75t_SL g1873 ( 
.A(n_1825),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1821),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1839),
.B(n_1786),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1839),
.B(n_1787),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1820),
.B(n_1787),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1851),
.B(n_1754),
.Y(n_1878)
);

INVxp67_ASAP7_75t_L g1879 ( 
.A(n_1854),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1852),
.B(n_1788),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1846),
.B(n_1780),
.Y(n_1881)
);

OAI22xp33_ASAP7_75t_L g1882 ( 
.A1(n_1868),
.A2(n_1836),
.B1(n_1795),
.B2(n_1855),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1860),
.Y(n_1883)
);

AOI311xp33_ASAP7_75t_L g1884 ( 
.A1(n_1865),
.A2(n_1838),
.A3(n_1845),
.B(n_1840),
.C(n_1844),
.Y(n_1884)
);

OAI32xp33_ASAP7_75t_L g1885 ( 
.A1(n_1866),
.A2(n_1795),
.A3(n_1838),
.B1(n_1833),
.B2(n_1832),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1862),
.A2(n_1772),
.B1(n_1830),
.B2(n_1827),
.Y(n_1886)
);

BUFx3_ASAP7_75t_L g1887 ( 
.A(n_1861),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1860),
.Y(n_1888)
);

AOI221x1_ASAP7_75t_SL g1889 ( 
.A1(n_1859),
.A2(n_1834),
.B1(n_1826),
.B2(n_1824),
.C(n_1822),
.Y(n_1889)
);

AOI21xp33_ASAP7_75t_L g1890 ( 
.A1(n_1856),
.A2(n_1765),
.B(n_1810),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1873),
.B(n_1808),
.Y(n_1891)
);

BUFx2_ASAP7_75t_L g1892 ( 
.A(n_1869),
.Y(n_1892)
);

O2A1O1Ixp33_ASAP7_75t_SL g1893 ( 
.A1(n_1863),
.A2(n_1810),
.B(n_1768),
.C(n_1769),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1864),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1870),
.B(n_1797),
.Y(n_1895)
);

OAI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1863),
.A2(n_1749),
.B1(n_1771),
.B2(n_1796),
.Y(n_1896)
);

AOI222xp33_ASAP7_75t_L g1897 ( 
.A1(n_1858),
.A2(n_1879),
.B1(n_1871),
.B2(n_1874),
.C1(n_1857),
.C2(n_1878),
.Y(n_1897)
);

OAI221xp5_ASAP7_75t_SL g1898 ( 
.A1(n_1870),
.A2(n_1733),
.B1(n_1750),
.B2(n_1788),
.C(n_1790),
.Y(n_1898)
);

O2A1O1Ixp5_ASAP7_75t_SL g1899 ( 
.A1(n_1874),
.A2(n_1817),
.B(n_1816),
.C(n_1811),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1857),
.B(n_1754),
.Y(n_1900)
);

AO22x1_ASAP7_75t_L g1901 ( 
.A1(n_1867),
.A2(n_1765),
.B1(n_1749),
.B2(n_1771),
.Y(n_1901)
);

AOI22xp33_ASAP7_75t_L g1902 ( 
.A1(n_1886),
.A2(n_1867),
.B1(n_1877),
.B2(n_1880),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1892),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1887),
.B(n_1877),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1894),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1891),
.B(n_1872),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1897),
.B(n_1875),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1889),
.B(n_1875),
.Y(n_1908)
);

HB1xp67_ASAP7_75t_L g1909 ( 
.A(n_1895),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1890),
.B(n_1876),
.Y(n_1910)
);

NOR2xp33_ASAP7_75t_L g1911 ( 
.A(n_1883),
.B(n_1864),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1888),
.Y(n_1912)
);

AOI211xp5_ASAP7_75t_L g1913 ( 
.A1(n_1908),
.A2(n_1885),
.B(n_1882),
.C(n_1898),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1906),
.B(n_1900),
.Y(n_1914)
);

AOI221xp5_ASAP7_75t_L g1915 ( 
.A1(n_1907),
.A2(n_1886),
.B1(n_1882),
.B2(n_1898),
.C(n_1893),
.Y(n_1915)
);

AOI31xp33_ASAP7_75t_SL g1916 ( 
.A1(n_1904),
.A2(n_1884),
.A3(n_1872),
.B(n_1881),
.Y(n_1916)
);

AOI221xp5_ASAP7_75t_L g1917 ( 
.A1(n_1907),
.A2(n_1896),
.B1(n_1901),
.B2(n_1880),
.C(n_1876),
.Y(n_1917)
);

NOR3xp33_ASAP7_75t_L g1918 ( 
.A(n_1903),
.B(n_1881),
.C(n_1771),
.Y(n_1918)
);

NAND3xp33_ASAP7_75t_SL g1919 ( 
.A(n_1902),
.B(n_1899),
.C(n_1796),
.Y(n_1919)
);

AOI211xp5_ASAP7_75t_L g1920 ( 
.A1(n_1909),
.A2(n_1774),
.B(n_1790),
.C(n_1803),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_SL g1921 ( 
.A(n_1902),
.B(n_1910),
.Y(n_1921)
);

NAND2xp33_ASAP7_75t_SL g1922 ( 
.A(n_1905),
.B(n_1749),
.Y(n_1922)
);

OAI221xp5_ASAP7_75t_L g1923 ( 
.A1(n_1911),
.A2(n_1771),
.B1(n_1772),
.B2(n_1803),
.C(n_1750),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1914),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1921),
.Y(n_1925)
);

A2O1A1Ixp33_ASAP7_75t_SL g1926 ( 
.A1(n_1913),
.A2(n_1911),
.B(n_1912),
.C(n_1805),
.Y(n_1926)
);

O2A1O1Ixp5_ASAP7_75t_L g1927 ( 
.A1(n_1922),
.A2(n_1783),
.B(n_1805),
.C(n_1750),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_SL g1928 ( 
.A(n_1919),
.B(n_1771),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1916),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1924),
.Y(n_1930)
);

INVxp67_ASAP7_75t_SL g1931 ( 
.A(n_1925),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_SL g1932 ( 
.A(n_1929),
.B(n_1918),
.Y(n_1932)
);

NAND2x1_ASAP7_75t_SL g1933 ( 
.A(n_1926),
.B(n_1917),
.Y(n_1933)
);

INVxp67_ASAP7_75t_SL g1934 ( 
.A(n_1928),
.Y(n_1934)
);

NOR3xp33_ASAP7_75t_L g1935 ( 
.A(n_1927),
.B(n_1915),
.C(n_1923),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1934),
.B(n_1931),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1933),
.B(n_1928),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1930),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1932),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1935),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1939),
.B(n_1920),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_SL g1942 ( 
.A(n_1937),
.B(n_1936),
.Y(n_1942)
);

HB1xp67_ASAP7_75t_L g1943 ( 
.A(n_1938),
.Y(n_1943)
);

XNOR2xp5_ASAP7_75t_L g1944 ( 
.A(n_1941),
.B(n_1940),
.Y(n_1944)
);

NOR2x1_ASAP7_75t_L g1945 ( 
.A(n_1944),
.B(n_1942),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1945),
.Y(n_1946)
);

CKINVDCx20_ASAP7_75t_R g1947 ( 
.A(n_1945),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1946),
.B(n_1943),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1947),
.B(n_1783),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1948),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1950),
.Y(n_1951)
);

OAI222xp33_ASAP7_75t_L g1952 ( 
.A1(n_1951),
.A2(n_1949),
.B1(n_1817),
.B2(n_1816),
.C1(n_1811),
.C2(n_1750),
.Y(n_1952)
);

AOI21xp5_ASAP7_75t_L g1953 ( 
.A1(n_1952),
.A2(n_1750),
.B(n_1757),
.Y(n_1953)
);

AOI22x1_ASAP7_75t_L g1954 ( 
.A1(n_1953),
.A2(n_1756),
.B1(n_1757),
.B2(n_1768),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1954),
.A2(n_1797),
.B1(n_1768),
.B2(n_1769),
.Y(n_1955)
);

AOI211xp5_ASAP7_75t_L g1956 ( 
.A1(n_1955),
.A2(n_1774),
.B(n_1768),
.C(n_1769),
.Y(n_1956)
);


endmodule