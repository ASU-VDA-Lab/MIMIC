module real_aes_1494_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_756, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_757, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_756;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_757;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g177 ( .A(n_0), .B(n_151), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_1), .B(n_108), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_2), .B(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_3), .B(n_135), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_4), .B(n_153), .Y(n_464) );
INVx1_ASAP7_75t_L g142 ( .A(n_5), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_6), .B(n_135), .Y(n_204) );
NAND2xp33_ASAP7_75t_SL g247 ( .A(n_7), .B(n_141), .Y(n_247) );
XNOR2xp5_ASAP7_75t_L g115 ( .A(n_8), .B(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g239 ( .A(n_9), .Y(n_239) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_10), .Y(n_108) );
AND2x2_ASAP7_75t_L g202 ( .A(n_11), .B(n_159), .Y(n_202) );
AND2x2_ASAP7_75t_L g466 ( .A(n_12), .B(n_155), .Y(n_466) );
AND2x2_ASAP7_75t_L g476 ( .A(n_13), .B(n_245), .Y(n_476) );
INVx2_ASAP7_75t_L g157 ( .A(n_14), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_15), .B(n_153), .Y(n_516) );
NOR3xp33_ASAP7_75t_L g106 ( .A(n_16), .B(n_107), .C(n_109), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g124 ( .A(n_16), .Y(n_124) );
AOI221x1_ASAP7_75t_L g242 ( .A1(n_17), .A2(n_144), .B1(n_243), .B2(n_245), .C(n_246), .Y(n_242) );
AOI22xp5_ASAP7_75t_SL g116 ( .A1(n_18), .A2(n_75), .B1(n_117), .B2(n_118), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_18), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g134 ( .A(n_19), .B(n_135), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_20), .B(n_135), .Y(n_521) );
INVx1_ASAP7_75t_L g112 ( .A(n_21), .Y(n_112) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_22), .A2(n_92), .B1(n_135), .B2(n_188), .Y(n_480) );
AOI221xp5_ASAP7_75t_SL g166 ( .A1(n_23), .A2(n_39), .B1(n_135), .B2(n_144), .C(n_167), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_24), .A2(n_144), .B(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_25), .B(n_151), .Y(n_207) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_26), .A2(n_91), .B(n_157), .Y(n_156) );
OR2x2_ASAP7_75t_L g160 ( .A(n_26), .B(n_91), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_27), .B(n_153), .Y(n_152) );
INVxp67_ASAP7_75t_L g241 ( .A(n_28), .Y(n_241) );
AND2x2_ASAP7_75t_L g228 ( .A(n_29), .B(n_165), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_30), .A2(n_144), .B(n_176), .Y(n_175) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_31), .A2(n_245), .B(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_32), .B(n_153), .Y(n_168) );
OAI22xp5_ASAP7_75t_SL g743 ( .A1(n_33), .A2(n_72), .B1(n_744), .B2(n_745), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_33), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_34), .A2(n_144), .B(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_35), .B(n_153), .Y(n_536) );
AND2x2_ASAP7_75t_L g141 ( .A(n_36), .B(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_L g145 ( .A(n_36), .B(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g196 ( .A(n_36), .Y(n_196) );
INVxp67_ASAP7_75t_L g109 ( .A(n_37), .Y(n_109) );
OR2x6_ASAP7_75t_L g125 ( .A(n_37), .B(n_126), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_38), .A2(n_741), .B1(n_742), .B2(n_746), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_38), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_40), .B(n_135), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_41), .A2(n_83), .B1(n_144), .B2(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_42), .B(n_153), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_43), .B(n_135), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_44), .B(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_45), .B(n_151), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_46), .A2(n_144), .B(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g180 ( .A(n_47), .B(n_165), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_48), .B(n_151), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_49), .B(n_165), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_50), .B(n_135), .Y(n_513) );
INVx1_ASAP7_75t_L g138 ( .A(n_51), .Y(n_138) );
INVx1_ASAP7_75t_L g148 ( .A(n_51), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_52), .B(n_153), .Y(n_474) );
AND2x2_ASAP7_75t_L g503 ( .A(n_53), .B(n_165), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_54), .B(n_135), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_55), .B(n_151), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_56), .B(n_151), .Y(n_535) );
AND2x2_ASAP7_75t_L g219 ( .A(n_57), .B(n_165), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_58), .B(n_135), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_59), .B(n_153), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_60), .B(n_135), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_61), .A2(n_144), .B(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_62), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_63), .B(n_151), .Y(n_216) );
AND2x2_ASAP7_75t_L g527 ( .A(n_64), .B(n_159), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_65), .A2(n_144), .B(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_66), .B(n_153), .Y(n_208) );
AND2x2_ASAP7_75t_SL g199 ( .A(n_67), .B(n_155), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_68), .B(n_151), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_69), .B(n_151), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_70), .A2(n_94), .B1(n_144), .B2(n_194), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_71), .B(n_153), .Y(n_524) );
INVx1_ASAP7_75t_L g744 ( .A(n_72), .Y(n_744) );
INVx1_ASAP7_75t_L g140 ( .A(n_73), .Y(n_140) );
INVx1_ASAP7_75t_L g146 ( .A(n_73), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_74), .B(n_151), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_75), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_76), .A2(n_144), .B(n_507), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_77), .A2(n_144), .B(n_454), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_78), .A2(n_144), .B(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g538 ( .A(n_79), .B(n_159), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_80), .B(n_165), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_81), .A2(n_85), .B1(n_135), .B2(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_82), .B(n_135), .Y(n_217) );
INVx1_ASAP7_75t_L g111 ( .A(n_84), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_86), .B(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_87), .B(n_151), .Y(n_169) );
AND2x2_ASAP7_75t_L g457 ( .A(n_88), .B(n_155), .Y(n_457) );
INVxp33_ASAP7_75t_L g753 ( .A(n_89), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_90), .A2(n_144), .B(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_93), .B(n_153), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_95), .A2(n_144), .B(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_96), .B(n_153), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_97), .B(n_135), .Y(n_179) );
INVxp67_ASAP7_75t_L g244 ( .A(n_98), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_99), .B(n_153), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_100), .A2(n_144), .B(n_149), .Y(n_143) );
BUFx2_ASAP7_75t_L g526 ( .A(n_101), .Y(n_526) );
NAND3xp33_ASAP7_75t_SL g731 ( .A(n_102), .B(n_732), .C(n_736), .Y(n_731) );
INVx1_ASAP7_75t_SL g748 ( .A(n_102), .Y(n_748) );
BUFx2_ASAP7_75t_L g751 ( .A(n_102), .Y(n_751) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_113), .B(n_752), .Y(n_103) );
CKINVDCx6p67_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
INVx3_ASAP7_75t_SL g754 ( .A(n_105), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g105 ( .A(n_106), .B(n_110), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_111), .B(n_112), .Y(n_126) );
OA331x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_729), .A3(n_731), .B1(n_739), .B2(n_740), .B3(n_747), .C1(n_749), .Y(n_113) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_119), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_115), .B(n_730), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_127), .B1(n_441), .B2(n_725), .Y(n_119) );
INVx4_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
INVx3_ASAP7_75t_SL g121 ( .A(n_122), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_123), .Y(n_122) );
AOI22xp5_ASAP7_75t_SL g730 ( .A1(n_123), .A2(n_127), .B1(n_441), .B2(n_726), .Y(n_730) );
AND2x6_ASAP7_75t_SL g123 ( .A(n_124), .B(n_125), .Y(n_123) );
OR2x6_ASAP7_75t_SL g727 ( .A(n_124), .B(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_124), .B(n_728), .Y(n_735) );
OR2x2_ASAP7_75t_L g738 ( .A(n_124), .B(n_125), .Y(n_738) );
CKINVDCx5p33_ASAP7_75t_R g728 ( .A(n_125), .Y(n_728) );
XNOR2xp5_ASAP7_75t_L g742 ( .A(n_127), .B(n_743), .Y(n_742) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_333), .Y(n_127) );
NOR3xp33_ASAP7_75t_L g128 ( .A(n_129), .B(n_261), .C(n_311), .Y(n_128) );
OAI211xp5_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_181), .B(n_229), .C(n_250), .Y(n_129) );
OR2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_161), .Y(n_130) );
AND2x2_ASAP7_75t_L g260 ( .A(n_131), .B(n_162), .Y(n_260) );
INVx1_ASAP7_75t_L g391 ( .A(n_131), .Y(n_391) );
NOR2x1p5_ASAP7_75t_L g423 ( .A(n_131), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g234 ( .A(n_132), .B(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g282 ( .A(n_132), .Y(n_282) );
OR2x2_ASAP7_75t_L g286 ( .A(n_132), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_132), .B(n_164), .Y(n_298) );
OR2x2_ASAP7_75t_L g320 ( .A(n_132), .B(n_164), .Y(n_320) );
AND2x4_ASAP7_75t_L g326 ( .A(n_132), .B(n_290), .Y(n_326) );
OR2x2_ASAP7_75t_L g343 ( .A(n_132), .B(n_236), .Y(n_343) );
INVx1_ASAP7_75t_L g378 ( .A(n_132), .Y(n_378) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_132), .Y(n_400) );
OR2x2_ASAP7_75t_L g414 ( .A(n_132), .B(n_347), .Y(n_414) );
AND2x4_ASAP7_75t_SL g418 ( .A(n_132), .B(n_236), .Y(n_418) );
OR2x6_ASAP7_75t_L g132 ( .A(n_133), .B(n_158), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_143), .B(n_155), .Y(n_133) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_141), .Y(n_135) );
INVx1_ASAP7_75t_L g248 ( .A(n_136), .Y(n_248) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
AND2x6_ASAP7_75t_L g151 ( .A(n_137), .B(n_146), .Y(n_151) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x4_ASAP7_75t_L g153 ( .A(n_139), .B(n_148), .Y(n_153) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx5_ASAP7_75t_L g154 ( .A(n_141), .Y(n_154) );
AND2x2_ASAP7_75t_L g147 ( .A(n_142), .B(n_148), .Y(n_147) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_142), .Y(n_191) );
AND2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
BUFx3_ASAP7_75t_L g192 ( .A(n_145), .Y(n_192) );
INVx2_ASAP7_75t_L g198 ( .A(n_146), .Y(n_198) );
AND2x4_ASAP7_75t_L g194 ( .A(n_147), .B(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g190 ( .A(n_148), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_152), .B(n_154), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_151), .B(n_526), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_154), .A2(n_168), .B(n_169), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_154), .A2(n_177), .B(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_154), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_154), .A2(n_215), .B(n_216), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_154), .A2(n_225), .B(n_226), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_154), .A2(n_455), .B(n_456), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_154), .A2(n_463), .B(n_464), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_154), .A2(n_473), .B(n_474), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_154), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_154), .A2(n_516), .B(n_517), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_154), .A2(n_524), .B(n_525), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_154), .A2(n_535), .B(n_536), .Y(n_534) );
INVx2_ASAP7_75t_SL g185 ( .A(n_155), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_155), .A2(n_521), .B(n_522), .Y(n_520) );
BUFx4f_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx3_ASAP7_75t_L g173 ( .A(n_156), .Y(n_173) );
AND2x2_ASAP7_75t_SL g159 ( .A(n_157), .B(n_160), .Y(n_159) );
AND2x4_ASAP7_75t_L g209 ( .A(n_157), .B(n_160), .Y(n_209) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_159), .Y(n_165) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g370 ( .A(n_162), .B(n_326), .Y(n_370) );
AND2x2_ASAP7_75t_L g417 ( .A(n_162), .B(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g162 ( .A(n_163), .B(n_171), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g233 ( .A(n_164), .Y(n_233) );
AND2x2_ASAP7_75t_L g280 ( .A(n_164), .B(n_171), .Y(n_280) );
INVx2_ASAP7_75t_L g287 ( .A(n_164), .Y(n_287) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_164), .Y(n_408) );
BUFx3_ASAP7_75t_L g424 ( .A(n_164), .Y(n_424) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_170), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_165), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_165), .A2(n_452), .B(n_453), .Y(n_451) );
AO21x2_ASAP7_75t_L g479 ( .A1(n_165), .A2(n_480), .B(n_481), .Y(n_479) );
INVx2_ASAP7_75t_L g249 ( .A(n_171), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_171), .B(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g347 ( .A(n_171), .B(n_287), .Y(n_347) );
INVx1_ASAP7_75t_L g365 ( .A(n_171), .Y(n_365) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_171), .Y(n_381) );
INVx1_ASAP7_75t_L g403 ( .A(n_171), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_171), .B(n_282), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_171), .B(n_236), .Y(n_440) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AOI21x1_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_180), .Y(n_172) );
INVx4_ASAP7_75t_L g245 ( .A(n_173), .Y(n_245) );
AO21x2_ASAP7_75t_L g469 ( .A1(n_173), .A2(n_470), .B(n_476), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_175), .B(n_179), .Y(n_174) );
INVx1_ASAP7_75t_SL g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_200), .Y(n_182) );
AND2x4_ASAP7_75t_L g254 ( .A(n_183), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g265 ( .A(n_183), .Y(n_265) );
AND2x2_ASAP7_75t_L g270 ( .A(n_183), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g305 ( .A(n_183), .B(n_210), .Y(n_305) );
AND2x2_ASAP7_75t_L g315 ( .A(n_183), .B(n_211), .Y(n_315) );
OR2x2_ASAP7_75t_L g395 ( .A(n_183), .B(n_310), .Y(n_395) );
OAI322xp33_ASAP7_75t_L g425 ( .A1(n_183), .A2(n_338), .A3(n_377), .B1(n_410), .B2(n_426), .C1(n_427), .C2(n_428), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_183), .B(n_408), .Y(n_426) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g259 ( .A(n_184), .Y(n_259) );
AOI21x1_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_199), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_193), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_188), .A2(n_194), .B1(n_238), .B2(n_240), .Y(n_237) );
AND2x4_ASAP7_75t_L g188 ( .A(n_189), .B(n_192), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
NOR2x1p5_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
INVx3_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_200), .A2(n_372), .B1(n_376), .B2(n_379), .Y(n_371) );
AOI211xp5_ASAP7_75t_L g431 ( .A1(n_200), .A2(n_432), .B(n_433), .C(n_436), .Y(n_431) );
AND2x4_ASAP7_75t_SL g200 ( .A(n_201), .B(n_210), .Y(n_200) );
AND2x4_ASAP7_75t_L g253 ( .A(n_201), .B(n_221), .Y(n_253) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_201), .Y(n_257) );
INVx5_ASAP7_75t_L g269 ( .A(n_201), .Y(n_269) );
INVx2_ASAP7_75t_L g278 ( .A(n_201), .Y(n_278) );
AND2x2_ASAP7_75t_L g301 ( .A(n_201), .B(n_211), .Y(n_301) );
AND2x2_ASAP7_75t_L g330 ( .A(n_201), .B(n_220), .Y(n_330) );
OR2x2_ASAP7_75t_L g339 ( .A(n_201), .B(n_259), .Y(n_339) );
OR2x2_ASAP7_75t_L g354 ( .A(n_201), .B(n_268), .Y(n_354) );
OR2x6_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_209), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_209), .B(n_239), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_209), .B(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_209), .B(n_244), .Y(n_243) );
NOR3xp33_ASAP7_75t_L g246 ( .A(n_209), .B(n_247), .C(n_248), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_209), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_209), .A2(n_513), .B(n_514), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_210), .B(n_230), .Y(n_229) );
INVx3_ASAP7_75t_SL g338 ( .A(n_210), .Y(n_338) );
AND2x2_ASAP7_75t_L g361 ( .A(n_210), .B(n_269), .Y(n_361) );
AND2x4_ASAP7_75t_L g210 ( .A(n_211), .B(n_220), .Y(n_210) );
INVx2_ASAP7_75t_L g255 ( .A(n_211), .Y(n_255) );
AND2x2_ASAP7_75t_L g258 ( .A(n_211), .B(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g272 ( .A(n_211), .B(n_221), .Y(n_272) );
INVx1_ASAP7_75t_L g276 ( .A(n_211), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_211), .B(n_221), .Y(n_310) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_211), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_211), .B(n_269), .Y(n_385) );
AO21x2_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_218), .B(n_219), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_213), .B(n_217), .Y(n_212) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_218), .A2(n_222), .B(n_228), .Y(n_221) );
AO21x2_ASAP7_75t_L g268 ( .A1(n_218), .A2(n_222), .B(n_228), .Y(n_268) );
AOI21x1_ASAP7_75t_L g459 ( .A1(n_218), .A2(n_460), .B(n_466), .Y(n_459) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_221), .Y(n_291) );
AND2x2_ASAP7_75t_L g375 ( .A(n_221), .B(n_259), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_227), .Y(n_222) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_234), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_231), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
OR2x6_ASAP7_75t_SL g439 ( .A(n_232), .B(n_440), .Y(n_439) );
INVxp67_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_233), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_233), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g387 ( .A(n_233), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_234), .A2(n_296), .B1(n_299), .B2(n_306), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_235), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g331 ( .A(n_235), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_235), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_SL g386 ( .A(n_235), .B(n_387), .Y(n_386) );
AND2x4_ASAP7_75t_L g235 ( .A(n_236), .B(n_249), .Y(n_235) );
AND2x2_ASAP7_75t_L g281 ( .A(n_236), .B(n_282), .Y(n_281) );
INVx3_ASAP7_75t_L g290 ( .A(n_236), .Y(n_290) );
OAI22xp33_ASAP7_75t_L g348 ( .A1(n_236), .A2(n_297), .B1(n_349), .B2(n_351), .Y(n_348) );
INVx1_ASAP7_75t_L g356 ( .A(n_236), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_236), .B(n_350), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_236), .B(n_280), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_236), .B(n_287), .Y(n_429) );
AND2x4_ASAP7_75t_L g236 ( .A(n_237), .B(n_242), .Y(n_236) );
INVx3_ASAP7_75t_L g531 ( .A(n_245), .Y(n_531) );
OAI21xp33_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_256), .B(n_260), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
NAND4xp25_ASAP7_75t_SL g299 ( .A(n_252), .B(n_300), .C(n_302), .D(n_304), .Y(n_299) );
INVx2_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_253), .B(n_360), .Y(n_389) );
AND2x2_ASAP7_75t_L g416 ( .A(n_253), .B(n_254), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_253), .B(n_276), .Y(n_427) );
INVx1_ASAP7_75t_L g292 ( .A(n_254), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g327 ( .A1(n_254), .A2(n_317), .B1(n_328), .B2(n_331), .Y(n_327) );
NAND3xp33_ASAP7_75t_L g349 ( .A(n_254), .B(n_267), .C(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_254), .B(n_269), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_254), .B(n_277), .Y(n_420) );
AND2x2_ASAP7_75t_L g352 ( .A(n_255), .B(n_259), .Y(n_352) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_255), .Y(n_413) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
INVx1_ASAP7_75t_L g308 ( .A(n_257), .Y(n_308) );
INVx1_ASAP7_75t_L g398 ( .A(n_258), .Y(n_398) );
AND2x2_ASAP7_75t_L g405 ( .A(n_258), .B(n_269), .Y(n_405) );
BUFx2_ASAP7_75t_L g360 ( .A(n_259), .Y(n_360) );
NAND3xp33_ASAP7_75t_SL g261 ( .A(n_262), .B(n_283), .C(n_295), .Y(n_261) );
OAI31xp33_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_270), .A3(n_273), .B(n_279), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_263), .A2(n_317), .B1(n_321), .B2(n_322), .Y(n_316) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
OR2x2_ASAP7_75t_L g302 ( .A(n_265), .B(n_303), .Y(n_302) );
NOR2x1_ASAP7_75t_L g328 ( .A(n_265), .B(n_329), .Y(n_328) );
O2A1O1Ixp33_ASAP7_75t_L g397 ( .A1(n_266), .A2(n_368), .B(n_398), .C(n_399), .Y(n_397) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_267), .B(n_413), .Y(n_412) );
AND2x4_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_268), .B(n_276), .Y(n_303) );
AND2x2_ASAP7_75t_L g321 ( .A(n_268), .B(n_301), .Y(n_321) );
AND2x2_ASAP7_75t_L g438 ( .A(n_271), .B(n_360), .Y(n_438) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g294 ( .A(n_272), .B(n_278), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_274), .B(n_277), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_277), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g369 ( .A(n_277), .B(n_352), .Y(n_369) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_278), .B(n_352), .Y(n_358) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx2_ASAP7_75t_L g350 ( .A(n_280), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_281), .B(n_381), .Y(n_380) );
AOI32xp33_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_291), .A3(n_292), .B1(n_293), .B2(n_756), .Y(n_283) );
AOI221xp5_ASAP7_75t_L g404 ( .A1(n_284), .A2(n_369), .B1(n_405), .B2(n_406), .C(n_409), .Y(n_404) );
AND2x4_ASAP7_75t_L g284 ( .A(n_285), .B(n_288), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_287), .Y(n_332) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g297 ( .A(n_289), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g402 ( .A(n_290), .B(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_291), .B(n_313), .Y(n_312) );
AOI221xp5_ASAP7_75t_L g335 ( .A1(n_293), .A2(n_336), .B1(n_340), .B2(n_344), .C(n_348), .Y(n_335) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OAI211xp5_ASAP7_75t_L g311 ( .A1(n_298), .A2(n_312), .B(n_316), .C(n_327), .Y(n_311) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OAI322xp33_ASAP7_75t_L g409 ( .A1(n_304), .A2(n_314), .A3(n_363), .B1(n_410), .B2(n_411), .C1(n_412), .C2(n_414), .Y(n_409) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AOI21xp33_ASAP7_75t_L g436 ( .A1(n_307), .A2(n_437), .B(n_439), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
O2A1O1Ixp33_ASAP7_75t_L g393 ( .A1(n_313), .A2(n_394), .B(n_396), .C(n_397), .Y(n_393) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g435 ( .A(n_320), .B(n_401), .Y(n_435) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
INVxp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_326), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g410 ( .A(n_326), .Y(n_410) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OAI31xp33_ASAP7_75t_L g366 ( .A1(n_330), .A2(n_367), .A3(n_369), .B(n_370), .Y(n_366) );
NOR2x1_ASAP7_75t_L g333 ( .A(n_334), .B(n_392), .Y(n_333) );
NAND5xp2_ASAP7_75t_L g334 ( .A(n_335), .B(n_355), .C(n_366), .D(n_371), .E(n_382), .Y(n_334) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
AOI21xp33_ASAP7_75t_L g433 ( .A1(n_338), .A2(n_434), .B(n_435), .Y(n_433) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g406 ( .A(n_342), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
A2O1A1Ixp33_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_357), .B(n_359), .C(n_362), .Y(n_355) );
INVxp33_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
OR2x2_ASAP7_75t_L g384 ( .A(n_360), .B(n_385), .Y(n_384) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_363), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_SL g372 ( .A(n_373), .B(n_375), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g434 ( .A(n_375), .Y(n_434) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_386), .B(n_388), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI21xp33_ASAP7_75t_L g388 ( .A1(n_384), .A2(n_389), .B(n_390), .Y(n_388) );
NAND4xp25_ASAP7_75t_L g392 ( .A(n_393), .B(n_404), .C(n_415), .D(n_431), .Y(n_392) );
INVx1_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_402), .B(n_423), .Y(n_422) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g432 ( .A(n_414), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_417), .B1(n_419), .B2(n_421), .C(n_425), .Y(n_415) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AND2x4_ASAP7_75t_L g441 ( .A(n_442), .B(n_638), .Y(n_441) );
NOR4xp75_ASAP7_75t_L g442 ( .A(n_443), .B(n_561), .C(n_586), .D(n_613), .Y(n_442) );
OAI21xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_498), .B(n_539), .Y(n_443) );
NOR4xp25_ASAP7_75t_L g444 ( .A(n_445), .B(n_482), .C(n_489), .D(n_493), .Y(n_444) );
INVx1_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_447), .B(n_467), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_458), .Y(n_448) );
NAND2x1p5_ASAP7_75t_L g601 ( .A(n_449), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_449), .B(n_486), .Y(n_632) );
AND2x2_ASAP7_75t_L g657 ( .A(n_449), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g682 ( .A(n_449), .B(n_477), .Y(n_682) );
AND2x2_ASAP7_75t_L g723 ( .A(n_449), .B(n_491), .Y(n_723) );
INVx4_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AND2x4_ASAP7_75t_SL g495 ( .A(n_450), .B(n_488), .Y(n_495) );
AND2x2_ASAP7_75t_L g497 ( .A(n_450), .B(n_469), .Y(n_497) );
NOR2x1_ASAP7_75t_L g547 ( .A(n_450), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g558 ( .A(n_450), .Y(n_558) );
AND2x2_ASAP7_75t_L g564 ( .A(n_450), .B(n_491), .Y(n_564) );
BUFx2_ASAP7_75t_L g577 ( .A(n_450), .Y(n_577) );
AND2x4_ASAP7_75t_L g608 ( .A(n_450), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g655 ( .A(n_450), .B(n_656), .Y(n_655) );
OR2x6_ASAP7_75t_L g450 ( .A(n_451), .B(n_457), .Y(n_450) );
INVx1_ASAP7_75t_L g649 ( .A(n_458), .Y(n_649) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx3_ASAP7_75t_L g488 ( .A(n_459), .Y(n_488) );
AND2x2_ASAP7_75t_L g491 ( .A(n_459), .B(n_469), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_465), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_467), .B(n_667), .Y(n_720) );
INVx2_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
OR2x2_ASAP7_75t_L g557 ( .A(n_468), .B(n_558), .Y(n_557) );
OR2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_477), .Y(n_468) );
INVx2_ASAP7_75t_L g487 ( .A(n_469), .Y(n_487) );
INVx2_ASAP7_75t_L g548 ( .A(n_469), .Y(n_548) );
AND2x2_ASAP7_75t_L g658 ( .A(n_469), .B(n_488), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_475), .Y(n_470) );
INVx2_ASAP7_75t_L g546 ( .A(n_477), .Y(n_546) );
BUFx3_ASAP7_75t_L g563 ( .A(n_477), .Y(n_563) );
AND2x2_ASAP7_75t_L g590 ( .A(n_477), .B(n_591), .Y(n_590) );
AND2x4_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
AND2x4_ASAP7_75t_L g484 ( .A(n_478), .B(n_479), .Y(n_484) );
NOR2x1_ASAP7_75t_L g482 ( .A(n_483), .B(n_485), .Y(n_482) );
INVx2_ASAP7_75t_L g492 ( .A(n_483), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_483), .B(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g661 ( .A(n_483), .B(n_601), .Y(n_661) );
AND2x2_ASAP7_75t_L g685 ( .A(n_483), .B(n_495), .Y(n_685) );
INVx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g581 ( .A(n_484), .B(n_487), .Y(n_581) );
AND2x2_ASAP7_75t_L g663 ( .A(n_484), .B(n_656), .Y(n_663) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_SL g706 ( .A(n_486), .Y(n_706) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g591 ( .A(n_487), .Y(n_591) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_488), .Y(n_595) );
INVx2_ASAP7_75t_L g603 ( .A(n_488), .Y(n_603) );
INVx1_ASAP7_75t_L g609 ( .A(n_488), .Y(n_609) );
AOI222xp33_ASAP7_75t_SL g539 ( .A1(n_489), .A2(n_540), .B1(n_544), .B2(n_549), .C1(n_556), .C2(n_559), .Y(n_539) );
INVx1_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g616 ( .A(n_491), .Y(n_616) );
BUFx2_ASAP7_75t_L g645 ( .A(n_491), .Y(n_645) );
OAI211xp5_ASAP7_75t_L g639 ( .A1(n_492), .A2(n_640), .B(n_644), .C(n_652), .Y(n_639) );
OR2x2_ASAP7_75t_L g710 ( .A(n_492), .B(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g718 ( .A(n_492), .B(n_623), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_496), .Y(n_493) );
INVx2_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_SL g675 ( .A(n_495), .B(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g693 ( .A(n_495), .B(n_581), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_495), .B(n_673), .Y(n_700) );
OR2x2_ASAP7_75t_L g701 ( .A(n_496), .B(n_563), .Y(n_701) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g623 ( .A(n_497), .B(n_595), .Y(n_623) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_518), .Y(n_499) );
INVx1_ASAP7_75t_L g717 ( .A(n_500), .Y(n_717) );
NOR2xp67_ASAP7_75t_L g500 ( .A(n_501), .B(n_510), .Y(n_500) );
AND2x2_ASAP7_75t_L g560 ( .A(n_501), .B(n_519), .Y(n_560) );
INVx1_ASAP7_75t_L g637 ( .A(n_501), .Y(n_637) );
OR2x2_ASAP7_75t_L g696 ( .A(n_501), .B(n_519), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_501), .B(n_568), .Y(n_702) );
INVx4_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g543 ( .A(n_502), .Y(n_543) );
OR2x2_ASAP7_75t_L g575 ( .A(n_502), .B(n_529), .Y(n_575) );
AND2x2_ASAP7_75t_L g584 ( .A(n_502), .B(n_511), .Y(n_584) );
NAND2x1_ASAP7_75t_L g612 ( .A(n_502), .B(n_519), .Y(n_612) );
AND2x2_ASAP7_75t_L g659 ( .A(n_502), .B(n_554), .Y(n_659) );
OR2x6_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g542 ( .A(n_511), .Y(n_542) );
INVx1_ASAP7_75t_L g552 ( .A(n_511), .Y(n_552) );
AND2x2_ASAP7_75t_L g568 ( .A(n_511), .B(n_555), .Y(n_568) );
INVx2_ASAP7_75t_L g573 ( .A(n_511), .Y(n_573) );
OR2x2_ASAP7_75t_L g669 ( .A(n_511), .B(n_519), .Y(n_669) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_528), .Y(n_518) );
NOR2x1_ASAP7_75t_SL g554 ( .A(n_519), .B(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g572 ( .A(n_519), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g585 ( .A(n_519), .B(n_529), .Y(n_585) );
BUFx2_ASAP7_75t_L g604 ( .A(n_519), .Y(n_604) );
INVx2_ASAP7_75t_SL g631 ( .A(n_519), .Y(n_631) );
OR2x6_ASAP7_75t_L g519 ( .A(n_520), .B(n_527), .Y(n_519) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g541 ( .A(n_529), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g687 ( .A(n_529), .B(n_629), .Y(n_687) );
INVx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_532), .B(n_538), .Y(n_530) );
AO21x1_ASAP7_75t_SL g555 ( .A1(n_531), .A2(n_532), .B(n_538), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_537), .Y(n_532) );
AOI211xp5_ASAP7_75t_L g703 ( .A1(n_540), .A2(n_564), .B(n_704), .C(n_708), .Y(n_703) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_541), .B(n_619), .Y(n_654) );
BUFx2_ASAP7_75t_L g618 ( .A(n_542), .Y(n_618) );
OR2x2_ASAP7_75t_L g566 ( .A(n_543), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g651 ( .A(n_543), .B(n_585), .Y(n_651) );
AND2x2_ASAP7_75t_L g672 ( .A(n_543), .B(n_628), .Y(n_672) );
INVx2_ASAP7_75t_L g679 ( .A(n_543), .Y(n_679) );
OAI21xp5_ASAP7_75t_SL g684 ( .A1(n_544), .A2(n_685), .B(n_686), .Y(n_684) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_547), .Y(n_544) );
AND2x2_ASAP7_75t_L g626 ( .A(n_545), .B(n_608), .Y(n_626) );
OR2x2_ASAP7_75t_L g705 ( .A(n_545), .B(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_546), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_548), .Y(n_579) );
AND2x2_ASAP7_75t_L g656 ( .A(n_548), .B(n_603), .Y(n_656) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_553), .Y(n_550) );
AND2x2_ASAP7_75t_L g641 ( .A(n_551), .B(n_642), .Y(n_641) );
AND2x4_ASAP7_75t_SL g650 ( .A(n_551), .B(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_551), .B(n_560), .Y(n_683) );
INVx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g559 ( .A(n_552), .B(n_560), .Y(n_559) );
OR2x2_ASAP7_75t_L g678 ( .A(n_553), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g628 ( .A(n_554), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g598 ( .A(n_555), .B(n_573), .Y(n_598) );
OAI31xp33_ASAP7_75t_L g605 ( .A1(n_556), .A2(n_606), .A3(n_608), .B(n_610), .Y(n_605) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_558), .B(n_581), .Y(n_607) );
AO21x1_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_565), .B(n_569), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
OR2x2_ASAP7_75t_L g617 ( .A(n_563), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g722 ( .A(n_563), .Y(n_722) );
INVx2_ASAP7_75t_SL g707 ( .A(n_564), .Y(n_707) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g611 ( .A(n_567), .B(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g695 ( .A(n_567), .B(n_696), .Y(n_695) );
INVx2_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_568), .B(n_631), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_576), .B1(n_580), .B2(n_582), .Y(n_569) );
AOI21xp33_ASAP7_75t_L g688 ( .A1(n_570), .A2(n_689), .B(n_690), .Y(n_688) );
INVx3_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
INVx1_ASAP7_75t_L g629 ( .A(n_573), .Y(n_629) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g643 ( .A(n_575), .B(n_604), .Y(n_643) );
OR2x2_ASAP7_75t_L g668 ( .A(n_575), .B(n_669), .Y(n_668) );
OR2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_577), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_577), .B(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g667 ( .A(n_577), .Y(n_667) );
INVx2_ASAP7_75t_L g596 ( .A(n_578), .Y(n_596) );
INVx1_ASAP7_75t_L g676 ( .A(n_579), .Y(n_676) );
AND2x2_ASAP7_75t_L g599 ( .A(n_581), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g673 ( .A(n_581), .Y(n_673) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_587), .B(n_605), .Y(n_586) );
OAI321xp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_592), .A3(n_597), .B1(n_598), .B2(n_599), .C(n_604), .Y(n_587) );
AOI322xp5_ASAP7_75t_L g713 ( .A1(n_588), .A2(n_619), .A3(n_714), .B1(n_716), .B2(n_718), .C1(n_719), .C2(n_724), .Y(n_713) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
BUFx2_ASAP7_75t_L g666 ( .A(n_591), .Y(n_666) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_596), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_593), .B(n_673), .Y(n_690) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g698 ( .A(n_596), .Y(n_698) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp33_ASAP7_75t_SL g630 ( .A(n_598), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OAI21xp33_ASAP7_75t_SL g697 ( .A1(n_601), .A2(n_607), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx3_ASAP7_75t_L g619 ( .A(n_612), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_633), .Y(n_613) );
AOI221xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_619), .B1(n_620), .B2(n_621), .C(n_624), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_616), .Y(n_635) );
AND2x2_ASAP7_75t_L g620 ( .A(n_618), .B(n_619), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OAI22xp33_ASAP7_75t_SL g624 ( .A1(n_625), .A2(n_627), .B1(n_630), .B2(n_632), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g636 ( .A(n_628), .B(n_637), .Y(n_636) );
OAI21xp33_ASAP7_75t_L g719 ( .A1(n_631), .A2(n_720), .B(n_721), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NOR3xp33_ASAP7_75t_SL g638 ( .A(n_639), .B(n_670), .C(n_691), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_643), .A2(n_678), .B1(n_705), .B2(n_707), .Y(n_704) );
OAI21xp33_ASAP7_75t_SL g644 ( .A1(n_645), .A2(n_646), .B(n_650), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_645), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_651), .A2(n_693), .B1(n_694), .B2(n_697), .C(n_699), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_655), .B1(n_657), .B2(n_659), .C(n_660), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g689 ( .A(n_655), .Y(n_689) );
INVx1_ASAP7_75t_L g711 ( .A(n_656), .Y(n_711) );
INVx1_ASAP7_75t_SL g709 ( .A(n_657), .Y(n_709) );
AOI31xp33_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_662), .A3(n_664), .B(n_668), .Y(n_660) );
OAI221xp5_ASAP7_75t_L g670 ( .A1(n_661), .A2(n_671), .B1(n_673), .B2(n_674), .C(n_757), .Y(n_670) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_667), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI211xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_677), .B(n_680), .C(n_688), .Y(n_674) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g686 ( .A(n_679), .B(n_687), .Y(n_686) );
OAI21xp5_ASAP7_75t_SL g680 ( .A1(n_681), .A2(n_683), .B(n_684), .Y(n_680) );
INVx1_ASAP7_75t_L g715 ( .A(n_687), .Y(n_715) );
BUFx2_ASAP7_75t_SL g724 ( .A(n_687), .Y(n_724) );
NAND3xp33_ASAP7_75t_SL g691 ( .A(n_692), .B(n_703), .C(n_713), .Y(n_691) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AOI21xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B(n_702), .Y(n_699) );
AOI21xp33_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_710), .B(n_712), .Y(n_708) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVxp67_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
CKINVDCx11_ASAP7_75t_R g726 ( .A(n_727), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_732), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_732), .B(n_750), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_734), .Y(n_733) );
BUFx3_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NOR2x1_ASAP7_75t_R g750 ( .A(n_735), .B(n_751), .Y(n_750) );
INVx3_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g746 ( .A(n_742), .Y(n_746) );
INVx2_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
endmodule