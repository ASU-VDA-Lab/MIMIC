module fake_jpeg_31018_n_535 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_535);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_535;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_54),
.Y(n_151)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_55),
.Y(n_152)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

HAxp5_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_0),
.CON(n_57),
.SN(n_57)
);

NAND2x1_ASAP7_75t_L g136 ( 
.A(n_57),
.B(n_38),
.Y(n_136)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_58),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_60),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_23),
.B(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_68),
.Y(n_106)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_23),
.B(n_17),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_69),
.Y(n_158)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_72),
.Y(n_163)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_24),
.B(n_17),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_75),
.B(n_102),
.Y(n_125)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_80),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_81),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_82),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_84),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g114 ( 
.A(n_89),
.Y(n_114)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_90),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_94),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

BUFx4f_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_96),
.Y(n_150)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_39),
.Y(n_100)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_24),
.B(n_18),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_105),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_45),
.Y(n_138)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_39),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_59),
.A2(n_26),
.B1(n_28),
.B2(n_43),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_120),
.A2(n_162),
.B1(n_44),
.B2(n_28),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_61),
.A2(n_33),
.B1(n_41),
.B2(n_52),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_130),
.A2(n_132),
.B1(n_164),
.B2(n_113),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_68),
.B(n_51),
.C(n_48),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_131),
.B(n_34),
.C(n_25),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_75),
.A2(n_52),
.B1(n_31),
.B2(n_32),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_138),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_25),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_149),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_91),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_143),
.A2(n_81),
.B1(n_87),
.B2(n_85),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_57),
.A2(n_45),
.B1(n_50),
.B2(n_49),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_43),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_L g146 ( 
.A1(n_96),
.A2(n_50),
.B(n_21),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_146),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_53),
.B(n_49),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_34),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_72),
.B(n_46),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_71),
.A2(n_21),
.B1(n_47),
.B2(n_26),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_74),
.A2(n_86),
.B1(n_78),
.B2(n_88),
.Y(n_164)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_168),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_167),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_169),
.Y(n_230)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_107),
.Y(n_170)
);

INVx13_ASAP7_75t_L g271 ( 
.A(n_170),
.Y(n_271)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_109),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_171),
.B(n_172),
.Y(n_234)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_173),
.B(n_180),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_114),
.A2(n_98),
.B1(n_66),
.B2(n_77),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_175),
.A2(n_212),
.B1(n_214),
.B2(n_218),
.Y(n_228)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_177),
.Y(n_272)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_178),
.Y(n_232)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_124),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_181),
.B(n_182),
.Y(n_241)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_183),
.B(n_190),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_184),
.A2(n_196),
.B1(n_207),
.B2(n_117),
.Y(n_239)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_107),
.Y(n_185)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_185),
.Y(n_244)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_187),
.B(n_209),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_118),
.A2(n_82),
.B1(n_51),
.B2(n_43),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_188),
.A2(n_193),
.B1(n_220),
.B2(n_162),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_108),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_189),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_166),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_125),
.B(n_31),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_191),
.B(n_195),
.Y(n_270)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_192),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_115),
.A2(n_26),
.B1(n_28),
.B2(n_47),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_194),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_114),
.Y(n_195)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_197),
.Y(n_268)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_150),
.Y(n_198)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_198),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_136),
.A2(n_44),
.B(n_47),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_199),
.A2(n_137),
.B(n_126),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_106),
.B(n_32),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_200),
.B(n_202),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_201),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_127),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_203),
.B(n_206),
.Y(n_275)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_150),
.Y(n_204)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_204),
.Y(n_265)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_111),
.Y(n_205)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_205),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_141),
.B(n_46),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_115),
.A2(n_44),
.B1(n_100),
.B2(n_104),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_146),
.B(n_18),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_208),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_134),
.A2(n_18),
.B1(n_16),
.B2(n_15),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_154),
.Y(n_210)
);

BUFx24_ASAP7_75t_L g254 ( 
.A(n_210),
.Y(n_254)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_110),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_211),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_166),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_160),
.B(n_151),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_213),
.Y(n_259)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_122),
.B(n_0),
.C(n_1),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_215),
.B(n_222),
.Y(n_247)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_157),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_216),
.Y(n_251)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_111),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_217),
.Y(n_267)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_121),
.Y(n_218)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_161),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_219),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_237)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_152),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_122),
.B(n_0),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_134),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_121),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_112),
.B(n_126),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_225),
.B(n_137),
.Y(n_253)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_117),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_226),
.A2(n_227),
.B1(n_128),
.B2(n_119),
.Y(n_243)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_120),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_199),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_231),
.B(n_261),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_179),
.A2(n_196),
.B1(n_220),
.B2(n_159),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_236),
.A2(n_249),
.B1(n_258),
.B2(n_9),
.Y(n_308)
);

OA22x2_ASAP7_75t_L g304 ( 
.A1(n_239),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_L g242 ( 
.A1(n_181),
.A2(n_152),
.B1(n_133),
.B2(n_119),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_242),
.A2(n_221),
.B1(n_170),
.B2(n_185),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_243),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_246),
.A2(n_239),
.B1(n_270),
.B2(n_253),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_176),
.B(n_1),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_248),
.B(n_275),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_197),
.A2(n_159),
.B1(n_113),
.B2(n_133),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_253),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_255),
.A2(n_225),
.B(n_224),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_219),
.A2(n_123),
.B1(n_116),
.B2(n_108),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_216),
.A2(n_112),
.B1(n_204),
.B2(n_198),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_260),
.A2(n_263),
.B1(n_169),
.B2(n_210),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_174),
.B(n_123),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_203),
.A2(n_128),
.B1(n_116),
.B2(n_5),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_174),
.B(n_14),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_3),
.Y(n_288)
);

OR2x4_ASAP7_75t_L g266 ( 
.A(n_187),
.B(n_3),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g276 ( 
.A1(n_266),
.A2(n_209),
.B(n_195),
.C(n_215),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_276),
.B(n_288),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_277),
.A2(n_287),
.B1(n_312),
.B2(n_256),
.Y(n_336)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_256),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_278),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_202),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_279),
.B(n_285),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_281),
.A2(n_296),
.B1(n_304),
.B2(n_308),
.Y(n_321)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_250),
.Y(n_282)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_282),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_283),
.A2(n_305),
.B1(n_311),
.B2(n_251),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_247),
.B(n_186),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_284),
.B(n_290),
.Y(n_319)
);

XNOR2x1_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_213),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_286),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_228),
.A2(n_205),
.B1(n_211),
.B2(n_214),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_178),
.C(n_177),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_168),
.C(n_192),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_291),
.B(n_300),
.Y(n_331)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_250),
.Y(n_292)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_292),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_234),
.B(n_226),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_293),
.B(n_302),
.Y(n_341)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_240),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_294),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_238),
.A2(n_189),
.B1(n_4),
.B2(n_6),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_265),
.Y(n_297)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_297),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_244),
.Y(n_298)
);

INVx5_ASAP7_75t_L g325 ( 
.A(n_298),
.Y(n_325)
);

INVx4_ASAP7_75t_SL g299 ( 
.A(n_232),
.Y(n_299)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_299),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_3),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_265),
.Y(n_301)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_301),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_235),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_230),
.Y(n_303)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_303),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_246),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_231),
.B(n_9),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_306),
.B(n_313),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_255),
.A2(n_238),
.B(n_264),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_307),
.A2(n_317),
.B(n_295),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_234),
.B(n_10),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_309),
.B(n_310),
.Y(n_342)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_256),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_241),
.A2(n_257),
.B1(n_230),
.B2(n_259),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_251),
.A2(n_11),
.B1(n_14),
.B2(n_268),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_238),
.A2(n_11),
.B1(n_14),
.B2(n_233),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_241),
.B(n_257),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_314),
.B(n_315),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_237),
.A2(n_266),
.B1(n_275),
.B2(n_235),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_316),
.B(n_244),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_230),
.A2(n_252),
.B(n_266),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_322),
.A2(n_328),
.B1(n_334),
.B2(n_339),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_323),
.A2(n_324),
.B(n_286),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_317),
.A2(n_248),
.B(n_245),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_284),
.A2(n_268),
.B1(n_262),
.B2(n_232),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_298),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_329),
.B(n_337),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_280),
.A2(n_262),
.B1(n_232),
.B2(n_245),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_336),
.A2(n_310),
.B1(n_278),
.B2(n_294),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_314),
.Y(n_337)
);

NOR2x1_ASAP7_75t_L g338 ( 
.A(n_315),
.B(n_254),
.Y(n_338)
);

OA21x2_ASAP7_75t_L g365 ( 
.A1(n_338),
.A2(n_303),
.B(n_304),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_280),
.A2(n_229),
.B1(n_272),
.B2(n_267),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_345),
.B(n_346),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_295),
.B(n_229),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_307),
.B(n_313),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_347),
.B(n_349),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_289),
.A2(n_272),
.B1(n_240),
.B2(n_269),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_348),
.A2(n_350),
.B1(n_308),
.B2(n_289),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_300),
.B(n_269),
.Y(n_349)
);

OAI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_302),
.A2(n_269),
.B1(n_240),
.B2(n_273),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_299),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_351),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_299),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_352),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_279),
.C(n_290),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_355),
.B(n_358),
.C(n_360),
.Y(n_389)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_318),
.Y(n_357)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_357),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_327),
.B(n_291),
.C(n_285),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_359),
.A2(n_365),
.B(n_344),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_319),
.B(n_306),
.C(n_276),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_343),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_361),
.B(n_362),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_351),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_318),
.Y(n_363)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_363),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_366),
.A2(n_368),
.B1(n_376),
.B2(n_381),
.Y(n_394)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_326),
.Y(n_367)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_367),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_322),
.A2(n_296),
.B1(n_304),
.B2(n_301),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_326),
.Y(n_369)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_369),
.Y(n_412)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_335),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_371),
.B(n_375),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_372),
.A2(n_378),
.B1(n_348),
.B2(n_339),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_319),
.B(n_288),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_373),
.B(n_354),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_323),
.B(n_282),
.C(n_292),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_374),
.B(n_333),
.C(n_332),
.Y(n_391)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_335),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_338),
.A2(n_304),
.B1(n_297),
.B2(n_273),
.Y(n_376)
);

BUFx8_ASAP7_75t_L g377 ( 
.A(n_343),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_377),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_321),
.A2(n_337),
.B1(n_333),
.B2(n_347),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_325),
.A2(n_254),
.B1(n_271),
.B2(n_329),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_353),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_382),
.B(n_387),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_338),
.A2(n_254),
.B1(n_271),
.B2(n_330),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_384),
.A2(n_386),
.B1(n_321),
.B2(n_352),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_341),
.B(n_254),
.Y(n_385)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_385),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_334),
.A2(n_271),
.B1(n_328),
.B2(n_320),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_353),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_346),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_388),
.B(n_340),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_383),
.B(n_341),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_390),
.B(n_398),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_391),
.B(n_392),
.C(n_393),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_355),
.B(n_331),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_358),
.B(n_331),
.C(n_320),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_360),
.B(n_332),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_397),
.B(n_399),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_347),
.C(n_324),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_400),
.B(n_402),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_376),
.A2(n_345),
.B1(n_342),
.B2(n_349),
.Y(n_401)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_401),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_368),
.A2(n_342),
.B1(n_354),
.B2(n_340),
.Y(n_403)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_403),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_359),
.B(n_373),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_405),
.B(n_409),
.Y(n_421)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_408),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_388),
.A2(n_325),
.B1(n_344),
.B2(n_365),
.Y(n_409)
);

AO21x1_ASAP7_75t_L g435 ( 
.A1(n_413),
.A2(n_417),
.B(n_363),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_380),
.B(n_385),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_414),
.B(n_415),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_380),
.B(n_370),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_364),
.A2(n_344),
.B1(n_386),
.B2(n_366),
.Y(n_416)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_416),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_384),
.A2(n_365),
.B(n_370),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_364),
.B(n_369),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_418),
.B(n_391),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_406),
.B(n_356),
.Y(n_424)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_424),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_398),
.B(n_401),
.Y(n_425)
);

MAJx2_ASAP7_75t_L g454 ( 
.A(n_425),
.B(n_393),
.C(n_389),
.Y(n_454)
);

BUFx12_ASAP7_75t_L g426 ( 
.A(n_407),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_426),
.B(n_445),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_396),
.B(n_379),
.Y(n_427)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_427),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_410),
.B(n_362),
.Y(n_428)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_428),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_435),
.A2(n_377),
.B(n_445),
.Y(n_467)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_404),
.Y(n_436)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_436),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_437),
.B(n_418),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_411),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_438),
.B(n_439),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_412),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_395),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_440),
.B(n_441),
.Y(n_451)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_415),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_419),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_443),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_409),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_414),
.B(n_362),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_444),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_403),
.B(n_367),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_392),
.C(n_389),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_447),
.B(n_425),
.C(n_423),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_438),
.A2(n_422),
.B1(n_443),
.B2(n_399),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_449),
.A2(n_450),
.B1(n_464),
.B2(n_467),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_422),
.A2(n_417),
.B1(n_413),
.B2(n_394),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_433),
.Y(n_453)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_453),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_454),
.B(n_455),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_430),
.B(n_397),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_437),
.B(n_405),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_457),
.B(n_461),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_420),
.B(n_402),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_458),
.B(n_421),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_434),
.A2(n_394),
.B1(n_416),
.B2(n_400),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_459),
.A2(n_434),
.B1(n_431),
.B2(n_436),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_421),
.B(n_371),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_463),
.B(n_420),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_433),
.A2(n_375),
.B1(n_361),
.B2(n_377),
.Y(n_464)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_467),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_468),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_469),
.B(n_472),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_448),
.B(n_426),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_470),
.B(n_481),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_452),
.A2(n_424),
.B1(n_431),
.B2(n_427),
.Y(n_473)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_473),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_457),
.B(n_429),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_474),
.B(n_477),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_446),
.A2(n_423),
.B1(n_439),
.B2(n_429),
.Y(n_476)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_476),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_478),
.B(n_465),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_447),
.B(n_444),
.C(n_432),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_455),
.C(n_461),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_446),
.Y(n_481)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_462),
.Y(n_483)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_483),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_458),
.B(n_435),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_484),
.B(n_472),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_486),
.B(n_484),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_478),
.B(n_466),
.Y(n_488)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_488),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_480),
.B(n_460),
.Y(n_489)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_489),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_479),
.B(n_426),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_491),
.B(n_495),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_468),
.B(n_440),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_497),
.B(n_471),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_474),
.B(n_469),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_498),
.B(n_499),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_500),
.B(n_502),
.Y(n_513)
);

OAI21xp33_ASAP7_75t_L g501 ( 
.A1(n_487),
.A2(n_482),
.B(n_451),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_501),
.B(n_428),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_485),
.A2(n_492),
.B1(n_490),
.B2(n_456),
.Y(n_502)
);

NOR2xp67_ASAP7_75t_L g505 ( 
.A(n_497),
.B(n_454),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_505),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_486),
.B(n_426),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_507),
.B(n_508),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_498),
.B(n_471),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_509),
.B(n_511),
.Y(n_516)
);

XNOR2x1_ASAP7_75t_L g511 ( 
.A(n_496),
.B(n_451),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_503),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_512),
.B(n_514),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_503),
.B(n_493),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_517),
.B(n_519),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_504),
.A2(n_490),
.B1(n_456),
.B2(n_435),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_513),
.B(n_510),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_520),
.A2(n_522),
.B(n_518),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_515),
.B(n_508),
.Y(n_521)
);

NOR2xp67_ASAP7_75t_SL g527 ( 
.A(n_521),
.B(n_475),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_516),
.B(n_506),
.Y(n_522)
);

OAI21xp33_ASAP7_75t_L g528 ( 
.A1(n_525),
.A2(n_526),
.B(n_524),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_523),
.A2(n_501),
.B(n_518),
.Y(n_526)
);

AOI21xp33_ASAP7_75t_L g529 ( 
.A1(n_527),
.A2(n_511),
.B(n_475),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_528),
.A2(n_529),
.B(n_521),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_530),
.Y(n_531)
);

AOI221xp5_ASAP7_75t_L g532 ( 
.A1(n_531),
.A2(n_519),
.B1(n_442),
.B2(n_459),
.C(n_441),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_532),
.A2(n_432),
.B(n_496),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_463),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_534),
.A2(n_494),
.B(n_522),
.Y(n_535)
);


endmodule