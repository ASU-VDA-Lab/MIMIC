module fake_jpeg_19188_n_161 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_161);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_161;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx11_ASAP7_75t_SL g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_8),
.Y(n_59)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_33),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_0),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_9),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_0),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_19),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_76),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_81),
.A2(n_62),
.B1(n_61),
.B2(n_56),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_88),
.A2(n_54),
.B1(n_60),
.B2(n_76),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_53),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_91),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_59),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_94),
.Y(n_102)
);

INVxp33_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_97),
.Y(n_119)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_99),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_93),
.B(n_86),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_86),
.C(n_76),
.Y(n_108)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_101),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_61),
.B1(n_54),
.B2(n_49),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_75),
.B1(n_73),
.B2(n_67),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_84),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_105),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_92),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_106),
.A2(n_69),
.B1(n_66),
.B2(n_64),
.Y(n_123)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_110),
.Y(n_132)
);

CKINVDCx12_ASAP7_75t_R g111 ( 
.A(n_98),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_71),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_116),
.Y(n_131)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_106),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_1),
.Y(n_128)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_120),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_70),
.B1(n_51),
.B2(n_52),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_121),
.A2(n_123),
.B1(n_58),
.B2(n_50),
.Y(n_124)
);

AO22x1_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_60),
.B1(n_63),
.B2(n_68),
.Y(n_122)
);

AO21x1_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_63),
.B(n_65),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_132),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_130),
.B(n_108),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_122),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_2),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_135),
.Y(n_137)
);

INVxp67_ASAP7_75t_SL g135 ( 
.A(n_117),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_3),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_136),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_138),
.A2(n_141),
.B(n_143),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_127),
.A2(n_121),
.B1(n_117),
.B2(n_109),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_139),
.A2(n_135),
.B1(n_125),
.B2(n_126),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_129),
.Y(n_141)
);

OAI32xp33_ASAP7_75t_L g143 ( 
.A1(n_131),
.A2(n_30),
.A3(n_46),
.B1(n_45),
.B2(n_44),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_134),
.C(n_137),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_147),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_28),
.C(n_43),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_148),
.Y(n_150)
);

XNOR2x2_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_146),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_150),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_140),
.C(n_144),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_27),
.Y(n_155)
);

OAI21x1_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_29),
.B(n_42),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_15),
.B1(n_40),
.B2(n_37),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_157),
.B(n_47),
.Y(n_158)
);

AOI321xp33_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_11),
.A3(n_35),
.B1(n_32),
.B2(n_12),
.C(n_36),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_4),
.C(n_5),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_5),
.B(n_6),
.Y(n_161)
);


endmodule