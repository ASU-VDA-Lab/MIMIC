module real_aes_15748_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_82;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_693;
wire n_496;
wire n_281;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_87;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
AOI22xp5_ASAP7_75t_L g243 ( .A1(n_0), .A2(n_2), .B1(n_244), .B2(n_245), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_0), .A2(n_150), .B1(n_663), .B2(n_665), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_0), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_1), .A2(n_16), .B1(n_171), .B2(n_180), .Y(n_188) );
INVx1_ASAP7_75t_L g505 ( .A(n_3), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_3), .B(n_466), .Y(n_571) );
XNOR2xp5_ASAP7_75t_L g669 ( .A(n_4), .B(n_27), .Y(n_669) );
INVx1_ASAP7_75t_L g573 ( .A(n_5), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_6), .A2(n_40), .B1(n_91), .B2(n_131), .Y(n_130) );
AOI22xp5_ASAP7_75t_L g108 ( .A1(n_7), .A2(n_10), .B1(n_109), .B2(n_110), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_8), .Y(n_179) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_9), .Y(n_93) );
INVx1_ASAP7_75t_L g520 ( .A(n_11), .Y(n_520) );
INVx1_ASAP7_75t_L g526 ( .A(n_11), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_12), .A2(n_674), .B1(n_675), .B2(n_676), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_12), .Y(n_675) );
INVx2_ASAP7_75t_L g516 ( .A(n_13), .Y(n_516) );
OAI21x1_ASAP7_75t_L g118 ( .A1(n_14), .A2(n_39), .B(n_119), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_15), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_17), .B(n_88), .Y(n_200) );
INVx4_ASAP7_75t_R g153 ( .A(n_18), .Y(n_153) );
OAI22xp33_ASAP7_75t_L g457 ( .A1(n_19), .A2(n_29), .B1(n_458), .B2(n_467), .Y(n_457) );
OAI22xp33_ASAP7_75t_L g547 ( .A1(n_19), .A2(n_29), .B1(n_548), .B2(n_551), .Y(n_547) );
INVx1_ASAP7_75t_L g488 ( .A(n_20), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_21), .B(n_171), .Y(n_206) );
INVx1_ASAP7_75t_L g249 ( .A(n_22), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_SL g177 ( .A1(n_23), .A2(n_87), .B(n_109), .C(n_178), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_24), .A2(n_36), .B1(n_109), .B2(n_113), .Y(n_189) );
INVx1_ASAP7_75t_L g674 ( .A(n_25), .Y(n_674) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_26), .Y(n_174) );
OAI22xp33_ASAP7_75t_SL g493 ( .A1(n_28), .A2(n_67), .B1(n_494), .B2(n_496), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_28), .A2(n_67), .B1(n_512), .B2(n_521), .Y(n_511) );
INVx1_ASAP7_75t_L g580 ( .A(n_30), .Y(n_580) );
INVx2_ASAP7_75t_L g560 ( .A(n_31), .Y(n_560) );
INVx1_ASAP7_75t_L g634 ( .A(n_31), .Y(n_634) );
INVx1_ASAP7_75t_L g203 ( .A(n_32), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_33), .B(n_109), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_34), .Y(n_222) );
INVx2_ASAP7_75t_L g651 ( .A(n_35), .Y(n_651) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_37), .Y(n_156) );
AOI22xp33_ASAP7_75t_L g112 ( .A1(n_38), .A2(n_66), .B1(n_109), .B2(n_113), .Y(n_112) );
BUFx3_ASAP7_75t_L g518 ( .A(n_41), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_42), .Y(n_121) );
AND2x4_ASAP7_75t_L g83 ( .A(n_43), .B(n_84), .Y(n_83) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_43), .Y(n_637) );
INVx1_ASAP7_75t_L g119 ( .A(n_44), .Y(n_119) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_45), .Y(n_463) );
OAI211xp5_ASAP7_75t_L g473 ( .A1(n_46), .A2(n_474), .B(n_479), .C(n_484), .Y(n_473) );
INVx1_ASAP7_75t_L g544 ( .A(n_46), .Y(n_544) );
INVx1_ASAP7_75t_L g492 ( .A(n_47), .Y(n_492) );
OAI211xp5_ASAP7_75t_L g527 ( .A1(n_47), .A2(n_528), .B(n_535), .C(n_539), .Y(n_527) );
INVx1_ASAP7_75t_L g575 ( .A(n_48), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_49), .A2(n_70), .B1(n_113), .B2(n_242), .Y(n_241) );
AO22x1_ASAP7_75t_L g134 ( .A1(n_50), .A2(n_58), .B1(n_135), .B2(n_137), .Y(n_134) );
INVx1_ASAP7_75t_L g84 ( .A(n_51), .Y(n_84) );
AND2x2_ASAP7_75t_L g181 ( .A(n_52), .B(n_182), .Y(n_181) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_53), .Y(n_462) );
INVx1_ASAP7_75t_L g586 ( .A(n_54), .Y(n_586) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_55), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_56), .B(n_131), .Y(n_228) );
INVx1_ASAP7_75t_L g592 ( .A(n_57), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_59), .B(n_171), .Y(n_223) );
INVx2_ASAP7_75t_L g88 ( .A(n_60), .Y(n_88) );
INVx1_ASAP7_75t_L g670 ( .A(n_61), .Y(n_670) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_62), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_63), .B(n_182), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_64), .B(n_117), .Y(n_132) );
BUFx3_ASAP7_75t_L g466 ( .A(n_65), .Y(n_466) );
INVx1_ASAP7_75t_L g470 ( .A(n_65), .Y(n_470) );
INVx1_ASAP7_75t_L g509 ( .A(n_68), .Y(n_509) );
INVx2_ASAP7_75t_L g570 ( .A(n_68), .Y(n_570) );
INVx1_ASAP7_75t_L g633 ( .A(n_68), .Y(n_633) );
XOR2xp5_ASAP7_75t_L g453 ( .A(n_69), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_71), .B(n_182), .Y(n_219) );
INVx1_ASAP7_75t_L g606 ( .A(n_72), .Y(n_606) );
A2O1A1Ixp33_ASAP7_75t_L g148 ( .A1(n_73), .A2(n_115), .B(n_131), .C(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g605 ( .A(n_74), .Y(n_605) );
AND2x2_ASAP7_75t_L g158 ( .A(n_75), .B(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g595 ( .A(n_76), .Y(n_595) );
NAND2xp33_ASAP7_75t_L g227 ( .A(n_77), .B(n_154), .Y(n_227) );
INVx1_ASAP7_75t_SL g683 ( .A(n_77), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_94), .B(n_452), .Y(n_78) );
CKINVDCx16_ASAP7_75t_R g79 ( .A(n_80), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
AND2x2_ASAP7_75t_L g81 ( .A(n_82), .B(n_85), .Y(n_81) );
AO31x2_ASAP7_75t_L g106 ( .A1(n_82), .A2(n_107), .A3(n_116), .B(n_120), .Y(n_106) );
INVx2_ASAP7_75t_L g157 ( .A(n_82), .Y(n_157) );
BUFx10_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
INVx1_ASAP7_75t_L g141 ( .A(n_83), .Y(n_141) );
BUFx10_ASAP7_75t_L g191 ( .A(n_83), .Y(n_191) );
INVx1_ASAP7_75t_L g247 ( .A(n_83), .Y(n_247) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_84), .Y(n_639) );
INVxp67_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AO21x1_ASAP7_75t_L g692 ( .A1(n_86), .A2(n_638), .B(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g86 ( .A(n_87), .B(n_89), .Y(n_86) );
INVx6_ASAP7_75t_L g111 ( .A(n_87), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_87), .B(n_134), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_87), .A2(n_227), .B(n_228), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g270 ( .A1(n_87), .A2(n_126), .B(n_134), .C(n_140), .Y(n_270) );
BUFx8_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx1_ASAP7_75t_L g115 ( .A(n_88), .Y(n_115) );
INVx2_ASAP7_75t_L g129 ( .A(n_88), .Y(n_129) );
INVx1_ASAP7_75t_L g176 ( .A(n_88), .Y(n_176) );
HB1xp67_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_92), .B(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx3_ASAP7_75t_L g109 ( .A(n_93), .Y(n_109) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_93), .Y(n_113) );
INVx1_ASAP7_75t_L g131 ( .A(n_93), .Y(n_131) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_93), .Y(n_136) );
INVx1_ASAP7_75t_L g138 ( .A(n_93), .Y(n_138) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_93), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_93), .Y(n_155) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_93), .Y(n_171) );
INVx1_ASAP7_75t_L g173 ( .A(n_93), .Y(n_173) );
INVx2_ASAP7_75t_L g180 ( .A(n_93), .Y(n_180) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
NOR2x2_ASAP7_75t_L g97 ( .A(n_98), .B(n_366), .Y(n_97) );
NAND4xp75_ASAP7_75t_L g98 ( .A(n_99), .B(n_271), .C(n_313), .D(n_337), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
OAI211xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_160), .B(n_208), .C(n_250), .Y(n_100) );
INVxp67_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
BUFx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g357 ( .A(n_103), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g451 ( .A(n_103), .B(n_388), .Y(n_451) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_123), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND2x2_ASAP7_75t_L g266 ( .A(n_105), .B(n_218), .Y(n_266) );
AND2x2_ASAP7_75t_L g307 ( .A(n_105), .B(n_268), .Y(n_307) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g214 ( .A(n_106), .B(n_143), .Y(n_214) );
OR2x2_ASAP7_75t_L g232 ( .A(n_106), .B(n_143), .Y(n_232) );
INVx2_ASAP7_75t_L g258 ( .A(n_106), .Y(n_258) );
AND2x2_ASAP7_75t_L g288 ( .A(n_106), .B(n_218), .Y(n_288) );
AND2x2_ASAP7_75t_L g317 ( .A(n_106), .B(n_142), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_106), .B(n_269), .Y(n_353) );
OAI22x1_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_111), .B1(n_112), .B2(n_114), .Y(n_107) );
INVx4_ASAP7_75t_L g110 ( .A(n_109), .Y(n_110) );
O2A1O1Ixp33_ASAP7_75t_L g221 ( .A1(n_110), .A2(n_222), .B(n_223), .C(n_224), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_111), .A2(n_127), .B1(n_188), .B2(n_189), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_111), .A2(n_114), .B1(n_241), .B2(n_243), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_113), .B(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g244 ( .A(n_113), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_114), .B(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g122 ( .A(n_117), .Y(n_122) );
OAI21xp33_ASAP7_75t_L g140 ( .A1(n_117), .A2(n_132), .B(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g146 ( .A(n_117), .Y(n_146) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_118), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
INVx2_ASAP7_75t_L g159 ( .A(n_122), .Y(n_159) );
BUFx2_ASAP7_75t_L g166 ( .A(n_122), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_122), .B(n_193), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_122), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g330 ( .A(n_123), .B(n_259), .Y(n_330) );
INVx2_ASAP7_75t_L g425 ( .A(n_123), .Y(n_425) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_142), .Y(n_123) );
INVx2_ASAP7_75t_L g213 ( .A(n_124), .Y(n_213) );
AND2x4_ASAP7_75t_L g256 ( .A(n_124), .B(n_143), .Y(n_256) );
AOI21x1_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_133), .B(n_139), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OAI21x1_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_130), .B(n_132), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_127), .A2(n_205), .B(n_206), .Y(n_204) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g225 ( .A(n_129), .Y(n_225) );
INVxp67_ASAP7_75t_SL g135 ( .A(n_136), .Y(n_135) );
OAI21xp33_ASAP7_75t_SL g199 ( .A1(n_137), .A2(n_200), .B(n_201), .Y(n_199) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_141), .A2(n_168), .B(n_177), .Y(n_167) );
AND2x2_ASAP7_75t_L g415 ( .A(n_142), .B(n_213), .Y(n_415) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g279 ( .A(n_143), .Y(n_279) );
AND2x2_ASAP7_75t_L g336 ( .A(n_143), .B(n_218), .Y(n_336) );
AND2x2_ASAP7_75t_L g351 ( .A(n_143), .B(n_259), .Y(n_351) );
AND2x2_ASAP7_75t_L g373 ( .A(n_143), .B(n_213), .Y(n_373) );
AO21x2_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_147), .B(n_158), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_151), .B(n_157), .Y(n_147) );
INVx2_ASAP7_75t_L g665 ( .A(n_150), .Y(n_665) );
OAI22xp33_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B1(n_155), .B2(n_156), .Y(n_152) );
INVx2_ASAP7_75t_L g242 ( .A(n_154), .Y(n_242) );
OAI211xp5_ASAP7_75t_SL g420 ( .A1(n_160), .A2(n_421), .B(n_423), .C(n_430), .Y(n_420) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_194), .Y(n_161) );
INVxp67_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
OR2x2_ASAP7_75t_L g407 ( .A(n_163), .B(n_343), .Y(n_407) );
OR2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_184), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_164), .B(n_196), .Y(n_306) );
INVxp67_ASAP7_75t_L g320 ( .A(n_164), .Y(n_320) );
AND2x2_ASAP7_75t_L g340 ( .A(n_164), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_164), .B(n_253), .Y(n_347) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g236 ( .A(n_165), .Y(n_236) );
AOI21x1_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_181), .Y(n_165) );
AO31x2_ASAP7_75t_L g239 ( .A1(n_166), .A2(n_240), .A3(n_246), .B(n_248), .Y(n_239) );
OAI21xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_172), .B(n_175), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
INVx2_ASAP7_75t_L g245 ( .A(n_173), .Y(n_245) );
BUFx4f_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_176), .B(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
INVx2_ASAP7_75t_L g190 ( .A(n_182), .Y(n_190) );
NOR2x1_ASAP7_75t_L g229 ( .A(n_182), .B(n_230), .Y(n_229) );
INVx4_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g207 ( .A(n_183), .B(n_191), .Y(n_207) );
OR2x2_ASAP7_75t_L g281 ( .A(n_184), .B(n_263), .Y(n_281) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
OR2x2_ASAP7_75t_L g329 ( .A(n_185), .B(n_236), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_185), .B(n_239), .Y(n_335) );
INVx2_ASAP7_75t_SL g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g235 ( .A(n_186), .B(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g304 ( .A(n_186), .B(n_239), .Y(n_304) );
BUFx2_ASAP7_75t_L g311 ( .A(n_186), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_186), .B(n_239), .Y(n_391) );
AO31x2_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_190), .A3(n_191), .B(n_192), .Y(n_186) );
INVx1_ASAP7_75t_L g230 ( .A(n_191), .Y(n_230) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x4_ASAP7_75t_L g321 ( .A(n_195), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g450 ( .A(n_195), .B(n_235), .Y(n_450) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx3_ASAP7_75t_L g253 ( .A(n_196), .Y(n_253) );
AND2x2_ASAP7_75t_L g264 ( .A(n_196), .B(n_239), .Y(n_264) );
AND2x2_ASAP7_75t_L g310 ( .A(n_196), .B(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g343 ( .A(n_196), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_196), .B(n_254), .Y(n_360) );
AND2x2_ASAP7_75t_L g399 ( .A(n_196), .B(n_400), .Y(n_399) );
AND2x4_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
OAI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_204), .B(n_207), .Y(n_198) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_215), .B(n_233), .Y(n_208) );
INVx2_ASAP7_75t_SL g209 ( .A(n_210), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_210), .A2(n_378), .B1(n_379), .B2(n_381), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_211), .B(n_214), .Y(n_210) );
AND2x2_ASAP7_75t_L g375 ( .A(n_211), .B(n_266), .Y(n_375) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g290 ( .A(n_212), .Y(n_290) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g439 ( .A(n_213), .B(n_259), .Y(n_439) );
AND2x2_ASAP7_75t_L g403 ( .A(n_214), .B(n_298), .Y(n_403) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_231), .Y(n_215) );
OR2x2_ASAP7_75t_L g300 ( .A(n_216), .B(n_277), .Y(n_300) );
OR2x2_ASAP7_75t_L g412 ( .A(n_216), .B(n_232), .Y(n_412) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g275 ( .A(n_217), .Y(n_275) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g259 ( .A(n_218), .Y(n_259) );
BUFx3_ASAP7_75t_L g341 ( .A(n_218), .Y(n_341) );
NAND2x1p5_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
OAI21x1_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_226), .B(n_229), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g689 ( .A(n_222), .Y(n_689) );
INVx2_ASAP7_75t_SL g224 ( .A(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g409 ( .A(n_232), .B(n_268), .Y(n_409) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_237), .Y(n_234) );
AND2x2_ASAP7_75t_L g251 ( .A(n_235), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g292 ( .A(n_235), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g429 ( .A(n_235), .Y(n_429) );
INVx1_ASAP7_75t_L g448 ( .A(n_235), .Y(n_448) );
INVx2_ASAP7_75t_L g263 ( .A(n_236), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_236), .B(n_239), .Y(n_312) );
INVx1_ASAP7_75t_L g376 ( .A(n_237), .Y(n_376) );
BUFx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g437 ( .A(n_238), .Y(n_437) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g254 ( .A(n_239), .Y(n_254) );
INVx1_ASAP7_75t_L g344 ( .A(n_239), .Y(n_344) );
INVx2_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_255), .B1(n_260), .B2(n_265), .Y(n_250) );
AND2x4_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
INVx2_ASAP7_75t_L g293 ( .A(n_253), .Y(n_293) );
AND2x2_ASAP7_75t_L g295 ( .A(n_253), .B(n_280), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_253), .B(n_263), .Y(n_355) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx3_ASAP7_75t_L g286 ( .A(n_256), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_256), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g380 ( .A(n_256), .B(n_364), .Y(n_380) );
INVx1_ASAP7_75t_L g284 ( .A(n_257), .Y(n_284) );
AOI222xp33_ASAP7_75t_L g294 ( .A1(n_257), .A2(n_295), .B1(n_296), .B2(n_301), .C1(n_307), .C2(n_308), .Y(n_294) );
OAI21xp33_ASAP7_75t_SL g324 ( .A1(n_257), .A2(n_325), .B(n_326), .Y(n_324) );
AND2x2_ASAP7_75t_L g348 ( .A(n_257), .B(n_267), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_257), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
OR2x2_ASAP7_75t_L g277 ( .A(n_258), .B(n_269), .Y(n_277) );
INVx1_ASAP7_75t_L g365 ( .A(n_258), .Y(n_365) );
BUFx2_ASAP7_75t_L g299 ( .A(n_259), .Y(n_299) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_264), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_262), .B(n_303), .Y(n_332) );
OR2x2_ASAP7_75t_L g444 ( .A(n_262), .B(n_304), .Y(n_444) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g327 ( .A(n_264), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g442 ( .A(n_264), .Y(n_442) );
OAI31xp33_ASAP7_75t_L g423 ( .A1(n_265), .A2(n_424), .A3(n_426), .B(n_427), .Y(n_423) );
AND2x4_ASAP7_75t_SL g265 ( .A(n_266), .B(n_267), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_266), .B(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_294), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_280), .B(n_282), .Y(n_272) );
NOR2x1_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x6_ASAP7_75t_L g393 ( .A(n_275), .B(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx1_ASAP7_75t_L g325 ( .A(n_278), .Y(n_325) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g416 ( .A(n_279), .B(n_353), .Y(n_416) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_281), .A2(n_370), .B1(n_372), .B2(n_374), .Y(n_369) );
A2O1A1Ixp33_ASAP7_75t_L g430 ( .A1(n_281), .A2(n_342), .B(n_404), .C(n_431), .Y(n_430) );
AOI21xp33_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_287), .B(n_291), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND4xp25_ASAP7_75t_L g383 ( .A(n_286), .B(n_384), .C(n_385), .D(n_387), .Y(n_383) );
NAND2x1_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_288), .B(n_290), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_288), .B(n_373), .Y(n_396) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g362 ( .A(n_293), .B(n_322), .Y(n_362) );
NAND2xp33_ASAP7_75t_L g296 ( .A(n_297), .B(n_300), .Y(n_296) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_300), .A2(n_444), .B1(n_445), .B2(n_447), .Y(n_443) );
AOI221x1_ASAP7_75t_L g382 ( .A1(n_301), .A2(n_383), .B1(n_389), .B2(n_392), .C(n_395), .Y(n_382) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g322 ( .A(n_304), .Y(n_322) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g334 ( .A(n_306), .B(n_335), .Y(n_334) );
NAND2x1p5_ASAP7_75t_L g397 ( .A(n_307), .B(n_388), .Y(n_397) );
O2A1O1Ixp5_ASAP7_75t_L g410 ( .A1(n_308), .A2(n_392), .B(n_411), .C(n_413), .Y(n_410) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx2_ASAP7_75t_L g359 ( .A(n_311), .Y(n_359) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_323), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_318), .Y(n_314) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_315), .A2(n_333), .B1(n_403), .B2(n_404), .C(n_406), .Y(n_402) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g339 ( .A(n_317), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_317), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g438 ( .A(n_317), .B(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
INVxp67_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
NAND2x1_ASAP7_75t_L g417 ( .A(n_320), .B(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g441 ( .A(n_320), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g381 ( .A(n_321), .Y(n_381) );
AOI222xp33_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_327), .B1(n_330), .B2(n_331), .C1(n_333), .C2(n_336), .Y(n_323) );
INVx1_ASAP7_75t_L g408 ( .A(n_327), .Y(n_408) );
INVx1_ASAP7_75t_L g371 ( .A(n_328), .Y(n_371) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g405 ( .A(n_329), .Y(n_405) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g346 ( .A(n_335), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g400 ( .A(n_335), .Y(n_400) );
AND2x2_ASAP7_75t_L g363 ( .A(n_336), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_356), .Y(n_337) );
AOI222xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_342), .B1(n_345), .B2(n_348), .C1(n_349), .C2(n_354), .Y(n_338) );
INVx3_ASAP7_75t_L g388 ( .A(n_341), .Y(n_388) );
BUFx2_ASAP7_75t_L g446 ( .A(n_341), .Y(n_446) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g418 ( .A(n_343), .Y(n_418) );
OR2x2_ASAP7_75t_L g428 ( .A(n_343), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
INVx2_ASAP7_75t_SL g386 ( .A(n_351), .Y(n_386) );
AND2x2_ASAP7_75t_L g431 ( .A(n_352), .B(n_388), .Y(n_431) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_353), .Y(n_384) );
INVxp67_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g390 ( .A(n_355), .B(n_391), .Y(n_390) );
NOR2x1_ASAP7_75t_L g356 ( .A(n_357), .B(n_361), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
OR2x2_ASAP7_75t_L g447 ( .A(n_360), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx1_ASAP7_75t_L g378 ( .A(n_362), .Y(n_378) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g385 ( .A(n_365), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g435 ( .A(n_365), .Y(n_435) );
NAND4xp75_ASAP7_75t_L g366 ( .A(n_367), .B(n_401), .C(n_419), .D(n_432), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_382), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_376), .B(n_377), .Y(n_368) );
INVxp33_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_371), .B(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g394 ( .A(n_373), .Y(n_394) );
AND2x2_ASAP7_75t_L g434 ( .A(n_373), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g404 ( .A(n_376), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g422 ( .A(n_387), .Y(n_422) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OAI22xp33_ASAP7_75t_SL g413 ( .A1(n_390), .A2(n_414), .B1(n_416), .B2(n_417), .Y(n_413) );
INVx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI21xp33_ASAP7_75t_SL g395 ( .A1(n_396), .A2(n_397), .B(n_398), .Y(n_395) );
INVx1_ASAP7_75t_L g426 ( .A(n_397), .Y(n_426) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_410), .Y(n_401) );
AOI21xp5_ASAP7_75t_SL g406 ( .A1(n_407), .A2(n_408), .B(n_409), .Y(n_406) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_449), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_436), .B1(n_438), .B2(n_440), .C(n_443), .Y(n_433) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
OAI221xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_636), .B1(n_640), .B2(n_684), .C(n_685), .Y(n_452) );
INVx1_ASAP7_75t_L g684 ( .A(n_454), .Y(n_684) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_510), .C(n_564), .Y(n_455) );
OAI31xp33_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_473), .A3(n_493), .B(n_502), .Y(n_456) );
OR2x6_ASAP7_75t_L g458 ( .A(n_459), .B(n_464), .Y(n_458) );
OR2x6_ASAP7_75t_L g495 ( .A(n_459), .B(n_469), .Y(n_495) );
BUFx4f_ASAP7_75t_L g574 ( .A(n_459), .Y(n_574) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx4f_ASAP7_75t_L g604 ( .A(n_460), .Y(n_604) );
INVx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
AND2x2_ASAP7_75t_L g471 ( .A(n_462), .B(n_472), .Y(n_471) );
NAND2x1_ASAP7_75t_L g478 ( .A(n_462), .B(n_463), .Y(n_478) );
AND2x2_ASAP7_75t_L g483 ( .A(n_462), .B(n_463), .Y(n_483) );
INVx1_ASAP7_75t_L g491 ( .A(n_462), .Y(n_491) );
INVx2_ASAP7_75t_L g501 ( .A(n_462), .Y(n_501) );
INVx2_ASAP7_75t_L g585 ( .A(n_462), .Y(n_585) );
INVx2_ASAP7_75t_L g472 ( .A(n_463), .Y(n_472) );
BUFx2_ASAP7_75t_L g487 ( .A(n_463), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_463), .B(n_501), .Y(n_500) );
OR2x2_ASAP7_75t_L g584 ( .A(n_463), .B(n_585), .Y(n_584) );
INVxp67_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g481 ( .A(n_465), .Y(n_481) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx2_ASAP7_75t_L g486 ( .A(n_466), .Y(n_486) );
AND2x4_ASAP7_75t_L g489 ( .A(n_466), .B(n_490), .Y(n_489) );
AND2x4_ASAP7_75t_L g598 ( .A(n_466), .B(n_505), .Y(n_598) );
CKINVDCx16_ASAP7_75t_R g467 ( .A(n_468), .Y(n_467) );
AND2x4_ASAP7_75t_L g468 ( .A(n_469), .B(n_471), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_SL g588 ( .A(n_477), .Y(n_588) );
BUFx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_478), .Y(n_594) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_488), .B1(n_489), .B2(n_492), .Y(n_484) );
AND2x4_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
OR2x2_ASAP7_75t_L g498 ( .A(n_486), .B(n_499), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_488), .A2(n_540), .B1(n_544), .B2(n_545), .Y(n_539) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx8_ASAP7_75t_L g578 ( .A(n_499), .Y(n_578) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx2_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
BUFx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g563 ( .A(n_508), .Y(n_563) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OAI31xp33_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_527), .A3(n_547), .B(n_557), .Y(n_510) );
BUFx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OR2x4_ASAP7_75t_L g513 ( .A(n_514), .B(n_517), .Y(n_513) );
AND2x4_ASAP7_75t_L g552 ( .A(n_514), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OR2x6_ASAP7_75t_L g523 ( .A(n_515), .B(n_524), .Y(n_523) );
AND2x4_ASAP7_75t_L g536 ( .A(n_515), .B(n_537), .Y(n_536) );
OR2x4_ASAP7_75t_L g550 ( .A(n_515), .B(n_517), .Y(n_550) );
NAND3x1_ASAP7_75t_L g631 ( .A(n_515), .B(n_632), .C(n_634), .Y(n_631) );
AND2x4_ASAP7_75t_L g649 ( .A(n_515), .B(n_650), .Y(n_649) );
INVx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx3_ASAP7_75t_L g542 ( .A(n_516), .Y(n_542) );
NAND2xp33_ASAP7_75t_SL g610 ( .A(n_516), .B(n_560), .Y(n_610) );
INVx2_ASAP7_75t_L g614 ( .A(n_517), .Y(n_614) );
OR2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_518), .B(n_526), .Y(n_525) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_518), .Y(n_534) );
AND2x4_ASAP7_75t_L g537 ( .A(n_518), .B(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g556 ( .A(n_518), .Y(n_556) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVxp67_ASAP7_75t_L g555 ( .A(n_520), .Y(n_555) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g623 ( .A(n_524), .Y(n_623) );
BUFx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g628 ( .A(n_525), .Y(n_628) );
INVx1_ASAP7_75t_L g533 ( .A(n_526), .Y(n_533) );
INVx2_ASAP7_75t_L g538 ( .A(n_526), .Y(n_538) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
OAI22xp33_ASAP7_75t_L g635 ( .A1(n_529), .A2(n_575), .B1(n_595), .B2(n_612), .Y(n_635) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx4_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx2_ASAP7_75t_L g617 ( .A(n_532), .Y(n_617) );
NAND2x1p5_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
BUFx2_ASAP7_75t_L g546 ( .A(n_533), .Y(n_546) );
BUFx2_ASAP7_75t_L g543 ( .A(n_534), .Y(n_543) );
INVx2_ASAP7_75t_L g648 ( .A(n_534), .Y(n_648) );
CKINVDCx8_ASAP7_75t_R g535 ( .A(n_536), .Y(n_535) );
AND2x4_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
AND2x4_ASAP7_75t_L g545 ( .A(n_541), .B(n_546), .Y(n_545) );
INVx3_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx6f_ASAP7_75t_L g620 ( .A(n_554), .Y(n_620) );
AND2x4_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_561), .Y(n_557) );
INVx1_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g650 ( .A(n_560), .Y(n_650) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g600 ( .A(n_563), .Y(n_600) );
OR2x2_ASAP7_75t_L g609 ( .A(n_563), .B(n_610), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_607), .Y(n_564) );
OAI33xp33_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_572), .A3(n_579), .B1(n_589), .B2(n_596), .B3(n_601), .Y(n_565) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x4_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
BUFx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OAI22xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_574), .B1(n_575), .B2(n_576), .Y(n_572) );
OAI22xp33_ASAP7_75t_L g611 ( .A1(n_573), .A2(n_592), .B1(n_612), .B2(n_615), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_576), .A2(n_602), .B1(n_605), .B2(n_606), .Y(n_601) );
INVx5_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_581), .B1(n_586), .B2(n_587), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_580), .A2(n_605), .B1(n_619), .B2(n_621), .Y(n_618) );
INVx4_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx4_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
BUFx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
BUFx3_ASAP7_75t_L g591 ( .A(n_584), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_586), .A2(n_606), .B1(n_625), .B2(n_626), .Y(n_624) );
INVx5_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OAI22xp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_592), .B1(n_593), .B2(n_595), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
BUFx4f_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g596 ( .A(n_597), .Y(n_596) );
AND2x4_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OAI33xp33_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_611), .A3(n_618), .B1(n_624), .B2(n_629), .B3(n_635), .Y(n_607) );
BUFx4f_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
BUFx2_ASAP7_75t_L g656 ( .A(n_610), .Y(n_656) );
BUFx4f_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
INVx3_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
INVx5_ASAP7_75t_L g625 ( .A(n_620), .Y(n_625) );
INVx3_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
BUFx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
CKINVDCx8_ASAP7_75t_R g626 ( .A(n_627), .Y(n_626) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_630), .Y(n_629) );
INVx3_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
INVx1_ASAP7_75t_L g658 ( .A(n_637), .Y(n_658) );
BUFx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_639), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g693 ( .A(n_639), .B(n_658), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_659), .B1(n_678), .B2(n_682), .Y(n_640) );
INVx3_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
BUFx12f_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
BUFx3_ASAP7_75t_L g687 ( .A(n_643), .Y(n_687) );
BUFx8_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI211xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_651), .B(n_652), .C(n_657), .Y(n_644) );
AND2x2_ASAP7_75t_L g681 ( .A(n_645), .B(n_652), .Y(n_681) );
INVx4_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x6_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .Y(n_646) );
NAND3xp33_ASAP7_75t_L g652 ( .A(n_647), .B(n_653), .C(n_656), .Y(n_652) );
INVx3_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx3_ASAP7_75t_L g655 ( .A(n_651), .Y(n_655) );
INVx2_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
BUFx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g680 ( .A(n_657), .Y(n_680) );
OAI22xp33_ASAP7_75t_L g686 ( .A1(n_659), .A2(n_682), .B1(n_687), .B2(n_688), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_661), .B1(n_673), .B2(n_677), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_666), .B1(n_667), .B2(n_672), .Y(n_661) );
INVx1_ASAP7_75t_L g672 ( .A(n_662), .Y(n_672) );
BUFx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B1(n_670), .B2(n_671), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_670), .Y(n_671) );
INVx1_ASAP7_75t_L g677 ( .A(n_673), .Y(n_677) );
INVx1_ASAP7_75t_L g676 ( .A(n_674), .Y(n_676) );
INVx2_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
BUFx2_ASAP7_75t_L g688 ( .A(n_679), .Y(n_688) );
OR2x6_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_684), .A2(n_686), .B1(n_689), .B2(n_690), .Y(n_685) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
endmodule