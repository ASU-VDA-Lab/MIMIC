module fake_jpeg_17261_n_360 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_360);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_360;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_31),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_21),
.B(n_10),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_21),
.B(n_10),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_60),
.Y(n_89)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_57),
.Y(n_72)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

BUFx2_ASAP7_75t_R g64 ( 
.A(n_60),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_64),
.B(n_70),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_41),
.B1(n_33),
.B2(n_38),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_20),
.B1(n_26),
.B2(n_31),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_44),
.B(n_43),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_55),
.A2(n_33),
.B1(n_41),
.B2(n_42),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_71),
.A2(n_83),
.B1(n_88),
.B2(n_26),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_78),
.B(n_31),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_81),
.Y(n_93)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_32),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_49),
.A2(n_33),
.B1(n_43),
.B2(n_42),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_85),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_33),
.B1(n_38),
.B2(n_30),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_91),
.A2(n_98),
.B1(n_106),
.B2(n_110),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_62),
.B(n_78),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_87),
.Y(n_144)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_65),
.A2(n_59),
.B1(n_58),
.B2(n_46),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_40),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_101),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_40),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_28),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_111),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_105),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_20),
.B1(n_37),
.B2(n_26),
.Y(n_106)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_40),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_71),
.A2(n_37),
.B1(n_39),
.B2(n_35),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_115),
.B1(n_30),
.B2(n_28),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_118),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_86),
.A2(n_37),
.B1(n_30),
.B2(n_28),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_40),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_116),
.B(n_87),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_35),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_121),
.Y(n_132)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_120),
.Y(n_151)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_124),
.B(n_137),
.Y(n_159)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

BUFx24_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_136),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_95),
.B1(n_98),
.B2(n_109),
.Y(n_154)
);

CKINVDCx12_ASAP7_75t_R g136 ( 
.A(n_121),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_99),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_72),
.Y(n_138)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_105),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_142),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_23),
.Y(n_141)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_104),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_147),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_152),
.Y(n_161)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_94),
.B(n_27),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_148),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_94),
.B(n_27),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_94),
.B(n_24),
.Y(n_150)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_100),
.B(n_75),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_101),
.A2(n_24),
.B(n_34),
.C(n_36),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_39),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_154),
.A2(n_120),
.B1(n_81),
.B2(n_76),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_122),
.A2(n_110),
.B1(n_113),
.B2(n_116),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_169),
.B1(n_173),
.B2(n_130),
.Y(n_178)
);

AO22x1_ASAP7_75t_SL g167 ( 
.A1(n_143),
.A2(n_111),
.B1(n_97),
.B2(n_90),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_137),
.B1(n_126),
.B2(n_112),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_168),
.A2(n_152),
.B(n_142),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_145),
.A2(n_84),
.B1(n_75),
.B2(n_92),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_128),
.A2(n_82),
.B1(n_102),
.B2(n_107),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_92),
.C(n_85),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_144),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_177),
.B(n_183),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_194),
.B1(n_197),
.B2(n_198),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_158),
.A2(n_144),
.B1(n_129),
.B2(n_127),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_179),
.A2(n_180),
.B(n_184),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_158),
.A2(n_138),
.B(n_150),
.Y(n_180)
);

BUFx12_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_134),
.Y(n_200)
);

OA22x2_ASAP7_75t_L g182 ( 
.A1(n_167),
.A2(n_174),
.B1(n_171),
.B2(n_155),
.Y(n_182)
);

OA21x2_ASAP7_75t_L g220 ( 
.A1(n_182),
.A2(n_77),
.B(n_97),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_160),
.A2(n_129),
.B(n_146),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_185),
.A2(n_186),
.B1(n_188),
.B2(n_193),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_175),
.A2(n_126),
.B1(n_130),
.B2(n_141),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_139),
.B1(n_140),
.B2(n_93),
.Y(n_188)
);

NOR2xp67_ASAP7_75t_R g189 ( 
.A(n_176),
.B(n_149),
.Y(n_189)
);

NOR2x1_ASAP7_75t_R g225 ( 
.A(n_189),
.B(n_180),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_148),
.Y(n_191)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_172),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_192),
.B(n_187),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_157),
.A2(n_139),
.B1(n_93),
.B2(n_112),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_132),
.B1(n_147),
.B2(n_153),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

OAI32xp33_ASAP7_75t_L g196 ( 
.A1(n_161),
.A2(n_165),
.A3(n_166),
.B1(n_124),
.B2(n_169),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_196),
.A2(n_176),
.B(n_163),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_166),
.A2(n_132),
.B1(n_147),
.B2(n_119),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_202),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_192),
.A2(n_171),
.B1(n_163),
.B2(n_165),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_205),
.A2(n_220),
.B1(n_223),
.B2(n_195),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_189),
.B(n_159),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_212),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_188),
.B(n_185),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_209),
.A2(n_214),
.B(n_216),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_210),
.B(n_36),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_156),
.Y(n_211)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_211),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_187),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_178),
.A2(n_164),
.B(n_162),
.Y(n_214)
);

MAJx2_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_177),
.C(n_191),
.Y(n_215)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_34),
.C(n_22),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_193),
.A2(n_182),
.B(n_179),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_219),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_190),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_199),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_222),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_184),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_182),
.A2(n_164),
.B1(n_123),
.B2(n_125),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_197),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_224),
.A2(n_226),
.B1(n_77),
.B2(n_131),
.Y(n_240)
);

AO21x1_ASAP7_75t_L g233 ( 
.A1(n_225),
.A2(n_97),
.B(n_36),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_179),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_186),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_231),
.C(n_234),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_228),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_224),
.A2(n_182),
.B1(n_198),
.B2(n_181),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_229),
.A2(n_230),
.B1(n_245),
.B2(n_226),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_222),
.A2(n_182),
.B1(n_181),
.B2(n_9),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_136),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_233),
.B(n_235),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_181),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_162),
.C(n_133),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_181),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_238),
.B(n_239),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_215),
.C(n_201),
.Y(n_239)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_243),
.Y(n_271)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_201),
.B(n_209),
.C(n_204),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_204),
.B(n_131),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_250),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_225),
.B(n_22),
.Y(n_246)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_246),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_212),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_223),
.Y(n_252)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_252),
.Y(n_258)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_260),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_220),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_252),
.A2(n_251),
.B1(n_216),
.B2(n_243),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_261),
.A2(n_262),
.B1(n_263),
.B2(n_264),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_237),
.A2(n_203),
.B1(n_214),
.B2(n_220),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_241),
.A2(n_203),
.B1(n_220),
.B2(n_221),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_235),
.A2(n_217),
.B1(n_207),
.B2(n_219),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_238),
.A2(n_208),
.B(n_207),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_SL g291 ( 
.A1(n_265),
.A2(n_269),
.B(n_1),
.C(n_2),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_249),
.A2(n_206),
.B1(n_125),
.B2(n_123),
.Y(n_266)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_266),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_232),
.A2(n_206),
.B1(n_162),
.B2(n_125),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_234),
.A2(n_123),
.B1(n_133),
.B2(n_39),
.Y(n_272)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_272),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_239),
.A2(n_131),
.B1(n_80),
.B2(n_76),
.Y(n_273)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_274),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_292),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_227),
.C(n_244),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_282),
.C(n_286),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g281 ( 
.A(n_266),
.Y(n_281)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_281),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_231),
.C(n_236),
.Y(n_282)
);

NOR3xp33_ASAP7_75t_SL g283 ( 
.A(n_256),
.B(n_233),
.C(n_242),
.Y(n_283)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_283),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_246),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_290),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_250),
.C(n_245),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_80),
.C(n_22),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_57),
.C(n_32),
.Y(n_308)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_12),
.C(n_16),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_291),
.A2(n_255),
.B1(n_260),
.B2(n_253),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_259),
.A2(n_12),
.B(n_19),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_264),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_281),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_295),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_306),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_276),
.A2(n_258),
.B(n_263),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_301),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_300),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_277),
.A2(n_261),
.B(n_262),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_279),
.A2(n_257),
.B1(n_267),
.B2(n_273),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_303),
.A2(n_286),
.B1(n_291),
.B2(n_282),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_284),
.A2(n_267),
.B1(n_12),
.B2(n_13),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_304),
.A2(n_305),
.B1(n_290),
.B2(n_15),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_288),
.A2(n_11),
.B1(n_18),
.B2(n_17),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_57),
.C(n_2),
.Y(n_322)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_309),
.Y(n_311)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_311),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_280),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_294),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_314),
.B(n_315),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_299),
.A2(n_278),
.B1(n_291),
.B2(n_283),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_317),
.C(n_319),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_285),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_309),
.A2(n_291),
.B1(n_8),
.B2(n_13),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_7),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_322),
.C(n_297),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_307),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_308),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_324),
.B(n_326),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_321),
.A2(n_301),
.B(n_298),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_325),
.A2(n_5),
.B(n_15),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_300),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_327),
.B(n_313),
.Y(n_337)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_318),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_329),
.B(n_14),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_332),
.B(n_333),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_321),
.A2(n_302),
.B1(n_8),
.B2(n_13),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_310),
.A2(n_302),
.B1(n_6),
.B2(n_14),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_334),
.B(n_320),
.C(n_322),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_331),
.B(n_310),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_337),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_338),
.B(n_341),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_339),
.A2(n_17),
.B(n_2),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_328),
.B(n_5),
.C(n_15),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_340),
.B(n_342),
.C(n_330),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_5),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_342),
.B(n_324),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_343),
.A2(n_336),
.B(n_335),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_344),
.B(n_345),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_348),
.B(n_326),
.Y(n_351)
);

OAI21xp33_ASAP7_75t_L g350 ( 
.A1(n_349),
.A2(n_17),
.B(n_2),
.Y(n_350)
);

NOR3xp33_ASAP7_75t_SL g354 ( 
.A(n_350),
.B(n_1),
.C(n_3),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_351),
.B(n_345),
.C(n_346),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_353),
.A2(n_354),
.B(n_352),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_355),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_356),
.A2(n_347),
.B(n_327),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_357),
.A2(n_1),
.B(n_4),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_358),
.B(n_4),
.C(n_345),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_359),
.B(n_4),
.Y(n_360)
);


endmodule