module real_aes_3454_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_374;
wire n_379;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_L g240 ( .A(n_0), .B(n_241), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_1), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g149 ( .A1(n_2), .A2(n_8), .B1(n_150), .B2(n_153), .Y(n_149) );
O2A1O1Ixp33_ASAP7_75t_SL g306 ( .A1(n_3), .A2(n_277), .B(n_307), .C(n_308), .Y(n_306) );
OAI22xp33_ASAP7_75t_L g251 ( .A1(n_4), .A2(n_61), .B1(n_248), .B2(n_252), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_5), .A2(n_29), .B1(n_193), .B2(n_196), .Y(n_192) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_6), .Y(n_83) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_7), .A2(n_158), .B(n_161), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_9), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g173 ( .A1(n_10), .A2(n_56), .B1(n_174), .B2(n_176), .Y(n_173) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_11), .A2(n_53), .B1(n_252), .B2(n_264), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_12), .Y(n_296) );
INVx1_ASAP7_75t_L g120 ( .A(n_13), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_13), .B(n_55), .Y(n_169) );
INVxp67_ASAP7_75t_L g184 ( .A(n_13), .Y(n_184) );
INVx1_ASAP7_75t_L g89 ( .A(n_14), .Y(n_89) );
AOI22xp5_ASAP7_75t_L g342 ( .A1(n_15), .A2(n_46), .B1(n_228), .B2(n_248), .Y(n_342) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_16), .A2(n_52), .B(n_244), .Y(n_243) );
OA21x2_ASAP7_75t_L g293 ( .A1(n_16), .A2(n_52), .B(n_244), .Y(n_293) );
NAND2xp5_ASAP7_75t_SL g116 ( .A(n_17), .B(n_105), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_18), .Y(n_372) );
BUFx3_ASAP7_75t_L g205 ( .A(n_19), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g312 ( .A1(n_20), .A2(n_227), .B(n_253), .C(n_313), .Y(n_312) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_20), .Y(n_641) );
OAI22xp33_ASAP7_75t_SL g247 ( .A1(n_21), .A2(n_33), .B1(n_248), .B2(n_249), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_22), .A2(n_26), .B1(n_249), .B2(n_260), .Y(n_259) );
BUFx6f_ASAP7_75t_L g105 ( .A(n_23), .Y(n_105) );
O2A1O1Ixp5_ASAP7_75t_L g323 ( .A1(n_24), .A2(n_277), .B(n_324), .C(n_326), .Y(n_323) );
INVx1_ASAP7_75t_L g106 ( .A(n_25), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_25), .B(n_54), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_27), .B(n_271), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_28), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g141 ( .A1(n_30), .A2(n_48), .B1(n_142), .B2(n_146), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_31), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_32), .A2(n_68), .B1(n_124), .B2(n_132), .Y(n_123) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_34), .A2(n_62), .B1(n_187), .B2(n_189), .Y(n_186) );
INVx1_ASAP7_75t_L g244 ( .A(n_35), .Y(n_244) );
INVx1_ASAP7_75t_L g162 ( .A(n_36), .Y(n_162) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_37), .Y(n_216) );
AND2x4_ASAP7_75t_L g220 ( .A(n_37), .B(n_214), .Y(n_220) );
AND2x4_ASAP7_75t_L g317 ( .A(n_37), .B(n_214), .Y(n_317) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_38), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_39), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_40), .Y(n_333) );
INVx2_ASAP7_75t_L g301 ( .A(n_41), .Y(n_301) );
O2A1O1Ixp33_ASAP7_75t_L g373 ( .A1(n_42), .A2(n_277), .B(n_374), .C(n_375), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_43), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_44), .B(n_285), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_45), .A2(n_59), .B1(n_263), .B2(n_265), .Y(n_262) );
OA22x2_ASAP7_75t_L g110 ( .A1(n_47), .A2(n_55), .B1(n_105), .B2(n_109), .Y(n_110) );
INVx1_ASAP7_75t_L g138 ( .A(n_47), .Y(n_138) );
HB1xp67_ASAP7_75t_L g84 ( .A(n_49), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_50), .Y(n_283) );
NAND2xp33_ASAP7_75t_R g346 ( .A(n_51), .B(n_293), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_51), .A2(n_76), .B1(n_271), .B2(n_403), .Y(n_402) );
HB1xp67_ASAP7_75t_L g93 ( .A(n_53), .Y(n_93) );
INVx1_ASAP7_75t_L g122 ( .A(n_54), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_54), .B(n_136), .Y(n_172) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_54), .Y(n_208) );
OAI21xp33_ASAP7_75t_L g139 ( .A1(n_55), .A2(n_60), .B(n_140), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_57), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_58), .Y(n_297) );
INVx1_ASAP7_75t_L g108 ( .A(n_60), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_60), .B(n_72), .Y(n_170) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_63), .Y(n_229) );
BUFx5_ASAP7_75t_L g248 ( .A(n_63), .Y(n_248) );
INVx1_ASAP7_75t_L g261 ( .A(n_63), .Y(n_261) );
INVx2_ASAP7_75t_L g319 ( .A(n_64), .Y(n_319) );
XNOR2xp5_ASAP7_75t_L g633 ( .A(n_65), .B(n_199), .Y(n_633) );
INVx2_ASAP7_75t_L g378 ( .A(n_66), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_67), .Y(n_314) );
INVx2_ASAP7_75t_SL g214 ( .A(n_69), .Y(n_214) );
INVx1_ASAP7_75t_L g331 ( .A(n_70), .Y(n_331) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_71), .Y(n_88) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_72), .B(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g97 ( .A(n_73), .B(n_98), .Y(n_97) );
INVx2_ASAP7_75t_L g336 ( .A(n_74), .Y(n_336) );
OAI21xp33_ASAP7_75t_SL g370 ( .A1(n_75), .A2(n_248), .B(n_371), .Y(n_370) );
INVxp67_ASAP7_75t_SL g303 ( .A(n_76), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_76), .B(n_271), .Y(n_352) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_200), .B1(n_217), .B2(n_230), .C(n_627), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_92), .Y(n_78) );
OAI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_81), .B1(n_86), .B2(n_87), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
OAI22xp5_ASAP7_75t_L g81 ( .A1(n_82), .A2(n_83), .B1(n_84), .B2(n_85), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_83), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_84), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_87), .Y(n_86) );
AOI22xp5_ASAP7_75t_L g87 ( .A1(n_88), .A2(n_89), .B1(n_90), .B2(n_91), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_88), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_89), .Y(n_90) );
AOI22xp5_ASAP7_75t_L g92 ( .A1(n_93), .A2(n_94), .B1(n_198), .B2(n_199), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_93), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_94), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_94), .A2(n_199), .B1(n_629), .B2(n_630), .Y(n_628) );
HB1xp67_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
NOR2x1_ASAP7_75t_L g95 ( .A(n_96), .B(n_155), .Y(n_95) );
NAND4xp25_ASAP7_75t_L g96 ( .A(n_97), .B(n_123), .C(n_141), .D(n_149), .Y(n_96) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
BUFx6f_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
AND2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_111), .Y(n_101) );
AND2x2_ASAP7_75t_L g175 ( .A(n_102), .B(n_152), .Y(n_175) );
AND2x2_ASAP7_75t_L g188 ( .A(n_102), .B(n_144), .Y(n_188) );
AND2x4_ASAP7_75t_L g190 ( .A(n_102), .B(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_110), .Y(n_102) );
INVx1_ASAP7_75t_L g127 ( .A(n_103), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
NAND2xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
INVx2_ASAP7_75t_L g109 ( .A(n_105), .Y(n_109) );
INVx3_ASAP7_75t_L g115 ( .A(n_105), .Y(n_115) );
NAND2xp33_ASAP7_75t_L g121 ( .A(n_105), .B(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g140 ( .A(n_105), .Y(n_140) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_105), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_106), .B(n_138), .Y(n_137) );
INVxp67_ASAP7_75t_L g209 ( .A(n_106), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
OAI21xp5_ASAP7_75t_L g183 ( .A1(n_108), .A2(n_140), .B(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g128 ( .A(n_110), .Y(n_128) );
AND2x2_ASAP7_75t_L g160 ( .A(n_110), .B(n_127), .Y(n_160) );
AND2x2_ASAP7_75t_L g182 ( .A(n_110), .B(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g154 ( .A(n_111), .B(n_126), .Y(n_154) );
AND2x4_ASAP7_75t_L g195 ( .A(n_111), .B(n_160), .Y(n_195) );
AND2x4_ASAP7_75t_L g197 ( .A(n_111), .B(n_134), .Y(n_197) );
AND2x4_ASAP7_75t_L g111 ( .A(n_112), .B(n_117), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OR2x2_ASAP7_75t_L g130 ( .A(n_113), .B(n_131), .Y(n_130) );
AND2x4_ASAP7_75t_L g144 ( .A(n_113), .B(n_145), .Y(n_144) );
AND2x4_ASAP7_75t_L g152 ( .A(n_113), .B(n_117), .Y(n_152) );
AND2x2_ASAP7_75t_L g179 ( .A(n_113), .B(n_180), .Y(n_179) );
AND2x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_116), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_115), .B(n_120), .Y(n_119) );
INVxp67_ASAP7_75t_L g136 ( .A(n_115), .Y(n_136) );
NAND3xp33_ASAP7_75t_L g171 ( .A(n_116), .B(n_135), .C(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g131 ( .A(n_118), .Y(n_131) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_121), .Y(n_118) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_129), .Y(n_125) );
AND2x4_ASAP7_75t_L g143 ( .A(n_126), .B(n_144), .Y(n_143) );
AND2x4_ASAP7_75t_L g151 ( .A(n_126), .B(n_152), .Y(n_151) );
AND2x4_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
AND2x4_ASAP7_75t_L g133 ( .A(n_129), .B(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g191 ( .A(n_130), .Y(n_191) );
INVx1_ASAP7_75t_L g145 ( .A(n_131), .Y(n_145) );
BUFx12f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g148 ( .A(n_134), .B(n_144), .Y(n_148) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_139), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_138), .Y(n_210) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx4_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx8_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x4_ASAP7_75t_L g159 ( .A(n_152), .B(n_160), .Y(n_159) );
BUFx5_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
OR2x2_ASAP7_75t_L g155 ( .A(n_156), .B(n_185), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_157), .B(n_173), .Y(n_156) );
BUFx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
INVx4_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AO21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_168), .B(n_171), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_167), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
BUFx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx5_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_179), .B(n_182), .Y(n_178) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_181), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_192), .Y(n_185) );
BUFx8_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_SL g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
BUFx3_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_203), .B(n_211), .Y(n_202) );
INVxp67_ASAP7_75t_SL g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g632 ( .A(n_204), .B(n_211), .Y(n_632) );
AOI211xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_207), .C(n_210), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_212), .B(n_215), .Y(n_211) );
OR2x2_ASAP7_75t_L g635 ( .A(n_212), .B(n_216), .Y(n_635) );
INVx1_ASAP7_75t_L g638 ( .A(n_212), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_212), .B(n_215), .Y(n_639) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
BUFx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_221), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_219), .B(n_291), .Y(n_290) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_220), .B(n_242), .Y(n_254) );
OAI221xp5_ASAP7_75t_L g276 ( .A1(n_220), .A2(n_253), .B1(n_277), .B2(n_278), .C(n_281), .Y(n_276) );
INVx1_ASAP7_75t_L g345 ( .A(n_220), .Y(n_345) );
OA21x2_ASAP7_75t_L g637 ( .A1(n_221), .A2(n_638), .B(n_639), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_222), .B(n_226), .Y(n_221) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx4_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
OA22x2_ASAP7_75t_L g258 ( .A1(n_224), .A2(n_259), .B1(n_262), .B2(n_266), .Y(n_258) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_225), .B(n_247), .Y(n_246) );
INVx3_ASAP7_75t_L g253 ( .A(n_225), .Y(n_253) );
INVx1_ASAP7_75t_L g266 ( .A(n_225), .Y(n_266) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_225), .Y(n_277) );
INVx4_ASAP7_75t_L g298 ( .A(n_225), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_225), .B(n_331), .Y(n_330) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_228), .A2(n_248), .B1(n_282), .B2(n_283), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_228), .A2(n_260), .B1(n_300), .B2(n_301), .Y(n_299) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx6_ASAP7_75t_L g249 ( .A(n_229), .Y(n_249) );
INVx2_ASAP7_75t_L g252 ( .A(n_229), .Y(n_252) );
INVx3_ASAP7_75t_L g325 ( .A(n_229), .Y(n_325) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
OR2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_518), .Y(n_233) );
NAND4xp25_ASAP7_75t_L g234 ( .A(n_235), .B(n_415), .C(n_455), .D(n_489), .Y(n_234) );
AOI211xp5_ASAP7_75t_SL g235 ( .A1(n_236), .A2(n_287), .B(n_347), .C(n_406), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_255), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_237), .A2(n_392), .B1(n_502), .B2(n_504), .Y(n_501) );
BUFx3_ASAP7_75t_L g515 ( .A(n_237), .Y(n_515) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g364 ( .A(n_238), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_238), .B(n_419), .Y(n_445) );
AND2x4_ASAP7_75t_L g487 ( .A(n_238), .B(n_409), .Y(n_487) );
INVx3_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g392 ( .A(n_239), .Y(n_392) );
AND2x2_ASAP7_75t_L g412 ( .A(n_239), .B(n_409), .Y(n_412) );
INVx2_ASAP7_75t_L g430 ( .A(n_239), .Y(n_430) );
AND2x2_ASAP7_75t_L g440 ( .A(n_239), .B(n_365), .Y(n_440) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_239), .Y(n_472) );
NAND2xp33_ASAP7_75t_R g568 ( .A(n_239), .B(n_365), .Y(n_568) );
AND2x4_ASAP7_75t_L g239 ( .A(n_240), .B(n_245), .Y(n_239) );
INVx2_ASAP7_75t_L g275 ( .A(n_241), .Y(n_275) );
NOR2xp33_ASAP7_75t_SL g315 ( .A(n_241), .B(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g271 ( .A(n_242), .Y(n_271) );
NOR2xp33_ASAP7_75t_SL g318 ( .A(n_242), .B(n_319), .Y(n_318) );
INVx4_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
BUFx3_ASAP7_75t_L g268 ( .A(n_243), .Y(n_268) );
INVx2_ASAP7_75t_L g286 ( .A(n_243), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_250), .Y(n_245) );
AOI22xp33_ASAP7_75t_SL g278 ( .A1(n_248), .A2(n_249), .B1(n_279), .B2(n_280), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_248), .A2(n_249), .B1(n_296), .B2(n_297), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_248), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_248), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_SL g371 ( .A(n_248), .B(n_372), .Y(n_371) );
INVx2_ASAP7_75t_SL g265 ( .A(n_249), .Y(n_265) );
INVx2_ASAP7_75t_L g309 ( .A(n_249), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_253), .B(n_254), .Y(n_250) );
INVx2_ASAP7_75t_L g469 ( .A(n_255), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_255), .A2(n_592), .B1(n_593), .B2(n_594), .Y(n_591) );
AND2x2_ASAP7_75t_L g623 ( .A(n_255), .B(n_624), .Y(n_623) );
AND2x4_ASAP7_75t_L g255 ( .A(n_256), .B(n_272), .Y(n_255) );
OR2x2_ASAP7_75t_L g439 ( .A(n_256), .B(n_409), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_267), .B(n_269), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OAI21x1_ASAP7_75t_L g381 ( .A1(n_258), .A2(n_270), .B(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_260), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g375 ( .A(n_260), .B(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g264 ( .A(n_261), .Y(n_264) );
INVx1_ASAP7_75t_L g307 ( .A(n_263), .Y(n_307) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g429 ( .A(n_272), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_273), .B(n_365), .Y(n_393) );
INVx2_ASAP7_75t_L g474 ( .A(n_273), .Y(n_474) );
OA21x2_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_276), .B(n_284), .Y(n_273) );
OA21x2_ASAP7_75t_L g409 ( .A1(n_274), .A2(n_276), .B(n_284), .Y(n_409) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g302 ( .A(n_275), .B(n_303), .Y(n_302) );
OAI22xp33_ASAP7_75t_L g294 ( .A1(n_277), .A2(n_295), .B1(n_298), .B2(n_299), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_277), .A2(n_298), .B1(n_342), .B2(n_343), .Y(n_341) );
INVx1_ASAP7_75t_L g358 ( .A(n_277), .Y(n_358) );
NOR2xp67_ASAP7_75t_L g344 ( .A(n_285), .B(n_345), .Y(n_344) );
INVx3_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
BUFx3_ASAP7_75t_L g334 ( .A(n_286), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_286), .B(n_378), .Y(n_377) );
AND2x4_ASAP7_75t_L g287 ( .A(n_288), .B(n_320), .Y(n_287) );
AND2x2_ASAP7_75t_L g414 ( .A(n_288), .B(n_359), .Y(n_414) );
INVx2_ASAP7_75t_SL g422 ( .A(n_288), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_288), .A2(n_424), .B1(n_431), .B2(n_436), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_288), .B(n_320), .Y(n_442) );
AND2x2_ASAP7_75t_L g498 ( .A(n_288), .B(n_493), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_288), .B(n_385), .Y(n_618) );
AND2x4_ASAP7_75t_L g288 ( .A(n_289), .B(n_304), .Y(n_288) );
INVx1_ASAP7_75t_L g506 ( .A(n_289), .Y(n_506) );
AND2x2_ASAP7_75t_L g583 ( .A(n_289), .B(n_339), .Y(n_583) );
OAI21x1_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_294), .B(n_302), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_291), .B(n_317), .Y(n_382) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
BUFx3_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g337 ( .A(n_293), .Y(n_337) );
INVx1_ASAP7_75t_L g368 ( .A(n_293), .Y(n_368) );
INVx2_ASAP7_75t_L g404 ( .A(n_293), .Y(n_404) );
INVx1_ASAP7_75t_L g356 ( .A(n_295), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_298), .A2(n_329), .B1(n_330), .B2(n_332), .Y(n_328) );
INVx2_ASAP7_75t_L g355 ( .A(n_298), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_299), .Y(n_357) );
AND2x2_ASAP7_75t_L g350 ( .A(n_304), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g388 ( .A(n_304), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_304), .B(n_321), .Y(n_405) );
INVx2_ASAP7_75t_L g435 ( .A(n_304), .Y(n_435) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_304), .Y(n_454) );
INVx1_ASAP7_75t_L g488 ( .A(n_304), .Y(n_488) );
OR2x2_ASAP7_75t_L g534 ( .A(n_304), .B(n_351), .Y(n_534) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_304), .Y(n_551) );
AO31x2_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_311), .A3(n_315), .B(n_318), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_310), .Y(n_630) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NOR3xp33_ASAP7_75t_L g322 ( .A(n_316), .B(n_323), .C(n_328), .Y(n_322) );
AOI221xp5_ASAP7_75t_L g354 ( .A1(n_316), .A2(n_355), .B1(n_356), .B2(n_357), .C(n_358), .Y(n_354) );
INVx4_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g367 ( .A(n_317), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g464 ( .A(n_320), .B(n_350), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_320), .B(n_387), .Y(n_475) );
AND2x4_ASAP7_75t_L g532 ( .A(n_320), .B(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_338), .Y(n_320) );
INVx2_ASAP7_75t_L g360 ( .A(n_321), .Y(n_360) );
AND2x2_ASAP7_75t_L g434 ( .A(n_321), .B(n_435), .Y(n_434) );
BUFx2_ASAP7_75t_R g452 ( .A(n_321), .Y(n_452) );
INVx2_ASAP7_75t_L g494 ( .A(n_321), .Y(n_494) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_321), .Y(n_511) );
AO21x2_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_334), .B(n_335), .Y(n_321) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g329 ( .A(n_325), .Y(n_329) );
INVx1_ASAP7_75t_L g374 ( .A(n_325), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g353 ( .A(n_334), .B(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g361 ( .A(n_339), .Y(n_361) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_339), .Y(n_386) );
AND2x2_ASAP7_75t_L g493 ( .A(n_339), .B(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_346), .Y(n_339) );
AND2x2_ASAP7_75t_L g401 ( .A(n_340), .B(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_344), .Y(n_340) );
OAI221xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_362), .B1(n_383), .B2(n_389), .C(n_394), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_359), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_350), .B(n_452), .Y(n_530) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_350), .Y(n_593) );
AND2x2_ASAP7_75t_L g387 ( .A(n_351), .B(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_351), .B(n_360), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_351), .B(n_541), .Y(n_606) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
AND2x2_ASAP7_75t_L g400 ( .A(n_353), .B(n_401), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g369 ( .A1(n_355), .A2(n_370), .B(n_373), .Y(n_369) );
AND2x2_ASAP7_75t_L g536 ( .A(n_359), .B(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g596 ( .A(n_359), .B(n_467), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_359), .B(n_453), .Y(n_626) );
AND2x4_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
OR2x2_ASAP7_75t_L g560 ( .A(n_360), .B(n_419), .Y(n_560) );
AND2x2_ASAP7_75t_L g481 ( .A(n_361), .B(n_435), .Y(n_481) );
INVx1_ASAP7_75t_SL g503 ( .A(n_361), .Y(n_503) );
INVx1_ASAP7_75t_L g542 ( .A(n_361), .Y(n_542) );
BUFx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_363), .B(n_485), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_379), .Y(n_363) );
INVx2_ASAP7_75t_L g396 ( .A(n_364), .Y(n_396) );
INVx2_ASAP7_75t_L g419 ( .A(n_365), .Y(n_419) );
INVx2_ASAP7_75t_L g428 ( .A(n_365), .Y(n_428) );
INVx1_ASAP7_75t_L g468 ( .A(n_365), .Y(n_468) );
AND2x2_ASAP7_75t_L g508 ( .A(n_365), .B(n_474), .Y(n_508) );
OR2x2_ASAP7_75t_L g579 ( .A(n_365), .B(n_430), .Y(n_579) );
BUFx2_ASAP7_75t_L g586 ( .A(n_365), .Y(n_586) );
INVx3_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AOI21x1_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_369), .B(n_377), .Y(n_366) );
AND2x4_ASAP7_75t_L g486 ( .A(n_379), .B(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_379), .B(n_443), .Y(n_499) );
INVx3_ASAP7_75t_L g509 ( .A(n_379), .Y(n_509) );
AND2x2_ASAP7_75t_L g543 ( .A(n_379), .B(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g620 ( .A(n_379), .B(n_440), .Y(n_620) );
INVx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g410 ( .A(n_380), .Y(n_410) );
AND2x2_ASAP7_75t_L g420 ( .A(n_380), .B(n_409), .Y(n_420) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g448 ( .A(n_381), .Y(n_448) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_384), .B(n_486), .Y(n_546) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
OR2x2_ASAP7_75t_L g421 ( .A(n_385), .B(n_422), .Y(n_421) );
NOR4xp25_ASAP7_75t_L g484 ( .A(n_385), .B(n_461), .C(n_485), .D(n_488), .Y(n_484) );
OR2x2_ASAP7_75t_L g571 ( .A(n_385), .B(n_572), .Y(n_571) );
INVx2_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
OR2x2_ASAP7_75t_L g611 ( .A(n_388), .B(n_550), .Y(n_611) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx2_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_391), .B(n_447), .Y(n_446) );
NOR2xp67_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_L g553 ( .A(n_392), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_397), .Y(n_394) );
O2A1O1Ixp33_ASAP7_75t_SL g456 ( .A1(n_395), .A2(n_457), .B(n_459), .C(n_463), .Y(n_456) );
INVx2_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g564 ( .A(n_396), .B(n_438), .Y(n_564) );
OAI21xp33_ASAP7_75t_L g574 ( .A1(n_397), .A2(n_575), .B(n_577), .Y(n_574) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_405), .Y(n_398) );
OR2x2_ASAP7_75t_L g432 ( .A(n_399), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g561 ( .A(n_399), .Y(n_561) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g517 ( .A(n_400), .B(n_494), .Y(n_517) );
INVx1_ASAP7_75t_L g550 ( .A(n_400), .Y(n_550) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g602 ( .A(n_405), .Y(n_602) );
AOI21xp33_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_411), .B(n_413), .Y(n_406) );
INVx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI32xp33_ASAP7_75t_L g441 ( .A1(n_408), .A2(n_442), .A3(n_443), .B1(n_446), .B2(n_449), .Y(n_441) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx1_ASAP7_75t_L g581 ( .A(n_411), .Y(n_581) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g544 ( .A(n_412), .B(n_428), .Y(n_544) );
OAI322xp33_ASAP7_75t_L g621 ( .A1(n_413), .A2(n_474), .A3(n_479), .B1(n_576), .B2(n_586), .C1(n_622), .C2(n_625), .Y(n_621) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_441), .Y(n_415) );
OAI21xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_421), .B(n_423), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_420), .Y(n_417) );
BUFx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g460 ( .A(n_420), .Y(n_460) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NAND2x1p5_ASAP7_75t_L g425 ( .A(n_426), .B(n_429), .Y(n_425) );
INVx2_ASAP7_75t_L g599 ( .A(n_426), .Y(n_599) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g462 ( .A(n_428), .Y(n_462) );
AND2x2_ASAP7_75t_L g567 ( .A(n_428), .B(n_448), .Y(n_567) );
AND2x2_ASAP7_75t_L g607 ( .A(n_429), .B(n_509), .Y(n_607) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g582 ( .A(n_434), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g492 ( .A(n_435), .Y(n_492) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_440), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g458 ( .A(n_439), .Y(n_458) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g479 ( .A(n_445), .B(n_448), .Y(n_479) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_448), .B(n_472), .Y(n_598) );
INVxp67_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_453), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g539 ( .A(n_454), .B(n_540), .Y(n_539) );
NOR4xp25_ASAP7_75t_L g455 ( .A(n_456), .B(n_465), .C(n_476), .D(n_484), .Y(n_455) );
INVx2_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
OAI221xp5_ASAP7_75t_L g526 ( .A1(n_460), .A2(n_527), .B1(n_528), .B2(n_531), .C(n_535), .Y(n_526) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_462), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AOI21xp33_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_470), .B(n_475), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_469), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_468), .B(n_474), .Y(n_473) );
OR2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_473), .Y(n_470) );
INVxp67_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g513 ( .A(n_474), .Y(n_513) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_480), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_481), .B(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g605 ( .A(n_481), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OR2x2_ASAP7_75t_L g572 ( .A(n_483), .B(n_492), .Y(n_572) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g522 ( .A(n_487), .B(n_509), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_487), .B(n_509), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_487), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_487), .B(n_586), .Y(n_585) );
NOR2xp67_ASAP7_75t_L g604 ( .A(n_487), .B(n_566), .Y(n_604) );
INVx1_ASAP7_75t_SL g612 ( .A(n_487), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_488), .B(n_503), .Y(n_502) );
INVx2_ASAP7_75t_SL g537 ( .A(n_488), .Y(n_537) );
INVx1_ASAP7_75t_L g594 ( .A(n_488), .Y(n_594) );
AOI211xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_495), .B(n_496), .C(n_512), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_493), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g589 ( .A(n_493), .Y(n_589) );
INVx1_ASAP7_75t_L g541 ( .A(n_494), .Y(n_541) );
OAI21xp33_ASAP7_75t_SL g496 ( .A1(n_497), .A2(n_499), .B(n_500), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NAND4xp25_ASAP7_75t_L g500 ( .A(n_501), .B(n_507), .C(n_509), .D(n_510), .Y(n_500) );
OR2x2_ASAP7_75t_L g504 ( .A(n_503), .B(n_505), .Y(n_504) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_505), .Y(n_525) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x4_ASAP7_75t_L g552 ( .A(n_508), .B(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g578 ( .A(n_509), .B(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g576 ( .A(n_510), .B(n_534), .Y(n_576) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NOR3xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .C(n_516), .Y(n_512) );
INVx1_ASAP7_75t_L g592 ( .A(n_513), .Y(n_592) );
INVxp67_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_515), .B(n_570), .Y(n_569) );
AOI21xp33_ASAP7_75t_SL g565 ( .A1(n_516), .A2(n_566), .B(n_568), .Y(n_565) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NAND3xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_554), .C(n_608), .Y(n_518) );
AOI211xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_523), .B(n_526), .C(n_545), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVxp67_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
INVxp67_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g562 ( .A(n_530), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g609 ( .A1(n_531), .A2(n_610), .B(n_612), .Y(n_609) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
OR2x2_ASAP7_75t_L g588 ( .A(n_534), .B(n_589), .Y(n_588) );
OAI21xp5_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_538), .B(n_543), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_538), .A2(n_604), .B1(n_605), .B2(n_607), .Y(n_603) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_552), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
NOR3xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_573), .C(n_590), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_569), .Y(n_555) );
AOI221xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_561), .B1(n_562), .B2(n_563), .C(n_565), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g615 ( .A(n_572), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_580), .Y(n_573) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g624 ( .A(n_579), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_582), .B1(n_584), .B2(n_587), .Y(n_580) );
AND2x4_ASAP7_75t_L g601 ( .A(n_583), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OAI221xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_595), .B1(n_597), .B2(n_600), .C(n_603), .Y(n_590) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NOR3xp33_ASAP7_75t_L g608 ( .A(n_609), .B(n_613), .C(n_621), .Y(n_608) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AOI21xp33_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_616), .B(n_619), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
BUFx3_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OAI222xp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_631), .B1(n_633), .B2(n_634), .C1(n_636), .C2(n_640), .Y(n_627) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_SL g631 ( .A(n_632), .Y(n_631) );
BUFx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
BUFx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
CKINVDCx5p33_ASAP7_75t_R g640 ( .A(n_641), .Y(n_640) );
endmodule