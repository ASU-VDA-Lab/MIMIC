module fake_netlist_1_888_n_1078 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1078);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1078;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_881;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_476;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_1012;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_769;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1024;
wire n_1016;
wire n_572;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_975;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_955;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_1011;
wire n_1025;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_844;
wire n_818;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_828;
wire n_767;
wire n_1063;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_950;
wire n_935;
wire n_460;
wire n_1046;
wire n_478;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_799;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_937;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_260;
wire n_806;
wire n_1066;
wire n_539;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_522;
wire n_264;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_924;
wire n_947;
wire n_1043;
wire n_912;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1027;
wire n_1007;
wire n_859;
wire n_1040;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_406;
wire n_395;
wire n_491;
wire n_385;
wire n_257;
wire n_992;
wire n_269;
INVx1_ASAP7_75t_L g253 ( .A(n_70), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_140), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_235), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_179), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_165), .Y(n_257) );
XNOR2xp5_ASAP7_75t_L g258 ( .A(n_201), .B(n_168), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_195), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_131), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_177), .Y(n_261) );
INVxp67_ASAP7_75t_SL g262 ( .A(n_101), .Y(n_262) );
BUFx5_ASAP7_75t_L g263 ( .A(n_215), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_143), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_220), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_141), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_226), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_216), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_155), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_229), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_223), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_125), .Y(n_272) );
BUFx6f_ASAP7_75t_L g273 ( .A(n_132), .Y(n_273) );
CKINVDCx20_ASAP7_75t_R g274 ( .A(n_72), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_37), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_159), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_63), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_14), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_14), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_66), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_40), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_76), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_37), .Y(n_283) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_180), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_19), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_114), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_54), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_120), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_227), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_244), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_203), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_171), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_138), .Y(n_293) );
CKINVDCx20_ASAP7_75t_R g294 ( .A(n_167), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_115), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_173), .Y(n_296) );
BUFx3_ASAP7_75t_L g297 ( .A(n_152), .Y(n_297) );
BUFx10_ASAP7_75t_L g298 ( .A(n_64), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_154), .Y(n_299) );
INVx2_ASAP7_75t_SL g300 ( .A(n_11), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_243), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_205), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_204), .Y(n_303) );
INVxp67_ASAP7_75t_L g304 ( .A(n_3), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_81), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_24), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_3), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_33), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_144), .Y(n_309) );
CKINVDCx14_ASAP7_75t_R g310 ( .A(n_225), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_169), .Y(n_311) );
INVx2_ASAP7_75t_SL g312 ( .A(n_98), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_27), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_51), .Y(n_314) );
CKINVDCx20_ASAP7_75t_R g315 ( .A(n_178), .Y(n_315) );
INVxp33_ASAP7_75t_SL g316 ( .A(n_157), .Y(n_316) );
CKINVDCx16_ASAP7_75t_R g317 ( .A(n_118), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_145), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_65), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_193), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_112), .Y(n_321) );
INVxp67_ASAP7_75t_L g322 ( .A(n_21), .Y(n_322) );
BUFx3_ASAP7_75t_L g323 ( .A(n_192), .Y(n_323) );
INVxp33_ASAP7_75t_L g324 ( .A(n_232), .Y(n_324) );
CKINVDCx20_ASAP7_75t_R g325 ( .A(n_133), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_122), .Y(n_326) );
INVx4_ASAP7_75t_R g327 ( .A(n_109), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_46), .Y(n_328) );
CKINVDCx20_ASAP7_75t_R g329 ( .A(n_224), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_209), .Y(n_330) );
CKINVDCx20_ASAP7_75t_R g331 ( .A(n_97), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_32), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_124), .Y(n_333) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_161), .Y(n_334) );
INVxp33_ASAP7_75t_SL g335 ( .A(n_39), .Y(n_335) );
CKINVDCx20_ASAP7_75t_R g336 ( .A(n_5), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_45), .Y(n_337) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_123), .Y(n_338) );
INVxp67_ASAP7_75t_L g339 ( .A(n_129), .Y(n_339) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_47), .Y(n_340) );
INVx3_ASAP7_75t_L g341 ( .A(n_16), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_91), .Y(n_342) );
BUFx3_ASAP7_75t_L g343 ( .A(n_32), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_90), .Y(n_344) );
BUFx2_ASAP7_75t_L g345 ( .A(n_119), .Y(n_345) );
INVxp67_ASAP7_75t_SL g346 ( .A(n_247), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_194), .Y(n_347) );
CKINVDCx20_ASAP7_75t_R g348 ( .A(n_7), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_142), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_59), .Y(n_350) );
CKINVDCx16_ASAP7_75t_R g351 ( .A(n_111), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_4), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_92), .Y(n_353) );
INVxp33_ASAP7_75t_SL g354 ( .A(n_93), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_230), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_75), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_126), .Y(n_357) );
BUFx3_ASAP7_75t_L g358 ( .A(n_51), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_245), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_181), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_162), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_82), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_234), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_134), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_238), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_40), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_153), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_151), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_218), .Y(n_369) );
BUFx3_ASAP7_75t_L g370 ( .A(n_104), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_41), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_206), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_188), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_100), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_187), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_86), .Y(n_376) );
CKINVDCx16_ASAP7_75t_R g377 ( .A(n_240), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_89), .Y(n_378) );
BUFx3_ASAP7_75t_L g379 ( .A(n_149), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_163), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_121), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_42), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_175), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_29), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_148), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_7), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_164), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_199), .B(n_25), .Y(n_388) );
INVxp33_ASAP7_75t_SL g389 ( .A(n_77), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_41), .Y(n_390) );
BUFx3_ASAP7_75t_L g391 ( .A(n_297), .Y(n_391) );
OAI22x1_ASAP7_75t_R g392 ( .A1(n_274), .A2(n_2), .B1(n_0), .B2(n_1), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_263), .Y(n_393) );
AND2x4_ASAP7_75t_L g394 ( .A(n_341), .B(n_0), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_335), .A2(n_4), .B1(n_1), .B2(n_2), .Y(n_395) );
NOR2x1_ASAP7_75t_L g396 ( .A(n_341), .B(n_5), .Y(n_396) );
AND2x6_ASAP7_75t_L g397 ( .A(n_297), .B(n_94), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_263), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_312), .B(n_6), .Y(n_399) );
AND2x4_ASAP7_75t_L g400 ( .A(n_341), .B(n_6), .Y(n_400) );
NAND2x1p5_ASAP7_75t_L g401 ( .A(n_345), .B(n_343), .Y(n_401) );
OAI22xp5_ASAP7_75t_SL g402 ( .A1(n_274), .A2(n_10), .B1(n_8), .B2(n_9), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_317), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_324), .B(n_8), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_263), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_263), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_390), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_335), .A2(n_12), .B1(n_9), .B2(n_11), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_300), .B(n_12), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_389), .A2(n_16), .B1(n_13), .B2(n_15), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_389), .A2(n_18), .B1(n_13), .B2(n_17), .Y(n_411) );
INVx2_ASAP7_75t_SL g412 ( .A(n_312), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_265), .A2(n_20), .B1(n_18), .B2(n_19), .Y(n_413) );
OAI21x1_ASAP7_75t_L g414 ( .A1(n_292), .A2(n_96), .B(n_95), .Y(n_414) );
OA21x2_ASAP7_75t_L g415 ( .A1(n_292), .A2(n_102), .B(n_99), .Y(n_415) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_273), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_277), .Y(n_417) );
AND2x6_ASAP7_75t_L g418 ( .A(n_323), .B(n_103), .Y(n_418) );
INVx3_ASAP7_75t_L g419 ( .A(n_343), .Y(n_419) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_273), .Y(n_420) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_273), .Y(n_421) );
XNOR2x2_ASAP7_75t_R g422 ( .A(n_336), .B(n_340), .Y(n_422) );
BUFx3_ASAP7_75t_L g423 ( .A(n_323), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_263), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_263), .Y(n_425) );
CKINVDCx8_ASAP7_75t_R g426 ( .A(n_351), .Y(n_426) );
BUFx3_ASAP7_75t_L g427 ( .A(n_391), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_412), .B(n_377), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_412), .B(n_300), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_416), .Y(n_430) );
INVx5_ASAP7_75t_L g431 ( .A(n_397), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_401), .B(n_254), .Y(n_432) );
AND2x6_ASAP7_75t_L g433 ( .A(n_394), .B(n_388), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_394), .A2(n_278), .B1(n_279), .B2(n_253), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_394), .A2(n_285), .B1(n_305), .B2(n_283), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_401), .B(n_267), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_393), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_426), .B(n_267), .Y(n_438) );
BUFx4f_ASAP7_75t_L g439 ( .A(n_397), .Y(n_439) );
BUFx10_ASAP7_75t_L g440 ( .A(n_394), .Y(n_440) );
INVx3_ASAP7_75t_L g441 ( .A(n_400), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_416), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_393), .Y(n_443) );
OR2x6_ASAP7_75t_L g444 ( .A(n_402), .B(n_277), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_426), .B(n_270), .Y(n_445) );
HB1xp67_ASAP7_75t_SL g446 ( .A(n_426), .Y(n_446) );
INVx5_ASAP7_75t_L g447 ( .A(n_397), .Y(n_447) );
INVx5_ASAP7_75t_L g448 ( .A(n_397), .Y(n_448) );
INVx3_ASAP7_75t_L g449 ( .A(n_400), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_404), .B(n_284), .Y(n_450) );
BUFx2_ASAP7_75t_L g451 ( .A(n_407), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_416), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_393), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_398), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_403), .B(n_339), .Y(n_455) );
NAND3xp33_ASAP7_75t_L g456 ( .A(n_404), .B(n_322), .C(n_304), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_398), .Y(n_457) );
INVx4_ASAP7_75t_L g458 ( .A(n_400), .Y(n_458) );
OR2x6_ASAP7_75t_L g459 ( .A(n_402), .B(n_282), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_400), .B(n_298), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_396), .B(n_358), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_398), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_399), .B(n_270), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_419), .B(n_298), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_409), .B(n_275), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_391), .B(n_275), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_413), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_405), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_419), .B(n_272), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_416), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_451), .B(n_409), .Y(n_471) );
INVx2_ASAP7_75t_SL g472 ( .A(n_465), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_429), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_SL g474 ( .A1(n_441), .A2(n_419), .B(n_406), .C(n_405), .Y(n_474) );
AND3x1_ASAP7_75t_SL g475 ( .A(n_444), .B(n_392), .C(n_422), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_433), .A2(n_397), .B1(n_418), .B2(n_406), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_464), .B(n_423), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_465), .B(n_423), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_439), .A2(n_414), .B(n_415), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_427), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_460), .A2(n_413), .B1(n_265), .B2(n_315), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_427), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_456), .A2(n_315), .B1(n_325), .B2(n_294), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_433), .A2(n_397), .B1(n_418), .B2(n_406), .Y(n_484) );
BUFx3_ASAP7_75t_L g485 ( .A(n_427), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_439), .B(n_272), .Y(n_486) );
INVx5_ASAP7_75t_L g487 ( .A(n_433), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_450), .B(n_286), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_429), .B(n_286), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_429), .B(n_289), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_429), .B(n_289), .Y(n_491) );
INVx2_ASAP7_75t_SL g492 ( .A(n_461), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_428), .B(n_316), .Y(n_493) );
BUFx5_ASAP7_75t_L g494 ( .A(n_440), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_466), .B(n_290), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_461), .B(n_291), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_461), .B(n_293), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_433), .A2(n_397), .B1(n_418), .B2(n_405), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_432), .B(n_395), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_441), .A2(n_424), .B(n_425), .C(n_414), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_440), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_439), .B(n_424), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_436), .B(n_298), .Y(n_503) );
O2A1O1Ixp5_ASAP7_75t_L g504 ( .A1(n_439), .A2(n_346), .B(n_262), .C(n_256), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_458), .B(n_424), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_434), .A2(n_435), .B1(n_446), .B2(n_467), .Y(n_506) );
NOR2xp33_ASAP7_75t_R g507 ( .A(n_440), .B(n_325), .Y(n_507) );
INVx8_ASAP7_75t_L g508 ( .A(n_433), .Y(n_508) );
OR2x6_ASAP7_75t_L g509 ( .A(n_444), .B(n_408), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_SL g510 ( .A1(n_441), .A2(n_449), .B(n_425), .C(n_310), .Y(n_510) );
INVx2_ASAP7_75t_SL g511 ( .A(n_440), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_458), .B(n_357), .Y(n_512) );
NOR3xp33_ASAP7_75t_L g513 ( .A(n_438), .B(n_410), .C(n_408), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_441), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_431), .B(n_357), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_431), .B(n_425), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_433), .A2(n_449), .B1(n_443), .B2(n_437), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_449), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_433), .B(n_360), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_449), .Y(n_520) );
BUFx2_ASAP7_75t_L g521 ( .A(n_444), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_463), .B(n_360), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_469), .B(n_361), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_437), .B(n_364), .Y(n_524) );
INVx3_ASAP7_75t_L g525 ( .A(n_443), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_445), .A2(n_331), .B1(n_334), .B2(n_329), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_431), .B(n_367), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_431), .B(n_255), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_431), .B(n_367), .Y(n_529) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_459), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_459), .Y(n_531) );
BUFx3_ASAP7_75t_L g532 ( .A(n_447), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_453), .A2(n_414), .B(n_417), .C(n_358), .Y(n_533) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_447), .Y(n_534) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_459), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_454), .B(n_368), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_447), .B(n_448), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_447), .B(n_375), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_455), .A2(n_459), .B1(n_331), .B2(n_334), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_457), .B(n_375), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_462), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_462), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_468), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_468), .B(n_380), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_447), .A2(n_281), .B1(n_287), .B2(n_280), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_447), .B(n_380), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_448), .B(n_257), .Y(n_547) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_448), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_448), .A2(n_418), .B1(n_417), .B2(n_314), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_473), .Y(n_550) );
OAI21xp5_ASAP7_75t_L g551 ( .A1(n_500), .A2(n_415), .B(n_448), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_472), .Y(n_552) );
AO21x1_ASAP7_75t_L g553 ( .A1(n_502), .A2(n_260), .B(n_259), .Y(n_553) );
OAI22xp5_ASAP7_75t_SL g554 ( .A1(n_509), .A2(n_348), .B1(n_340), .B2(n_411), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_505), .A2(n_448), .B(n_415), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_471), .B(n_316), .Y(n_556) );
A2O1A1Ixp33_ASAP7_75t_L g557 ( .A1(n_493), .A2(n_319), .B(n_328), .C(n_313), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_492), .B(n_281), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_525), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_481), .B(n_348), .Y(n_560) );
INVx1_ASAP7_75t_SL g561 ( .A(n_494), .Y(n_561) );
BUFx4f_ASAP7_75t_L g562 ( .A(n_508), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_543), .Y(n_563) );
O2A1O1Ixp33_ASAP7_75t_L g564 ( .A1(n_513), .A2(n_344), .B(n_352), .C(n_342), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_514), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_499), .A2(n_354), .B1(n_418), .B2(n_362), .Y(n_566) );
AO32x1_ASAP7_75t_L g567 ( .A1(n_541), .A2(n_268), .A3(n_276), .B1(n_271), .B2(n_269), .Y(n_567) );
NAND2x1p5_ASAP7_75t_L g568 ( .A(n_487), .B(n_415), .Y(n_568) );
AOI21x1_ASAP7_75t_L g569 ( .A1(n_502), .A2(n_442), .B(n_430), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_505), .A2(n_295), .B(n_288), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_478), .B(n_287), .Y(n_571) );
NAND3xp33_ASAP7_75t_L g572 ( .A(n_533), .B(n_366), .C(n_356), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_518), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_474), .A2(n_301), .B(n_296), .Y(n_574) );
O2A1O1Ixp33_ASAP7_75t_L g575 ( .A1(n_506), .A2(n_376), .B(n_378), .C(n_371), .Y(n_575) );
NAND2x1p5_ASAP7_75t_L g576 ( .A(n_487), .B(n_282), .Y(n_576) );
INVx2_ASAP7_75t_SL g577 ( .A(n_503), .Y(n_577) );
A2O1A1Ixp33_ASAP7_75t_L g578 ( .A1(n_542), .A2(n_384), .B(n_382), .C(n_307), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_474), .A2(n_303), .B(n_302), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_520), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_496), .B(n_350), .Y(n_581) );
NAND2xp33_ASAP7_75t_SL g582 ( .A(n_517), .B(n_258), .Y(n_582) );
INVx2_ASAP7_75t_SL g583 ( .A(n_489), .Y(n_583) );
NAND2x1p5_ASAP7_75t_L g584 ( .A(n_487), .B(n_306), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_497), .B(n_353), .Y(n_585) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_508), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_480), .Y(n_587) );
NOR2xp33_ASAP7_75t_R g588 ( .A(n_531), .B(n_381), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_494), .B(n_381), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_477), .A2(n_320), .B(n_318), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_517), .A2(n_306), .B1(n_308), .B2(n_307), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_490), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_482), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_509), .A2(n_308), .B1(n_333), .B2(n_321), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_491), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_488), .B(n_332), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_485), .Y(n_597) );
BUFx3_ASAP7_75t_L g598 ( .A(n_521), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_485), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_539), .A2(n_359), .B1(n_365), .B2(n_347), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_508), .A2(n_372), .B1(n_373), .B2(n_369), .Y(n_601) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_494), .B(n_261), .Y(n_602) );
INVx3_ASAP7_75t_L g603 ( .A(n_494), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_524), .B(n_337), .Y(n_604) );
BUFx12f_ASAP7_75t_L g605 ( .A(n_475), .Y(n_605) );
O2A1O1Ixp33_ASAP7_75t_L g606 ( .A1(n_530), .A2(n_385), .B(n_387), .C(n_383), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_536), .Y(n_607) );
BUFx2_ASAP7_75t_L g608 ( .A(n_526), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_476), .A2(n_309), .B1(n_326), .B2(n_311), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_535), .B(n_386), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_540), .Y(n_611) );
AND2x4_ASAP7_75t_L g612 ( .A(n_511), .B(n_418), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_544), .Y(n_613) );
BUFx2_ASAP7_75t_L g614 ( .A(n_483), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_495), .B(n_512), .Y(n_615) );
BUFx6f_ASAP7_75t_L g616 ( .A(n_534), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_476), .A2(n_330), .B1(n_374), .B2(n_355), .Y(n_617) );
AO32x2_ASAP7_75t_L g618 ( .A1(n_510), .A2(n_418), .A3(n_263), .B1(n_421), .B2(n_416), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_501), .A2(n_442), .B(n_430), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_523), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_522), .B(n_264), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_545), .Y(n_622) );
A2O1A1Ixp33_ASAP7_75t_SL g623 ( .A1(n_484), .A2(n_430), .B(n_452), .C(n_442), .Y(n_623) );
INVx3_ASAP7_75t_L g624 ( .A(n_494), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_519), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_484), .B(n_266), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_486), .A2(n_470), .B(n_452), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_504), .Y(n_628) );
O2A1O1Ixp33_ASAP7_75t_L g629 ( .A1(n_515), .A2(n_363), .B(n_379), .C(n_370), .Y(n_629) );
INVx3_ASAP7_75t_L g630 ( .A(n_532), .Y(n_630) );
NAND2x1_ASAP7_75t_L g631 ( .A(n_498), .B(n_327), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_498), .B(n_299), .Y(n_632) );
BUFx2_ASAP7_75t_L g633 ( .A(n_546), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_528), .Y(n_634) );
AND2x4_ASAP7_75t_SL g635 ( .A(n_549), .B(n_273), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_516), .A2(n_470), .B(n_349), .Y(n_636) );
AOI21x1_ASAP7_75t_L g637 ( .A1(n_528), .A2(n_547), .B(n_529), .Y(n_637) );
INVx1_ASAP7_75t_SL g638 ( .A(n_527), .Y(n_638) );
AND3x1_ASAP7_75t_SL g639 ( .A(n_549), .B(n_22), .C(n_23), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_538), .B(n_23), .Y(n_640) );
BUFx12f_ASAP7_75t_L g641 ( .A(n_534), .Y(n_641) );
BUFx6f_ASAP7_75t_L g642 ( .A(n_534), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_547), .Y(n_643) );
NOR2xp67_ASAP7_75t_L g644 ( .A(n_537), .B(n_25), .Y(n_644) );
NOR2xp33_ASAP7_75t_R g645 ( .A(n_548), .B(n_26), .Y(n_645) );
AND2x4_ASAP7_75t_L g646 ( .A(n_548), .B(n_26), .Y(n_646) );
A2O1A1Ixp33_ASAP7_75t_L g647 ( .A1(n_473), .A2(n_338), .B(n_421), .C(n_420), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_472), .B(n_27), .Y(n_648) );
AOI21xp5_ASAP7_75t_L g649 ( .A1(n_479), .A2(n_421), .B(n_420), .Y(n_649) );
BUFx2_ASAP7_75t_L g650 ( .A(n_507), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_517), .A2(n_421), .B1(n_420), .B2(n_30), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_479), .A2(n_106), .B(n_105), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_479), .A2(n_108), .B(n_107), .Y(n_653) );
CKINVDCx14_ASAP7_75t_R g654 ( .A(n_507), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_473), .Y(n_655) );
OA22x2_ASAP7_75t_L g656 ( .A1(n_509), .A2(n_28), .B1(n_29), .B2(n_30), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_473), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_472), .B(n_31), .Y(n_658) );
AO32x1_ASAP7_75t_L g659 ( .A1(n_492), .A2(n_31), .A3(n_33), .B1(n_34), .B2(n_35), .Y(n_659) );
AND2x4_ASAP7_75t_L g660 ( .A(n_583), .B(n_34), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_646), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_608), .B(n_36), .Y(n_662) );
OA21x2_ASAP7_75t_L g663 ( .A1(n_551), .A2(n_113), .B(n_110), .Y(n_663) );
OAI21x1_ASAP7_75t_L g664 ( .A1(n_551), .A2(n_117), .B(n_116), .Y(n_664) );
INVx3_ASAP7_75t_L g665 ( .A(n_641), .Y(n_665) );
AO31x2_ASAP7_75t_L g666 ( .A1(n_553), .A2(n_38), .A3(n_42), .B(n_43), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_622), .B(n_43), .Y(n_667) );
AND2x4_ASAP7_75t_L g668 ( .A(n_563), .B(n_44), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_552), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_658), .Y(n_670) );
AND2x4_ASAP7_75t_L g671 ( .A(n_592), .B(n_44), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_646), .Y(n_672) );
INVx4_ASAP7_75t_L g673 ( .A(n_562), .Y(n_673) );
INVx4_ASAP7_75t_SL g674 ( .A(n_605), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_565), .Y(n_675) );
BUFx2_ASAP7_75t_L g676 ( .A(n_588), .Y(n_676) );
CKINVDCx12_ASAP7_75t_R g677 ( .A(n_554), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_573), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_648), .Y(n_679) );
AO31x2_ASAP7_75t_L g680 ( .A1(n_609), .A2(n_48), .A3(n_49), .B(n_50), .Y(n_680) );
O2A1O1Ixp33_ASAP7_75t_SL g681 ( .A1(n_623), .A2(n_170), .B(n_251), .C(n_250), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_619), .A2(n_128), .B(n_127), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_582), .A2(n_49), .B1(n_52), .B2(n_53), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_614), .B(n_52), .Y(n_684) );
O2A1O1Ixp33_ASAP7_75t_SL g685 ( .A1(n_561), .A2(n_172), .B(n_249), .C(n_248), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_594), .A2(n_55), .B1(n_56), .B2(n_57), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_595), .B(n_57), .Y(n_687) );
INVx3_ASAP7_75t_L g688 ( .A(n_586), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_556), .B(n_58), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_611), .A2(n_135), .B(n_130), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_613), .A2(n_137), .B(n_136), .Y(n_691) );
AO31x2_ASAP7_75t_L g692 ( .A1(n_609), .A2(n_60), .A3(n_61), .B(n_62), .Y(n_692) );
AOI21xp5_ASAP7_75t_L g693 ( .A1(n_568), .A2(n_627), .B(n_626), .Y(n_693) );
O2A1O1Ixp33_ASAP7_75t_SL g694 ( .A1(n_561), .A2(n_631), .B(n_628), .C(n_647), .Y(n_694) );
OR2x2_ASAP7_75t_L g695 ( .A(n_600), .B(n_62), .Y(n_695) );
AO31x2_ASAP7_75t_L g696 ( .A1(n_617), .A2(n_63), .A3(n_64), .B(n_65), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_550), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_557), .B(n_67), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g699 ( .A1(n_625), .A2(n_183), .B(n_246), .Y(n_699) );
AO32x2_ASAP7_75t_L g700 ( .A1(n_594), .A2(n_67), .A3(n_68), .B1(n_69), .B2(n_70), .Y(n_700) );
BUFx2_ASAP7_75t_L g701 ( .A(n_598), .Y(n_701) );
AOI221x1_ASAP7_75t_L g702 ( .A1(n_572), .A2(n_71), .B1(n_72), .B2(n_73), .C(n_74), .Y(n_702) );
AND2x4_ASAP7_75t_L g703 ( .A(n_577), .B(n_73), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_639), .A2(n_78), .B1(n_79), .B2(n_80), .Y(n_704) );
A2O1A1Ixp33_ASAP7_75t_L g705 ( .A1(n_620), .A2(n_78), .B(n_79), .C(n_80), .Y(n_705) );
AO32x2_ASAP7_75t_L g706 ( .A1(n_651), .A2(n_617), .A3(n_591), .B1(n_601), .B2(n_567), .Y(n_706) );
AO31x2_ASAP7_75t_L g707 ( .A1(n_652), .A2(n_83), .A3(n_84), .B(n_85), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_655), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_610), .B(n_87), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_632), .A2(n_190), .B(n_242), .Y(n_710) );
INVxp67_ASAP7_75t_SL g711 ( .A(n_586), .Y(n_711) );
AND2x6_ASAP7_75t_L g712 ( .A(n_586), .B(n_88), .Y(n_712) );
O2A1O1Ixp33_ASAP7_75t_SL g713 ( .A1(n_578), .A2(n_191), .B(n_241), .C(n_239), .Y(n_713) );
BUFx2_ASAP7_75t_L g714 ( .A(n_650), .Y(n_714) );
NAND2x1_ASAP7_75t_L g715 ( .A(n_603), .B(n_139), .Y(n_715) );
A2O1A1Ixp33_ASAP7_75t_L g716 ( .A1(n_590), .A2(n_146), .B(n_147), .C(n_150), .Y(n_716) );
A2O1A1Ixp33_ASAP7_75t_L g717 ( .A1(n_606), .A2(n_156), .B(n_158), .C(n_160), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_656), .Y(n_718) );
AND2x4_ASAP7_75t_L g719 ( .A(n_603), .B(n_252), .Y(n_719) );
NAND2x1p5_ASAP7_75t_L g720 ( .A(n_562), .B(n_166), .Y(n_720) );
INVx5_ASAP7_75t_L g721 ( .A(n_616), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_604), .A2(n_174), .B(n_176), .Y(n_722) );
A2O1A1Ixp33_ASAP7_75t_L g723 ( .A1(n_570), .A2(n_182), .B(n_184), .C(n_185), .Y(n_723) );
INVxp67_ASAP7_75t_SL g724 ( .A(n_576), .Y(n_724) );
OAI21x1_ASAP7_75t_L g725 ( .A1(n_637), .A2(n_186), .B(n_189), .Y(n_725) );
A2O1A1Ixp33_ASAP7_75t_L g726 ( .A1(n_574), .A2(n_196), .B(n_197), .C(n_198), .Y(n_726) );
AOI21xp5_ASAP7_75t_L g727 ( .A1(n_559), .A2(n_200), .B(n_202), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g728 ( .A1(n_596), .A2(n_207), .B(n_208), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_581), .A2(n_210), .B(n_211), .Y(n_729) );
AO31x2_ASAP7_75t_L g730 ( .A1(n_579), .A2(n_212), .A3(n_213), .B(n_214), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_585), .B(n_217), .Y(n_731) );
AOI221xp5_ASAP7_75t_L g732 ( .A1(n_571), .A2(n_219), .B1(n_221), .B2(n_222), .C(n_228), .Y(n_732) );
A2O1A1Ixp33_ASAP7_75t_L g733 ( .A1(n_566), .A2(n_231), .B(n_233), .C(n_236), .Y(n_733) );
INVx1_ASAP7_75t_SL g734 ( .A(n_645), .Y(n_734) );
A2O1A1Ixp33_ASAP7_75t_L g735 ( .A1(n_657), .A2(n_237), .B(n_580), .C(n_629), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_640), .A2(n_558), .B1(n_633), .B2(n_621), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_584), .B(n_644), .Y(n_737) );
INVx1_ASAP7_75t_SL g738 ( .A(n_584), .Y(n_738) );
O2A1O1Ixp5_ASAP7_75t_SL g739 ( .A1(n_567), .A2(n_659), .B(n_602), .C(n_589), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g740 ( .A1(n_612), .A2(n_636), .B(n_634), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_624), .B(n_638), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_597), .A2(n_599), .B1(n_587), .B2(n_593), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g743 ( .A1(n_643), .A2(n_638), .B(n_630), .Y(n_743) );
AND2x4_ASAP7_75t_L g744 ( .A(n_635), .B(n_630), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_616), .B(n_642), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_567), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_618), .B(n_659), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g748 ( .A1(n_659), .A2(n_555), .B(n_615), .Y(n_748) );
A2O1A1Ixp33_ASAP7_75t_L g749 ( .A1(n_618), .A2(n_615), .B(n_607), .C(n_613), .Y(n_749) );
O2A1O1Ixp33_ASAP7_75t_L g750 ( .A1(n_557), .A2(n_564), .B(n_594), .C(n_575), .Y(n_750) );
AOI21xp5_ASAP7_75t_L g751 ( .A1(n_555), .A2(n_615), .B(n_479), .Y(n_751) );
AO21x1_ASAP7_75t_L g752 ( .A1(n_649), .A2(n_653), .B(n_652), .Y(n_752) );
OAI21x1_ASAP7_75t_L g753 ( .A1(n_649), .A2(n_551), .B(n_569), .Y(n_753) );
AND2x6_ASAP7_75t_L g754 ( .A(n_561), .B(n_586), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_552), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g756 ( .A1(n_555), .A2(n_615), .B(n_479), .Y(n_756) );
OA21x2_ASAP7_75t_L g757 ( .A1(n_551), .A2(n_533), .B(n_500), .Y(n_757) );
OAI21x1_ASAP7_75t_L g758 ( .A1(n_649), .A2(n_551), .B(n_569), .Y(n_758) );
NOR2xp33_ASAP7_75t_SL g759 ( .A(n_562), .B(n_508), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_560), .B(n_472), .Y(n_760) );
INVx2_ASAP7_75t_L g761 ( .A(n_697), .Y(n_761) );
OAI221xp5_ASAP7_75t_L g762 ( .A1(n_750), .A2(n_704), .B1(n_695), .B2(n_683), .C(n_684), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_755), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_668), .Y(n_764) );
BUFx3_ASAP7_75t_L g765 ( .A(n_665), .Y(n_765) );
AO21x2_ASAP7_75t_L g766 ( .A1(n_748), .A2(n_746), .B(n_747), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_708), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_718), .B(n_679), .Y(n_768) );
INVx2_ASAP7_75t_SL g769 ( .A(n_665), .Y(n_769) );
A2O1A1Ixp33_ASAP7_75t_L g770 ( .A1(n_704), .A2(n_709), .B(n_683), .C(n_749), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_668), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_760), .B(n_736), .Y(n_772) );
BUFx2_ASAP7_75t_SL g773 ( .A(n_712), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_689), .B(n_667), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_670), .B(n_687), .Y(n_775) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_662), .A2(n_671), .B1(n_660), .B2(n_677), .Y(n_776) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_686), .A2(n_671), .B1(n_660), .B2(n_738), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_675), .Y(n_778) );
AO31x2_ASAP7_75t_L g779 ( .A1(n_752), .A2(n_702), .A3(n_735), .B(n_693), .Y(n_779) );
INVx3_ASAP7_75t_L g780 ( .A(n_673), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_678), .Y(n_781) );
AOI21xp5_ASAP7_75t_L g782 ( .A1(n_694), .A2(n_757), .B(n_731), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_703), .B(n_686), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_661), .B(n_672), .Y(n_784) );
AND2x4_ASAP7_75t_L g785 ( .A(n_673), .B(n_724), .Y(n_785) );
OAI21xp5_ASAP7_75t_L g786 ( .A1(n_739), .A2(n_740), .B(n_757), .Y(n_786) );
INVxp67_ASAP7_75t_L g787 ( .A(n_676), .Y(n_787) );
AO21x2_ASAP7_75t_L g788 ( .A1(n_681), .A2(n_664), .B(n_743), .Y(n_788) );
AND3x2_ASAP7_75t_L g789 ( .A(n_714), .B(n_759), .C(n_674), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_698), .Y(n_790) );
BUFx2_ASAP7_75t_L g791 ( .A(n_712), .Y(n_791) );
AND2x4_ASAP7_75t_L g792 ( .A(n_674), .B(n_721), .Y(n_792) );
AOI21x1_ASAP7_75t_L g793 ( .A1(n_663), .A2(n_710), .B(n_725), .Y(n_793) );
AO31x2_ASAP7_75t_L g794 ( .A1(n_726), .A2(n_733), .A3(n_716), .B(n_717), .Y(n_794) );
AO21x2_ASAP7_75t_L g795 ( .A1(n_699), .A2(n_685), .B(n_713), .Y(n_795) );
OAI21xp5_ASAP7_75t_L g796 ( .A1(n_729), .A2(n_722), .B(n_728), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_738), .B(n_737), .Y(n_797) );
AO21x2_ASAP7_75t_L g798 ( .A1(n_741), .A2(n_682), .B(n_690), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_707), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_700), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_700), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_680), .Y(n_802) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_734), .Y(n_803) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_744), .A2(n_720), .B1(n_719), .B2(n_705), .Y(n_804) );
OR2x6_ASAP7_75t_L g805 ( .A(n_744), .B(n_719), .Y(n_805) );
OAI21x1_ASAP7_75t_L g806 ( .A1(n_715), .A2(n_745), .B(n_727), .Y(n_806) );
OA21x2_ASAP7_75t_L g807 ( .A1(n_691), .A2(n_723), .B(n_732), .Y(n_807) );
BUFx2_ASAP7_75t_L g808 ( .A(n_712), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_680), .B(n_692), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_688), .B(n_711), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_666), .Y(n_811) );
AO21x1_ASAP7_75t_SL g812 ( .A1(n_754), .A2(n_742), .B(n_759), .Y(n_812) );
AND2x2_ASAP7_75t_L g813 ( .A(n_680), .B(n_692), .Y(n_813) );
OR2x2_ASAP7_75t_L g814 ( .A(n_692), .B(n_696), .Y(n_814) );
BUFx12f_ASAP7_75t_L g815 ( .A(n_754), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_688), .B(n_721), .Y(n_816) );
INVx2_ASAP7_75t_L g817 ( .A(n_666), .Y(n_817) );
A2O1A1Ixp33_ASAP7_75t_L g818 ( .A1(n_721), .A2(n_706), .B(n_696), .C(n_666), .Y(n_818) );
OR2x6_ASAP7_75t_L g819 ( .A(n_706), .B(n_696), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_706), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_730), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_730), .A2(n_509), .B1(n_554), .B2(n_513), .Y(n_822) );
AOI22xp33_ASAP7_75t_SL g823 ( .A1(n_730), .A2(n_507), .B1(n_654), .B2(n_554), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_669), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_669), .Y(n_825) );
A2O1A1Ixp33_ASAP7_75t_L g826 ( .A1(n_750), .A2(n_718), .B(n_704), .C(n_709), .Y(n_826) );
BUFx6f_ASAP7_75t_L g827 ( .A(n_721), .Y(n_827) );
AOI21xp5_ASAP7_75t_L g828 ( .A1(n_751), .A2(n_756), .B(n_748), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_750), .B(n_592), .Y(n_829) );
OA21x2_ASAP7_75t_L g830 ( .A1(n_753), .A2(n_758), .B(n_748), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_750), .B(n_592), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_750), .B(n_592), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_750), .B(n_592), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_669), .Y(n_834) );
INVx2_ASAP7_75t_L g835 ( .A(n_697), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_750), .B(n_592), .Y(n_836) );
INVx2_ASAP7_75t_L g837 ( .A(n_697), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_750), .B(n_592), .Y(n_838) );
A2O1A1Ixp33_ASAP7_75t_L g839 ( .A1(n_750), .A2(n_718), .B(n_704), .C(n_709), .Y(n_839) );
AOI21xp5_ASAP7_75t_L g840 ( .A1(n_751), .A2(n_756), .B(n_748), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_750), .B(n_592), .Y(n_841) );
BUFx3_ASAP7_75t_L g842 ( .A(n_665), .Y(n_842) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_704), .A2(n_683), .B1(n_686), .B2(n_671), .Y(n_843) );
AOI21xp5_ASAP7_75t_L g844 ( .A1(n_751), .A2(n_756), .B(n_748), .Y(n_844) );
BUFx2_ASAP7_75t_L g845 ( .A(n_701), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_669), .Y(n_846) );
AOI21xp5_ASAP7_75t_L g847 ( .A1(n_751), .A2(n_756), .B(n_748), .Y(n_847) );
OAI22xp5_ASAP7_75t_L g848 ( .A1(n_704), .A2(n_683), .B1(n_686), .B2(n_671), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_669), .Y(n_849) );
INVx2_ASAP7_75t_SL g850 ( .A(n_665), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_669), .Y(n_851) );
AOI21xp5_ASAP7_75t_L g852 ( .A1(n_751), .A2(n_756), .B(n_748), .Y(n_852) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_704), .A2(n_683), .B1(n_686), .B2(n_671), .Y(n_853) );
AOI21xp5_ASAP7_75t_L g854 ( .A1(n_751), .A2(n_756), .B(n_748), .Y(n_854) );
AND2x4_ASAP7_75t_L g855 ( .A(n_673), .B(n_665), .Y(n_855) );
HB1xp67_ASAP7_75t_L g856 ( .A(n_701), .Y(n_856) );
OAI22x1_ASAP7_75t_L g857 ( .A1(n_686), .A2(n_481), .B1(n_704), .B2(n_683), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_802), .Y(n_858) );
OR2x2_ASAP7_75t_L g859 ( .A(n_772), .B(n_777), .Y(n_859) );
INVx3_ASAP7_75t_L g860 ( .A(n_827), .Y(n_860) );
OR2x2_ASAP7_75t_L g861 ( .A(n_772), .B(n_777), .Y(n_861) );
OR2x2_ASAP7_75t_L g862 ( .A(n_783), .B(n_797), .Y(n_862) );
AO21x2_ASAP7_75t_L g863 ( .A1(n_828), .A2(n_844), .B(n_840), .Y(n_863) );
OAI222xp33_ASAP7_75t_L g864 ( .A1(n_843), .A2(n_853), .B1(n_848), .B2(n_762), .C1(n_822), .C2(n_776), .Y(n_864) );
AO21x2_ASAP7_75t_L g865 ( .A1(n_847), .A2(n_854), .B(n_852), .Y(n_865) );
HB1xp67_ASAP7_75t_L g866 ( .A(n_845), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_761), .B(n_767), .Y(n_867) );
OR2x6_ASAP7_75t_L g868 ( .A(n_773), .B(n_791), .Y(n_868) );
HB1xp67_ASAP7_75t_L g869 ( .A(n_856), .Y(n_869) );
OR2x6_ASAP7_75t_L g870 ( .A(n_808), .B(n_805), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_835), .B(n_837), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_768), .Y(n_872) );
INVx2_ASAP7_75t_L g873 ( .A(n_766), .Y(n_873) );
INVx3_ASAP7_75t_L g874 ( .A(n_827), .Y(n_874) );
AND2x2_ASAP7_75t_L g875 ( .A(n_778), .B(n_781), .Y(n_875) );
NAND3xp33_ASAP7_75t_L g876 ( .A(n_823), .B(n_818), .C(n_770), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_768), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_799), .Y(n_878) );
OA21x2_ASAP7_75t_L g879 ( .A1(n_786), .A2(n_782), .B(n_821), .Y(n_879) );
INVx3_ASAP7_75t_L g880 ( .A(n_815), .Y(n_880) );
AND2x4_ASAP7_75t_L g881 ( .A(n_805), .B(n_797), .Y(n_881) );
INVx2_ASAP7_75t_L g882 ( .A(n_830), .Y(n_882) );
BUFx3_ASAP7_75t_L g883 ( .A(n_785), .Y(n_883) );
AND2x4_ASAP7_75t_L g884 ( .A(n_805), .B(n_806), .Y(n_884) );
AO21x2_ASAP7_75t_L g885 ( .A1(n_811), .A2(n_817), .B(n_809), .Y(n_885) );
AND2x2_ASAP7_75t_L g886 ( .A(n_790), .B(n_829), .Y(n_886) );
HB1xp67_ASAP7_75t_L g887 ( .A(n_785), .Y(n_887) );
BUFx3_ASAP7_75t_L g888 ( .A(n_855), .Y(n_888) );
OR2x2_ASAP7_75t_L g889 ( .A(n_819), .B(n_814), .Y(n_889) );
AO21x2_ASAP7_75t_L g890 ( .A1(n_813), .A2(n_793), .B(n_788), .Y(n_890) );
OR2x2_ASAP7_75t_L g891 ( .A(n_819), .B(n_829), .Y(n_891) );
AND2x2_ASAP7_75t_L g892 ( .A(n_831), .B(n_832), .Y(n_892) );
OAI211xp5_ASAP7_75t_L g893 ( .A1(n_774), .A2(n_839), .B(n_826), .C(n_803), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_800), .Y(n_894) );
AND2x2_ASAP7_75t_L g895 ( .A(n_831), .B(n_832), .Y(n_895) );
OR2x2_ASAP7_75t_L g896 ( .A(n_819), .B(n_833), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_801), .Y(n_897) );
HB1xp67_ASAP7_75t_L g898 ( .A(n_765), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_763), .Y(n_899) );
AND2x2_ASAP7_75t_L g900 ( .A(n_833), .B(n_838), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_836), .B(n_841), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_824), .Y(n_902) );
OAI22xp33_ASAP7_75t_L g903 ( .A1(n_857), .A2(n_804), .B1(n_764), .B2(n_771), .Y(n_903) );
OR2x6_ASAP7_75t_L g904 ( .A(n_836), .B(n_841), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_825), .Y(n_905) );
AO21x2_ASAP7_75t_L g906 ( .A1(n_796), .A2(n_820), .B(n_795), .Y(n_906) );
AO21x2_ASAP7_75t_L g907 ( .A1(n_798), .A2(n_775), .B(n_784), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_834), .Y(n_908) );
HB1xp67_ASAP7_75t_L g909 ( .A(n_842), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_846), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_849), .B(n_851), .Y(n_911) );
AOI21xp5_ASAP7_75t_SL g912 ( .A1(n_807), .A2(n_812), .B(n_792), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_779), .Y(n_913) );
BUFx3_ASAP7_75t_L g914 ( .A(n_855), .Y(n_914) );
HB1xp67_ASAP7_75t_L g915 ( .A(n_769), .Y(n_915) );
OA21x2_ASAP7_75t_L g916 ( .A1(n_779), .A2(n_816), .B(n_810), .Y(n_916) );
INVx2_ASAP7_75t_L g917 ( .A(n_779), .Y(n_917) );
OAI221xp5_ASAP7_75t_L g918 ( .A1(n_787), .A2(n_850), .B1(n_780), .B2(n_789), .C(n_794), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_794), .Y(n_919) );
AO21x2_ASAP7_75t_L g920 ( .A1(n_828), .A2(n_844), .B(n_840), .Y(n_920) );
NAND3xp33_ASAP7_75t_L g921 ( .A(n_823), .B(n_818), .C(n_770), .Y(n_921) );
AND2x2_ASAP7_75t_L g922 ( .A(n_761), .B(n_718), .Y(n_922) );
INVx4_ASAP7_75t_L g923 ( .A(n_868), .Y(n_923) );
OR2x2_ASAP7_75t_L g924 ( .A(n_859), .B(n_861), .Y(n_924) );
BUFx2_ASAP7_75t_L g925 ( .A(n_884), .Y(n_925) );
INVx2_ASAP7_75t_L g926 ( .A(n_882), .Y(n_926) );
AND2x2_ASAP7_75t_L g927 ( .A(n_892), .B(n_895), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_895), .B(n_900), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_900), .B(n_901), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_901), .B(n_862), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_858), .Y(n_931) );
HB1xp67_ASAP7_75t_L g932 ( .A(n_869), .Y(n_932) );
NOR2x1_ASAP7_75t_L g933 ( .A(n_918), .B(n_868), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_872), .B(n_877), .Y(n_934) );
AND2x4_ASAP7_75t_L g935 ( .A(n_884), .B(n_889), .Y(n_935) );
OR2x2_ASAP7_75t_L g936 ( .A(n_889), .B(n_891), .Y(n_936) );
OR2x6_ASAP7_75t_SL g937 ( .A(n_876), .B(n_921), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_858), .Y(n_938) );
NOR2x1_ASAP7_75t_SL g939 ( .A(n_868), .B(n_870), .Y(n_939) );
HB1xp67_ASAP7_75t_L g940 ( .A(n_866), .Y(n_940) );
AND2x2_ASAP7_75t_L g941 ( .A(n_904), .B(n_907), .Y(n_941) );
AND2x4_ASAP7_75t_L g942 ( .A(n_884), .B(n_885), .Y(n_942) );
NOR2x1_ASAP7_75t_L g943 ( .A(n_868), .B(n_883), .Y(n_943) );
INVx3_ASAP7_75t_L g944 ( .A(n_884), .Y(n_944) );
HB1xp67_ASAP7_75t_L g945 ( .A(n_916), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_907), .B(n_894), .Y(n_946) );
OR2x2_ASAP7_75t_L g947 ( .A(n_891), .B(n_896), .Y(n_947) );
AND2x2_ASAP7_75t_L g948 ( .A(n_907), .B(n_897), .Y(n_948) );
HB1xp67_ASAP7_75t_L g949 ( .A(n_916), .Y(n_949) );
BUFx3_ASAP7_75t_L g950 ( .A(n_883), .Y(n_950) );
AND2x2_ASAP7_75t_L g951 ( .A(n_897), .B(n_899), .Y(n_951) );
AND2x2_ASAP7_75t_L g952 ( .A(n_899), .B(n_902), .Y(n_952) );
AND2x2_ASAP7_75t_L g953 ( .A(n_902), .B(n_905), .Y(n_953) );
AND2x2_ASAP7_75t_L g954 ( .A(n_908), .B(n_910), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_878), .Y(n_955) );
AND2x2_ASAP7_75t_L g956 ( .A(n_867), .B(n_871), .Y(n_956) );
INVx1_ASAP7_75t_SL g957 ( .A(n_887), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_871), .B(n_886), .Y(n_958) );
NOR2xp33_ASAP7_75t_L g959 ( .A(n_898), .B(n_909), .Y(n_959) );
AOI211xp5_ASAP7_75t_L g960 ( .A1(n_864), .A2(n_903), .B(n_893), .C(n_921), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_875), .B(n_922), .Y(n_961) );
AND2x2_ASAP7_75t_L g962 ( .A(n_927), .B(n_919), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_927), .B(n_913), .Y(n_963) );
INVx1_ASAP7_75t_L g964 ( .A(n_931), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_924), .B(n_876), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_938), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_938), .Y(n_967) );
INVxp67_ASAP7_75t_L g968 ( .A(n_959), .Y(n_968) );
AND2x4_ASAP7_75t_L g969 ( .A(n_944), .B(n_873), .Y(n_969) );
INVx6_ASAP7_75t_L g970 ( .A(n_923), .Y(n_970) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_932), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_958), .B(n_917), .Y(n_972) );
OR2x2_ASAP7_75t_L g973 ( .A(n_947), .B(n_920), .Y(n_973) );
AND2x2_ASAP7_75t_L g974 ( .A(n_930), .B(n_879), .Y(n_974) );
AND2x2_ASAP7_75t_L g975 ( .A(n_951), .B(n_879), .Y(n_975) );
INVx2_ASAP7_75t_L g976 ( .A(n_926), .Y(n_976) );
AND2x2_ASAP7_75t_L g977 ( .A(n_951), .B(n_879), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_946), .B(n_879), .Y(n_978) );
BUFx3_ASAP7_75t_L g979 ( .A(n_950), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_956), .B(n_911), .Y(n_980) );
AND2x2_ASAP7_75t_L g981 ( .A(n_946), .B(n_906), .Y(n_981) );
OR2x2_ASAP7_75t_L g982 ( .A(n_947), .B(n_920), .Y(n_982) );
AND2x2_ASAP7_75t_L g983 ( .A(n_948), .B(n_906), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_952), .B(n_863), .Y(n_984) );
HB1xp67_ASAP7_75t_L g985 ( .A(n_957), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_955), .Y(n_986) );
OR2x2_ASAP7_75t_L g987 ( .A(n_936), .B(n_863), .Y(n_987) );
AND2x2_ASAP7_75t_L g988 ( .A(n_961), .B(n_890), .Y(n_988) );
AND2x2_ASAP7_75t_L g989 ( .A(n_961), .B(n_890), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_935), .B(n_865), .Y(n_990) );
AND2x2_ASAP7_75t_L g991 ( .A(n_978), .B(n_941), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_978), .B(n_941), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_964), .Y(n_993) );
INVx2_ASAP7_75t_L g994 ( .A(n_976), .Y(n_994) );
INVx6_ASAP7_75t_L g995 ( .A(n_970), .Y(n_995) );
INVxp67_ASAP7_75t_L g996 ( .A(n_985), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_965), .B(n_953), .Y(n_997) );
AND2x2_ASAP7_75t_L g998 ( .A(n_974), .B(n_942), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_965), .B(n_953), .Y(n_999) );
AND2x4_ASAP7_75t_L g1000 ( .A(n_990), .B(n_944), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_974), .B(n_942), .Y(n_1001) );
INVx1_ASAP7_75t_L g1002 ( .A(n_966), .Y(n_1002) );
INVx1_ASAP7_75t_SL g1003 ( .A(n_979), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_990), .B(n_942), .Y(n_1004) );
BUFx2_ASAP7_75t_L g1005 ( .A(n_979), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_988), .B(n_925), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_966), .Y(n_1007) );
INVx1_ASAP7_75t_SL g1008 ( .A(n_979), .Y(n_1008) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_988), .B(n_942), .Y(n_1009) );
INVx1_ASAP7_75t_SL g1010 ( .A(n_971), .Y(n_1010) );
OR2x2_ASAP7_75t_L g1011 ( .A(n_989), .B(n_936), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_967), .Y(n_1012) );
OR2x2_ASAP7_75t_L g1013 ( .A(n_989), .B(n_928), .Y(n_1013) );
NOR2x1_ASAP7_75t_L g1014 ( .A(n_986), .B(n_933), .Y(n_1014) );
NOR2xp33_ASAP7_75t_L g1015 ( .A(n_968), .B(n_940), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_975), .B(n_944), .Y(n_1016) );
OR2x2_ASAP7_75t_L g1017 ( .A(n_973), .B(n_929), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_975), .B(n_945), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_977), .B(n_945), .Y(n_1019) );
NOR3xp33_ASAP7_75t_L g1020 ( .A(n_984), .B(n_960), .C(n_880), .Y(n_1020) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_977), .B(n_949), .Y(n_1021) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_981), .B(n_949), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_993), .Y(n_1023) );
NOR2xp33_ASAP7_75t_L g1024 ( .A(n_1010), .B(n_880), .Y(n_1024) );
NAND2xp5_ASAP7_75t_SL g1025 ( .A(n_1020), .B(n_943), .Y(n_1025) );
AND2x4_ASAP7_75t_L g1026 ( .A(n_1000), .B(n_969), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_997), .B(n_963), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_997), .B(n_963), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_999), .B(n_962), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_998), .B(n_981), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_1001), .B(n_991), .Y(n_1031) );
NAND2xp5_ASAP7_75t_L g1032 ( .A(n_1022), .B(n_972), .Y(n_1032) );
INVxp33_ASAP7_75t_L g1033 ( .A(n_1015), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_1001), .B(n_983), .Y(n_1034) );
INVx2_ASAP7_75t_L g1035 ( .A(n_994), .Y(n_1035) );
INVxp67_ASAP7_75t_L g1036 ( .A(n_1010), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_1018), .B(n_1019), .Y(n_1037) );
OR2x2_ASAP7_75t_L g1038 ( .A(n_1011), .B(n_982), .Y(n_1038) );
OR2x2_ASAP7_75t_L g1039 ( .A(n_1013), .B(n_987), .Y(n_1039) );
INVx2_ASAP7_75t_L g1040 ( .A(n_1035), .Y(n_1040) );
INVx1_ASAP7_75t_SL g1041 ( .A(n_1024), .Y(n_1041) );
INVx2_ASAP7_75t_L g1042 ( .A(n_1035), .Y(n_1042) );
INVx1_ASAP7_75t_SL g1043 ( .A(n_1037), .Y(n_1043) );
XNOR2xp5_ASAP7_75t_L g1044 ( .A(n_1033), .B(n_980), .Y(n_1044) );
INVxp67_ASAP7_75t_L g1045 ( .A(n_1036), .Y(n_1045) );
OAI221xp5_ASAP7_75t_L g1046 ( .A1(n_1025), .A2(n_1014), .B1(n_996), .B2(n_1005), .C(n_1008), .Y(n_1046) );
INVxp33_ASAP7_75t_L g1047 ( .A(n_1032), .Y(n_1047) );
AOI22xp5_ASAP7_75t_L g1048 ( .A1(n_1027), .A2(n_1000), .B1(n_1021), .B2(n_1018), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1023), .Y(n_1049) );
AOI222xp33_ASAP7_75t_L g1050 ( .A1(n_1028), .A2(n_1021), .B1(n_1018), .B2(n_1019), .C1(n_1006), .C2(n_991), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1023), .Y(n_1051) );
AOI22xp5_ASAP7_75t_L g1052 ( .A1(n_1029), .A2(n_1000), .B1(n_1021), .B2(n_1019), .Y(n_1052) );
NAND2xp5_ASAP7_75t_SL g1053 ( .A(n_1026), .B(n_1003), .Y(n_1053) );
OAI22xp5_ASAP7_75t_L g1054 ( .A1(n_1038), .A2(n_937), .B1(n_995), .B2(n_1003), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1049), .Y(n_1055) );
AOI21xp5_ASAP7_75t_L g1056 ( .A1(n_1053), .A2(n_939), .B(n_1026), .Y(n_1056) );
OAI32xp33_ASAP7_75t_L g1057 ( .A1(n_1053), .A2(n_1038), .A3(n_1039), .B1(n_1008), .B2(n_1031), .Y(n_1057) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_1050), .B(n_1030), .Y(n_1058) );
OAI31xp33_ASAP7_75t_SL g1059 ( .A1(n_1054), .A2(n_1026), .A3(n_1034), .B(n_992), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_1041), .B(n_1009), .Y(n_1060) );
INVxp67_ASAP7_75t_SL g1061 ( .A(n_1045), .Y(n_1061) );
OAI22xp5_ASAP7_75t_L g1062 ( .A1(n_1058), .A2(n_1052), .B1(n_1048), .B2(n_1046), .Y(n_1062) );
AOI221xp5_ASAP7_75t_L g1063 ( .A1(n_1057), .A2(n_1044), .B1(n_1047), .B2(n_1043), .C(n_1051), .Y(n_1063) );
O2A1O1Ixp33_ASAP7_75t_L g1064 ( .A1(n_1061), .A2(n_915), .B(n_1042), .C(n_1040), .Y(n_1064) );
INVx2_ASAP7_75t_L g1065 ( .A(n_1055), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1065), .Y(n_1066) );
AOI221xp5_ASAP7_75t_SL g1067 ( .A1(n_1062), .A2(n_1056), .B1(n_1060), .B2(n_1059), .C(n_1004), .Y(n_1067) );
AND4x1_ASAP7_75t_L g1068 ( .A(n_1063), .B(n_912), .C(n_1004), .D(n_1016), .Y(n_1068) );
NOR2xp67_ASAP7_75t_L g1069 ( .A(n_1066), .B(n_1064), .Y(n_1069) );
NOR4xp25_ASAP7_75t_L g1070 ( .A(n_1067), .B(n_1002), .C(n_1012), .D(n_1007), .Y(n_1070) );
NOR3xp33_ASAP7_75t_SL g1071 ( .A(n_1070), .B(n_1068), .C(n_934), .Y(n_1071) );
OR2x2_ASAP7_75t_L g1072 ( .A(n_1069), .B(n_1017), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1072), .Y(n_1073) );
A2O1A1Ixp33_ASAP7_75t_L g1074 ( .A1(n_1073), .A2(n_1071), .B(n_914), .C(n_888), .Y(n_1074) );
AOI221xp5_ASAP7_75t_L g1075 ( .A1(n_1074), .A2(n_914), .B1(n_888), .B2(n_881), .C(n_874), .Y(n_1075) );
AOI21xp5_ASAP7_75t_L g1076 ( .A1(n_1075), .A2(n_881), .B(n_860), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_1076), .B(n_954), .Y(n_1077) );
AOI21xp33_ASAP7_75t_L g1078 ( .A1(n_1077), .A2(n_860), .B(n_874), .Y(n_1078) );
endmodule