module fake_jpeg_29670_n_392 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_392);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_392;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_22),
.B(n_9),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_64),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_54),
.B(n_83),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_22),
.B(n_8),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_23),
.B(n_10),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_76),
.Y(n_110)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_69),
.Y(n_101)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_81),
.A2(n_84),
.B1(n_42),
.B2(n_39),
.Y(n_100)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_42),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_26),
.B(n_10),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_33),
.B1(n_32),
.B2(n_41),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_86),
.A2(n_107),
.B1(n_29),
.B2(n_28),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_103),
.B(n_104),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_67),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_48),
.A2(n_31),
.B1(n_26),
.B2(n_33),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_113),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_63),
.A2(n_42),
.B1(n_19),
.B2(n_37),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_32),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_120),
.B(n_124),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_31),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_59),
.B(n_41),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_29),
.B(n_28),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_133),
.Y(n_168)
);

NOR2x1_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_161),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_74),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_20),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_135),
.C(n_160),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_20),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_117),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_138),
.A2(n_145),
.B1(n_157),
.B2(n_159),
.Y(n_182)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_142),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_121),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_148),
.Y(n_169)
);

BUFx8_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_144),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_97),
.A2(n_38),
.B1(n_65),
.B2(n_53),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_109),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_149),
.B(n_158),
.Y(n_166)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_151),
.Y(n_171)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_85),
.A2(n_50),
.B1(n_61),
.B2(n_57),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_153),
.A2(n_100),
.B1(n_114),
.B2(n_98),
.Y(n_176)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_156),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_105),
.Y(n_156)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_90),
.Y(n_157)
);

AOI21xp33_ASAP7_75t_L g158 ( 
.A1(n_118),
.A2(n_110),
.B(n_89),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_97),
.A2(n_49),
.B1(n_51),
.B2(n_77),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_93),
.A2(n_27),
.B1(n_44),
.B2(n_3),
.Y(n_160)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_139),
.A2(n_90),
.B1(n_95),
.B2(n_98),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_172),
.A2(n_153),
.B1(n_182),
.B2(n_95),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_134),
.B(n_110),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_135),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_176),
.A2(n_154),
.B1(n_133),
.B2(n_99),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_154),
.A2(n_126),
.B(n_108),
.C(n_125),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_178),
.A2(n_125),
.B(n_136),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_183),
.A2(n_198),
.B1(n_182),
.B2(n_178),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_184),
.B(n_192),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_133),
.C(n_152),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_162),
.C(n_176),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_168),
.B(n_132),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_193),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_189),
.A2(n_171),
.B(n_178),
.Y(n_209)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_190),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_192),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_169),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_137),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_168),
.B(n_146),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_194),
.B(n_196),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_195),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_162),
.B(n_170),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_169),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_197),
.Y(n_215)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_141),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_170),
.Y(n_212)
);

NAND3xp33_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_166),
.C(n_175),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_216),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_210),
.C(n_187),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_209),
.A2(n_218),
.B(n_183),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_180),
.C(n_166),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_219),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_213),
.B(n_190),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_214),
.A2(n_183),
.B1(n_193),
.B2(n_197),
.Y(n_228)
);

AOI32xp33_ASAP7_75t_L g216 ( 
.A1(n_196),
.A2(n_171),
.A3(n_172),
.B1(n_164),
.B2(n_163),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_200),
.A2(n_177),
.B(n_163),
.Y(n_218)
);

NOR2x1_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_177),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_203),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_220),
.Y(n_247)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_204),
.Y(n_221)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_221),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_213),
.B(n_184),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_223),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_234),
.C(n_207),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_198),
.B1(n_219),
.B2(n_188),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_225),
.A2(n_214),
.B1(n_206),
.B2(n_218),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_203),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_227),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_235),
.B1(n_209),
.B2(n_219),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_186),
.Y(n_229)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_230),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_231),
.A2(n_232),
.B(n_219),
.Y(n_246)
);

XOR2x2_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_198),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_173),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_233),
.B(n_236),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_199),
.C(n_174),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_214),
.A2(n_164),
.B1(n_185),
.B2(n_195),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_167),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_206),
.Y(n_237)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_238),
.A2(n_205),
.B1(n_179),
.B2(n_167),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_239),
.A2(n_221),
.B1(n_217),
.B2(n_205),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_215),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_240),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_241),
.B(n_243),
.C(n_242),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_201),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_179),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_210),
.C(n_218),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_220),
.B(n_216),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_245),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_246),
.A2(n_232),
.B(n_211),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_225),
.A2(n_226),
.B1(n_227),
.B2(n_231),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_250),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_226),
.A2(n_210),
.B1(n_211),
.B2(n_208),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_208),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_230),
.Y(n_259)
);

OAI32xp33_ASAP7_75t_L g258 ( 
.A1(n_249),
.A2(n_222),
.A3(n_228),
.B1(n_237),
.B2(n_232),
.Y(n_258)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_259),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_255),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_260),
.B(n_264),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_262),
.A2(n_263),
.B(n_256),
.Y(n_285)
);

OA21x2_ASAP7_75t_L g263 ( 
.A1(n_246),
.A2(n_235),
.B(n_204),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_255),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_266),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_238),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_269),
.A2(n_239),
.B1(n_244),
.B2(n_254),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_195),
.Y(n_270)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_251),
.Y(n_271)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_167),
.Y(n_272)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

AND2x2_ASAP7_75t_SL g273 ( 
.A(n_254),
.B(n_195),
.Y(n_273)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_248),
.A2(n_252),
.B1(n_245),
.B2(n_251),
.Y(n_274)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

BUFx12f_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_275),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_241),
.C(n_243),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_279),
.B(n_286),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_284),
.C(n_292),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_283),
.A2(n_288),
.B1(n_273),
.B2(n_263),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_250),
.C(n_256),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_285),
.A2(n_101),
.B(n_142),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_267),
.B(n_160),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_265),
.A2(n_185),
.B1(n_165),
.B2(n_140),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_261),
.B(n_144),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_290),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_185),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_150),
.C(n_161),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_258),
.B(n_144),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_94),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_278),
.A2(n_295),
.B1(n_281),
.B2(n_257),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_300),
.A2(n_303),
.B1(n_316),
.B2(n_318),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_287),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_301),
.B(n_304),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_268),
.C(n_269),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_306),
.C(n_313),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_277),
.A2(n_259),
.B1(n_264),
.B2(n_260),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_296),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_305),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_270),
.C(n_273),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_291),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_309),
.B(n_310),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_298),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_283),
.B(n_263),
.Y(n_311)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_311),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_277),
.A2(n_275),
.B1(n_157),
.B2(n_130),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_314),
.C(n_290),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_279),
.B(n_275),
.C(n_148),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_275),
.C(n_151),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_129),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_315),
.B(n_319),
.Y(n_323)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_294),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_317),
.B(n_320),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_297),
.A2(n_122),
.B1(n_155),
.B2(n_102),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_293),
.B(n_147),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_322),
.B(n_336),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_299),
.A2(n_285),
.B(n_282),
.Y(n_327)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_327),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_289),
.Y(n_330)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_330),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_299),
.B(n_286),
.C(n_99),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_331),
.B(n_332),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_306),
.B(n_116),
.C(n_122),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_307),
.B(n_112),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_333),
.B(n_335),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_112),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_308),
.B(n_123),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_317),
.B(n_101),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_337),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_321),
.A2(n_313),
.B(n_314),
.Y(n_338)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_338),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_321),
.B(n_308),
.C(n_105),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_339),
.B(n_116),
.C(n_84),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_329),
.A2(n_13),
.B1(n_17),
.B2(n_3),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_342),
.A2(n_49),
.B1(n_12),
.B2(n_4),
.Y(n_360)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_325),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_344),
.B(n_347),
.Y(n_355)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_326),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_328),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_348),
.B(n_336),
.Y(n_352)
);

AOI21x1_ASAP7_75t_L g350 ( 
.A1(n_323),
.A2(n_330),
.B(n_329),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_350),
.A2(n_341),
.B(n_349),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_339),
.B(n_324),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_351),
.B(n_352),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_345),
.B(n_334),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_353),
.B(n_356),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_345),
.B(n_334),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_354),
.B(n_6),
.C(n_16),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_343),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_357),
.B(n_360),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_358),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_340),
.B(n_12),
.Y(n_359)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_359),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_349),
.B(n_81),
.C(n_11),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_361),
.B(n_13),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_362),
.A2(n_346),
.B(n_13),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_363),
.A2(n_367),
.B(n_4),
.Y(n_375)
);

AOI21xp33_ASAP7_75t_L g367 ( 
.A1(n_355),
.A2(n_7),
.B(n_17),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_368),
.B(n_369),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_354),
.B(n_44),
.C(n_6),
.Y(n_369)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_371),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_365),
.B(n_356),
.C(n_357),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_374),
.A2(n_379),
.B(n_370),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_375),
.B(n_377),
.C(n_378),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_372),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_366),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_364),
.B(n_4),
.C(n_5),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_380),
.A2(n_16),
.B1(n_1),
.B2(n_0),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_373),
.A2(n_368),
.B(n_369),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_381),
.A2(n_5),
.B(n_14),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_376),
.A2(n_5),
.B(n_14),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_383),
.A2(n_16),
.B(n_1),
.Y(n_386)
);

AO21x1_ASAP7_75t_L g388 ( 
.A1(n_384),
.A2(n_385),
.B(n_386),
.Y(n_388)
);

NOR3xp33_ASAP7_75t_SL g387 ( 
.A(n_384),
.B(n_382),
.C(n_44),
.Y(n_387)
);

INVx11_ASAP7_75t_L g389 ( 
.A(n_387),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_389),
.B(n_388),
.C(n_44),
.Y(n_390)
);

AOI21x1_ASAP7_75t_L g391 ( 
.A1(n_390),
.A2(n_389),
.B(n_1),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_391),
.B(n_1),
.Y(n_392)
);


endmodule