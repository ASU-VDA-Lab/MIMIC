module fake_jpeg_6949_n_289 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_289);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVxp33_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_2),
.B(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_28),
.A2(n_30),
.B1(n_34),
.B2(n_37),
.Y(n_41)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g37 ( 
.A(n_23),
.B(n_13),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_37),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_46),
.Y(n_67)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_47),
.B(n_23),
.Y(n_68)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_53),
.Y(n_79)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_37),
.B(n_30),
.C(n_33),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_30),
.B1(n_29),
.B2(n_33),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_37),
.B1(n_29),
.B2(n_33),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_31),
.B1(n_30),
.B2(n_28),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_46),
.B(n_41),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_68),
.B(n_18),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_33),
.B1(n_31),
.B2(n_29),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_15),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_34),
.Y(n_78)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_13),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_66),
.B(n_26),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_69),
.A2(n_70),
.B1(n_72),
.B2(n_81),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_29),
.B1(n_31),
.B2(n_28),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_54),
.B(n_30),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_80),
.C(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_83),
.Y(n_89)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_49),
.C(n_42),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_54),
.A2(n_31),
.B1(n_28),
.B2(n_49),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_28),
.B1(n_38),
.B2(n_34),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_15),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_64),
.Y(n_88)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_63),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_88),
.B(n_96),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_90),
.Y(n_124)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_93),
.Y(n_121)
);

AO22x1_ASAP7_75t_SL g92 ( 
.A1(n_71),
.A2(n_55),
.B1(n_68),
.B2(n_66),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_92),
.A2(n_59),
.B1(n_60),
.B2(n_75),
.Y(n_122)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_94),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_104),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_59),
.Y(n_100)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_85),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_66),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_106),
.Y(n_125)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_70),
.C(n_71),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_116),
.C(n_117),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_80),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_114),
.B(n_119),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_91),
.A2(n_84),
.B(n_69),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_74),
.C(n_84),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_51),
.C(n_61),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_91),
.A2(n_77),
.B(n_65),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_36),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_122),
.Y(n_137)
);

FAx1_ASAP7_75t_SL g123 ( 
.A(n_89),
.B(n_36),
.CI(n_26),
.CON(n_123),
.SN(n_123)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_128),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_34),
.Y(n_128)
);

OAI32xp33_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_106),
.A3(n_102),
.B1(n_95),
.B2(n_99),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_149),
.Y(n_159)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_131),
.Y(n_154)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_127),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_132),
.B(n_111),
.Y(n_166)
);

AOI21xp33_ASAP7_75t_L g133 ( 
.A1(n_125),
.A2(n_88),
.B(n_104),
.Y(n_133)
);

NOR4xp25_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_17),
.C(n_25),
.D(n_14),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_122),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_135),
.Y(n_163)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_119),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_141),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_101),
.Y(n_139)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_101),
.Y(n_140)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_75),
.Y(n_142)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_146),
.Y(n_170)
);

OA22x2_ASAP7_75t_SL g145 ( 
.A1(n_120),
.A2(n_102),
.B1(n_32),
.B2(n_35),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_SL g172 ( 
.A1(n_145),
.A2(n_23),
.B(n_35),
.Y(n_172)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_90),
.Y(n_148)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_103),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_36),
.C(n_97),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_151),
.C(n_26),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_116),
.C(n_114),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_18),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_19),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_134),
.A2(n_112),
.B1(n_117),
.B2(n_124),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_153),
.A2(n_151),
.B1(n_150),
.B2(n_143),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_149),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_152),
.Y(n_199)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_148),
.A2(n_123),
.B(n_126),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_162),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_126),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_164),
.C(n_171),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_115),
.Y(n_162)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_108),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_169),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_147),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_108),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_93),
.C(n_53),
.Y(n_171)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_172),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_131),
.B(n_17),
.Y(n_173)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_15),
.Y(n_175)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_141),
.Y(n_176)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_129),
.Y(n_180)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_163),
.A2(n_138),
.B1(n_130),
.B2(n_135),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_182),
.A2(n_190),
.B1(n_159),
.B2(n_177),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_154),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_192),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_86),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_189),
.Y(n_205)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

XOR2x2_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_145),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_158),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_53),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_198),
.Y(n_212)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_145),
.C(n_147),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_164),
.C(n_153),
.Y(n_204)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_168),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_180),
.A2(n_159),
.B1(n_165),
.B2(n_169),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_202),
.A2(n_197),
.B1(n_181),
.B2(n_191),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_203),
.B(n_187),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_207),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_21),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_145),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_211),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_185),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_175),
.C(n_132),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_213),
.A2(n_191),
.B(n_178),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_52),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_216),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_193),
.A2(n_14),
.B1(n_18),
.B2(n_25),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_215),
.A2(n_217),
.B1(n_186),
.B2(n_205),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_21),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_179),
.A2(n_14),
.B1(n_25),
.B2(n_27),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_198),
.Y(n_218)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_218),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_213),
.B(n_184),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_219),
.B(n_233),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_235),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_225),
.C(n_204),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_212),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_223),
.A2(n_22),
.B1(n_27),
.B2(n_20),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_188),
.Y(n_224)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_234),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_206),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_232),
.A2(n_22),
.B1(n_19),
.B2(n_16),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_216),
.B(n_16),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_200),
.B(n_16),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_21),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_237),
.A2(n_245),
.B(n_246),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_206),
.C(n_207),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_241),
.C(n_226),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_201),
.C(n_214),
.Y(n_241)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_243),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_232),
.A2(n_27),
.B1(n_22),
.B2(n_19),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_244),
.A2(n_10),
.B1(n_11),
.B2(n_8),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_221),
.Y(n_245)
);

BUFx4f_ASAP7_75t_SL g249 ( 
.A(n_229),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_249),
.A2(n_231),
.B(n_21),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_235),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_250),
.A2(n_255),
.B(n_259),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_261),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_256),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_242),
.A2(n_231),
.B1(n_226),
.B2(n_62),
.Y(n_253)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_20),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_249),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_257),
.B(n_240),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_62),
.C(n_1),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_35),
.Y(n_260)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_260),
.Y(n_271)
);

NOR3xp33_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_7),
.C(n_11),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_254),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_0),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_236),
.Y(n_266)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_266),
.Y(n_273)
);

AOI222xp33_ASAP7_75t_L g267 ( 
.A1(n_259),
.A2(n_249),
.B1(n_240),
.B2(n_246),
.C1(n_8),
.C2(n_10),
.Y(n_267)
);

AOI322xp5_ASAP7_75t_L g272 ( 
.A1(n_267),
.A2(n_7),
.A3(n_1),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_269),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_258),
.A2(n_252),
.B1(n_7),
.B2(n_2),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_0),
.C(n_1),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_265),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_35),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_275),
.A2(n_277),
.B(n_269),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_264),
.B(n_20),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_276),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_263),
.Y(n_282)
);

AOI322xp5_ASAP7_75t_L g283 ( 
.A1(n_279),
.A2(n_280),
.A3(n_282),
.B1(n_274),
.B2(n_273),
.C1(n_275),
.C2(n_268),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_283),
.A2(n_284),
.B(n_3),
.Y(n_285)
);

AOI322xp5_ASAP7_75t_L g284 ( 
.A1(n_281),
.A2(n_32),
.A3(n_35),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_0),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_4),
.Y(n_286)
);

OAI321xp33_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_32),
.C(n_249),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_5),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_288),
.A2(n_6),
.B(n_32),
.Y(n_289)
);


endmodule