module fake_jpeg_2679_n_57 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_57);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_57;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_5),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

NAND2xp33_ASAP7_75t_SL g10 ( 
.A(n_1),
.B(n_0),
.Y(n_10)
);

BUFx24_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_5),
.B(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_6),
.B(n_1),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_0),
.Y(n_19)
);

AND2x2_ASAP7_75t_SL g27 ( 
.A(n_19),
.B(n_16),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_21),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_3),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_24),
.Y(n_30)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_11),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_4),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_22),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_19),
.A2(n_16),
.B1(n_9),
.B2(n_8),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_28),
.A2(n_31),
.B1(n_23),
.B2(n_11),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_19),
.A2(n_9),
.B1(n_8),
.B2(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_24),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_38),
.C(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_21),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_31),
.B(n_28),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_18),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_27),
.C(n_29),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_29),
.C(n_23),
.Y(n_47)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_30),
.B(n_39),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_11),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_6),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_46),
.B(n_47),
.Y(n_51)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_49),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_41),
.B1(n_45),
.B2(n_17),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_49),
.B(n_18),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_55),
.C(n_53),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_7),
.B(n_51),
.Y(n_55)
);

NAND2xp33_ASAP7_75t_R g57 ( 
.A(n_56),
.B(n_7),
.Y(n_57)
);


endmodule