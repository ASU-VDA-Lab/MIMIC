module fake_jpeg_7301_n_261 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_261);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_261;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_34),
.Y(n_40)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_18),
.B1(n_26),
.B2(n_16),
.Y(n_39)
);

AND2x4_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_20),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_17),
.Y(n_57)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_48),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_29),
.A2(n_18),
.B1(n_26),
.B2(n_16),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_18),
.B1(n_16),
.B2(n_26),
.Y(n_66)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g76 ( 
.A(n_57),
.B(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_13),
.Y(n_61)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_13),
.Y(n_63)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_14),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_67),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_73),
.B1(n_35),
.B2(n_40),
.Y(n_84)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_36),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVxp67_ASAP7_75t_SL g92 ( 
.A(n_70),
.Y(n_92)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_36),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_14),
.C(n_40),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_74),
.Y(n_100)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_80),
.Y(n_96)
);

AO22x2_ASAP7_75t_L g79 ( 
.A1(n_73),
.A2(n_14),
.B1(n_25),
.B2(n_37),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_73),
.B1(n_62),
.B2(n_70),
.Y(n_99)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_85),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_84),
.A2(n_64),
.B1(n_40),
.B2(n_53),
.Y(n_103)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_87),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_69),
.Y(n_104)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_93),
.Y(n_108)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_94),
.B(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_60),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_109),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_73),
.B1(n_64),
.B2(n_66),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_73),
.B1(n_64),
.B2(n_51),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_112),
.C(n_34),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_79),
.A2(n_57),
.B1(n_72),
.B2(n_41),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_105),
.A2(n_76),
.B1(n_77),
.B2(n_89),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_77),
.A2(n_14),
.B1(n_53),
.B2(n_68),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_67),
.B(n_65),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_63),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_75),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_92),
.Y(n_130)
);

XNOR2x1_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_56),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_61),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_114),
.A2(n_133),
.B1(n_106),
.B2(n_127),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_111),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_116),
.B(n_119),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_68),
.B1(n_50),
.B2(n_54),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_81),
.B1(n_108),
.B2(n_75),
.Y(n_148)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_88),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_127),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_96),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_129),
.Y(n_153)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_132),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_125),
.A2(n_134),
.B(n_25),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_101),
.A2(n_82),
.B1(n_45),
.B2(n_50),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_126),
.A2(n_123),
.B1(n_97),
.B2(n_100),
.Y(n_138)
);

INVx3_ASAP7_75t_SL g128 ( 
.A(n_107),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_128),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_109),
.Y(n_129)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_131),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_85),
.C(n_80),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_45),
.B1(n_54),
.B2(n_68),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_129),
.A2(n_134),
.B1(n_133),
.B2(n_103),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_136),
.A2(n_117),
.B1(n_126),
.B2(n_123),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_113),
.B(n_102),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_137),
.A2(n_141),
.B(n_145),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_138),
.A2(n_148),
.B1(n_19),
.B2(n_25),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_99),
.B(n_97),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_146),
.B1(n_155),
.B2(n_116),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_121),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_147),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_125),
.A2(n_94),
.B1(n_95),
.B2(n_110),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_114),
.A2(n_108),
.B1(n_93),
.B2(n_86),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_128),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_150),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_128),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_154),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_131),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_117),
.A2(n_91),
.B1(n_47),
.B2(n_49),
.Y(n_155)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_159),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_158),
.A2(n_149),
.B1(n_135),
.B2(n_154),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_153),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_162),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_142),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_132),
.C(n_120),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_170),
.C(n_172),
.Y(n_178)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_166),
.Y(n_186)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_167),
.A2(n_138),
.B1(n_141),
.B2(n_145),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_124),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_137),
.Y(n_187)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_122),
.C(n_91),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_78),
.C(n_25),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_146),
.A2(n_27),
.B1(n_21),
.B2(n_22),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_173),
.A2(n_175),
.B1(n_21),
.B2(n_27),
.Y(n_183)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_144),
.A2(n_27),
.B1(n_23),
.B2(n_22),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_176),
.B(n_143),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_187),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_183),
.B(n_195),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_171),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_185),
.A2(n_189),
.B(n_177),
.Y(n_210)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_171),
.Y(n_189)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_135),
.B1(n_139),
.B2(n_22),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_191),
.A2(n_194),
.B1(n_183),
.B2(n_166),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_158),
.A2(n_23),
.B1(n_21),
.B2(n_24),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_165),
.A2(n_23),
.B1(n_24),
.B2(n_15),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_181),
.A2(n_164),
.B(n_176),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_196),
.A2(n_200),
.B(n_206),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_199),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_180),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_181),
.A2(n_164),
.B(n_160),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_193),
.A2(n_160),
.B(n_170),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_168),
.C(n_163),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_209),
.C(n_211),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g208 ( 
.A(n_187),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_210),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_178),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_167),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_203),
.A2(n_192),
.B1(n_193),
.B2(n_157),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_213),
.A2(n_201),
.B1(n_205),
.B2(n_202),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_200),
.A2(n_186),
.B(n_172),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_217),
.C(n_218),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_191),
.Y(n_216)
);

OA21x2_ASAP7_75t_L g228 ( 
.A1(n_216),
.A2(n_8),
.B(n_12),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_194),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_192),
.C(n_175),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_204),
.A2(n_9),
.B(n_12),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_223),
.C(n_224),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_15),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_17),
.C(n_19),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_212),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_231),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_228),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_24),
.C(n_15),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_232),
.C(n_234),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_19),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_220),
.B(n_11),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g233 ( 
.A1(n_219),
.A2(n_11),
.B(n_10),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_233),
.A2(n_0),
.B(n_2),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_11),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_0),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_2),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_214),
.C(n_221),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_238),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_224),
.C(n_10),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_10),
.C(n_8),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_241),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_0),
.C(n_2),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_7),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_244),
.B(n_3),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_228),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_236),
.C(n_4),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_249),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_242),
.A2(n_7),
.B(n_4),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_250),
.A2(n_3),
.B(n_4),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_251),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_252),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_3),
.C(n_5),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_256),
.A2(n_247),
.B(n_253),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_257),
.A2(n_255),
.B1(n_254),
.B2(n_249),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_258),
.B(n_5),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_259),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_6),
.Y(n_261)
);


endmodule