module real_aes_10774_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_733;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_756;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
INVx1_ASAP7_75t_L g196 ( .A(n_0), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_1), .B(n_252), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_2), .B(n_177), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_3), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_4), .B(n_176), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_5), .A2(n_102), .B1(n_114), .B2(n_880), .Y(n_101) );
INVx1_ASAP7_75t_L g113 ( .A(n_6), .Y(n_113) );
NOR2xp67_ASAP7_75t_L g121 ( .A(n_6), .B(n_85), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_7), .B(n_150), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_8), .B(n_143), .Y(n_598) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_9), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_10), .Y(n_326) );
NAND2x1p5_ASAP7_75t_L g552 ( .A(n_11), .B(n_143), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_12), .B(n_274), .Y(n_622) );
CKINVDCx5p33_ASAP7_75t_R g876 ( .A(n_13), .Y(n_876) );
AOI22xp5_ASAP7_75t_L g871 ( .A1(n_14), .A2(n_98), .B1(n_872), .B2(n_873), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_14), .Y(n_872) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_15), .B(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g579 ( .A(n_16), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_17), .B(n_159), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_18), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_19), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_20), .B(n_150), .Y(n_242) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_21), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_22), .B(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_23), .B(n_168), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_24), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_25), .B(n_190), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_26), .B(n_159), .Y(n_255) );
NAND2xp33_ASAP7_75t_L g548 ( .A(n_27), .B(n_176), .Y(n_548) );
NAND2xp33_ASAP7_75t_L g597 ( .A(n_28), .B(n_176), .Y(n_597) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_29), .Y(n_151) );
OAI21xp33_ASAP7_75t_L g273 ( .A1(n_30), .A2(n_184), .B(n_274), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_31), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_32), .B(n_150), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_33), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_34), .B(n_187), .Y(n_551) );
INVx1_ASAP7_75t_L g110 ( .A(n_35), .Y(n_110) );
OAI21x1_ASAP7_75t_L g145 ( .A1(n_36), .A2(n_67), .B(n_146), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_L g582 ( .A1(n_37), .A2(n_155), .B(n_583), .C(n_585), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_38), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_39), .B(n_150), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_40), .Y(n_321) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_41), .B(n_160), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_42), .Y(n_528) );
NAND2xp33_ASAP7_75t_L g625 ( .A(n_43), .B(n_238), .Y(n_625) );
AND2x6_ASAP7_75t_L g165 ( .A(n_44), .B(n_166), .Y(n_165) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_45), .A2(n_81), .B1(n_176), .B2(n_240), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_46), .B(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_47), .B(n_159), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_48), .B(n_584), .Y(n_596) );
NAND2xp33_ASAP7_75t_L g608 ( .A(n_49), .B(n_238), .Y(n_608) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_50), .Y(n_178) );
INVx1_ASAP7_75t_L g166 ( .A(n_51), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_52), .Y(n_569) );
OAI22x1_ASAP7_75t_R g859 ( .A1(n_53), .A2(n_89), .B1(n_860), .B2(n_861), .Y(n_859) );
INVx1_ASAP7_75t_L g861 ( .A(n_53), .Y(n_861) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_54), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_55), .B(n_240), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_56), .B(n_238), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_57), .B(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_58), .B(n_168), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_59), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_60), .B(n_190), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_61), .B(n_252), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g523 ( .A(n_62), .Y(n_523) );
AND2x2_ASAP7_75t_L g108 ( .A(n_63), .B(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g587 ( .A(n_64), .B(n_190), .Y(n_587) );
INVx2_ASAP7_75t_L g208 ( .A(n_65), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_66), .B(n_240), .Y(n_538) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_68), .Y(n_550) );
NAND2xp33_ASAP7_75t_L g537 ( .A(n_69), .B(n_206), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_70), .B(n_160), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_71), .Y(n_116) );
INVx1_ASAP7_75t_L g200 ( .A(n_72), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_73), .B(n_252), .Y(n_624) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_74), .Y(n_329) );
BUFx10_ASAP7_75t_L g127 ( .A(n_75), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_76), .B(n_525), .Y(n_594) );
NAND2xp33_ASAP7_75t_L g541 ( .A(n_77), .B(n_150), .Y(n_541) );
INVx1_ASAP7_75t_L g323 ( .A(n_78), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_79), .B(n_160), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_80), .B(n_176), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_82), .B(n_190), .Y(n_245) );
INVx1_ASAP7_75t_L g211 ( .A(n_83), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g586 ( .A(n_84), .Y(n_586) );
AND2x2_ASAP7_75t_L g112 ( .A(n_85), .B(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g146 ( .A(n_86), .Y(n_146) );
INVx1_ASAP7_75t_L g111 ( .A(n_87), .Y(n_111) );
OR2x2_ASAP7_75t_L g118 ( .A(n_87), .B(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g511 ( .A(n_87), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_87), .B(n_120), .Y(n_879) );
CKINVDCx5p33_ASAP7_75t_R g566 ( .A(n_88), .Y(n_566) );
INVx1_ASAP7_75t_L g860 ( .A(n_89), .Y(n_860) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_90), .B(n_187), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g603 ( .A(n_91), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_92), .B(n_168), .Y(n_627) );
INVx1_ASAP7_75t_L g109 ( .A(n_93), .Y(n_109) );
INVx1_ASAP7_75t_L g578 ( .A(n_94), .Y(n_578) );
CKINVDCx5p33_ASAP7_75t_R g563 ( .A(n_95), .Y(n_563) );
NOR2xp67_ASAP7_75t_L g270 ( .A(n_96), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g570 ( .A(n_97), .B(n_143), .Y(n_570) );
INVx1_ASAP7_75t_L g873 ( .A(n_98), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_99), .B(n_190), .Y(n_542) );
NAND2xp33_ASAP7_75t_L g216 ( .A(n_100), .B(n_190), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
BUFx12f_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g881 ( .A(n_104), .Y(n_881) );
INVx4_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND2x2_ASAP7_75t_SL g105 ( .A(n_106), .B(n_112), .Y(n_105) );
NOR3xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .C(n_111), .Y(n_106) );
INVx4_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x4_ASAP7_75t_L g120 ( .A(n_110), .B(n_121), .Y(n_120) );
OR2x6_ASAP7_75t_L g114 ( .A(n_115), .B(n_122), .Y(n_114) );
INVx1_ASAP7_75t_L g874 ( .A(n_115), .Y(n_874) );
NOR2xp67_ASAP7_75t_SL g115 ( .A(n_116), .B(n_117), .Y(n_115) );
INVx4_ASAP7_75t_L g869 ( .A(n_117), .Y(n_869) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OR2x6_ASAP7_75t_L g125 ( .A(n_120), .B(n_126), .Y(n_125) );
OAI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_128), .B(n_863), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g878 ( .A(n_126), .B(n_879), .Y(n_878) );
INVx2_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
BUFx12f_ASAP7_75t_L g867 ( .A(n_127), .Y(n_867) );
INVx2_ASAP7_75t_SL g128 ( .A(n_129), .Y(n_128) );
OAI22x1_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_858), .B1(n_859), .B2(n_862), .Y(n_129) );
INVx2_ASAP7_75t_L g862 ( .A(n_130), .Y(n_862) );
OAI22x1_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_510), .B1(n_512), .B2(n_857), .Y(n_130) );
XNOR2x1_ASAP7_75t_L g870 ( .A(n_131), .B(n_871), .Y(n_870) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_447), .Y(n_131) );
NOR2x1_ASAP7_75t_L g132 ( .A(n_133), .B(n_374), .Y(n_132) );
NAND3xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_307), .C(n_354), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_289), .Y(n_134) );
OAI21xp33_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_213), .B(n_259), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AOI322xp5_ASAP7_75t_L g455 ( .A1(n_137), .A2(n_304), .A3(n_456), .B1(n_458), .B2(n_460), .C1(n_464), .C2(n_466), .Y(n_455) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_170), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AOI322xp5_ASAP7_75t_L g307 ( .A1(n_139), .A2(n_308), .A3(n_332), .B1(n_335), .B2(n_337), .C1(n_342), .C2(n_346), .Y(n_307) );
AND2x2_ASAP7_75t_L g424 ( .A(n_139), .B(n_170), .Y(n_424) );
AND2x2_ASAP7_75t_L g426 ( .A(n_139), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g476 ( .A(n_139), .Y(n_476) );
OR2x2_ASAP7_75t_L g494 ( .A(n_139), .B(n_470), .Y(n_494) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x4_ASAP7_75t_L g298 ( .A(n_140), .B(n_299), .Y(n_298) );
AND2x4_ASAP7_75t_L g343 ( .A(n_140), .B(n_267), .Y(n_343) );
BUFx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g262 ( .A(n_141), .Y(n_262) );
OAI21x1_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_147), .B(n_167), .Y(n_141) );
OAI21x1_ASAP7_75t_SL g247 ( .A1(n_142), .A2(n_248), .B(n_258), .Y(n_247) );
OAI21x1_ASAP7_75t_L g520 ( .A1(n_142), .A2(n_521), .B(n_530), .Y(n_520) );
OA21x2_ASAP7_75t_L g544 ( .A1(n_142), .A2(n_545), .B(n_552), .Y(n_544) );
OA21x2_ASAP7_75t_L g600 ( .A1(n_142), .A2(n_601), .B(n_609), .Y(n_600) );
OAI21x1_ASAP7_75t_L g617 ( .A1(n_142), .A2(n_521), .B(n_530), .Y(n_617) );
OAI21x1_ASAP7_75t_L g646 ( .A1(n_142), .A2(n_545), .B(n_552), .Y(n_646) );
BUFx4f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_143), .B(n_182), .Y(n_181) );
INVx3_ASAP7_75t_L g234 ( .A(n_143), .Y(n_234) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_143), .A2(n_535), .B(n_542), .Y(n_534) );
INVx4_ASAP7_75t_L g557 ( .A(n_143), .Y(n_557) );
OA21x2_ASAP7_75t_L g640 ( .A1(n_143), .A2(n_535), .B(n_542), .Y(n_640) );
OA21x2_ASAP7_75t_L g672 ( .A1(n_143), .A2(n_535), .B(n_542), .Y(n_672) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g169 ( .A(n_144), .Y(n_169) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g191 ( .A(n_145), .Y(n_191) );
OAI21x1_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_157), .B(n_163), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_152), .B(n_155), .Y(n_148) );
INVx2_ASAP7_75t_L g198 ( .A(n_150), .Y(n_198) );
INVx2_ASAP7_75t_L g252 ( .A(n_150), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_150), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_SL g584 ( .A(n_150), .Y(n_584) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_151), .Y(n_154) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_151), .Y(n_160) );
INVx2_ASAP7_75t_L g177 ( .A(n_151), .Y(n_177) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_151), .Y(n_206) );
INVx1_ASAP7_75t_L g320 ( .A(n_151), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_153), .B(n_200), .Y(n_199) );
INVxp67_ASAP7_75t_L g224 ( .A(n_153), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_153), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g179 ( .A(n_154), .Y(n_179) );
INVx2_ASAP7_75t_L g568 ( .A(n_154), .Y(n_568) );
INVx2_ASAP7_75t_SL g162 ( .A(n_155), .Y(n_162) );
CKINVDCx6p67_ASAP7_75t_R g218 ( .A(n_155), .Y(n_218) );
INVx2_ASAP7_75t_SL g226 ( .A(n_155), .Y(n_226) );
INVx5_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx5_ASAP7_75t_L g174 ( .A(n_156), .Y(n_174) );
BUFx12f_ASAP7_75t_L g184 ( .A(n_156), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_156), .A2(n_523), .B(n_524), .C(n_526), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_161), .B(n_162), .Y(n_157) );
OAI22xp5_ASAP7_75t_L g203 ( .A1(n_159), .A2(n_204), .B1(n_207), .B2(n_208), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_159), .A2(n_176), .B1(n_220), .B2(n_221), .Y(n_219) );
NOR2xp67_ASAP7_75t_L g562 ( .A(n_159), .B(n_563), .Y(n_562) );
INVx5_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
OR2x2_ASAP7_75t_L g325 ( .A(n_160), .B(n_326), .Y(n_325) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_162), .A2(n_560), .B(n_562), .Y(n_559) );
INVx2_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
INVx8_ASAP7_75t_L g244 ( .A(n_164), .Y(n_244) );
OAI21xp5_ASAP7_75t_L g330 ( .A1(n_164), .A2(n_168), .B(n_331), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_164), .A2(n_559), .B(n_564), .Y(n_558) );
NOR2xp67_ASAP7_75t_L g573 ( .A(n_164), .B(n_574), .Y(n_573) );
INVx8_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g182 ( .A(n_165), .Y(n_182) );
AOI21xp33_ASAP7_75t_L g212 ( .A1(n_165), .A2(n_169), .B(n_210), .Y(n_212) );
INVx1_ASAP7_75t_L g228 ( .A(n_165), .Y(n_228) );
BUFx2_ASAP7_75t_L g626 ( .A(n_165), .Y(n_626) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_169), .B(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_169), .B(n_323), .Y(n_322) );
AND2x4_ASAP7_75t_SL g297 ( .A(n_170), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_192), .Y(n_170) );
AND2x2_ASAP7_75t_L g261 ( .A(n_171), .B(n_262), .Y(n_261) );
INVx2_ASAP7_75t_SL g171 ( .A(n_172), .Y(n_171) );
AND2x4_ASAP7_75t_L g283 ( .A(n_172), .B(n_266), .Y(n_283) );
AND2x2_ASAP7_75t_L g334 ( .A(n_172), .B(n_281), .Y(n_334) );
OR2x2_ASAP7_75t_L g345 ( .A(n_172), .B(n_282), .Y(n_345) );
INVx1_ASAP7_75t_L g365 ( .A(n_172), .Y(n_365) );
AND2x2_ASAP7_75t_L g373 ( .A(n_172), .B(n_282), .Y(n_373) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_172), .Y(n_383) );
AND2x2_ASAP7_75t_L g436 ( .A(n_172), .B(n_262), .Y(n_436) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_183), .B(n_189), .Y(n_172) );
OAI21xp33_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_181), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_174), .A2(n_242), .B(n_243), .Y(n_241) );
INVx1_ASAP7_75t_L g257 ( .A(n_174), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_174), .A2(n_540), .B(n_541), .Y(n_539) );
AOI21x1_ASAP7_75t_L g620 ( .A1(n_174), .A2(n_621), .B(n_622), .Y(n_620) );
OAI22xp33_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_178), .B1(n_179), .B2(n_180), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_176), .B(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g187 ( .A(n_177), .Y(n_187) );
INVx2_ASAP7_75t_L g238 ( .A(n_177), .Y(n_238) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_179), .A2(n_186), .B1(n_187), .B2(n_188), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_184), .B(n_185), .Y(n_183) );
BUFx2_ASAP7_75t_L g201 ( .A(n_184), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_184), .Y(n_209) );
INVx3_ASAP7_75t_L g253 ( .A(n_184), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_184), .A2(n_270), .B1(n_273), .B2(n_275), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_184), .A2(n_624), .B(n_625), .Y(n_623) );
NOR2x1p5_ASAP7_75t_SL g227 ( .A(n_190), .B(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g268 ( .A(n_190), .Y(n_268) );
BUFx5_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g278 ( .A(n_191), .Y(n_278) );
INVx2_ASAP7_75t_L g264 ( .A(n_192), .Y(n_264) );
AND2x2_ASAP7_75t_L g363 ( .A(n_192), .B(n_262), .Y(n_363) );
AND2x2_ASAP7_75t_L g440 ( .A(n_192), .B(n_404), .Y(n_440) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g282 ( .A(n_193), .Y(n_282) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_202), .B(n_212), .Y(n_193) );
OAI21xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_199), .B(n_201), .Y(n_194) );
NOR2x1_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_197), .A2(n_253), .B(n_528), .C(n_529), .Y(n_527) );
O2A1O1Ixp5_ASAP7_75t_L g549 ( .A1(n_197), .A2(n_253), .B(n_550), .C(n_551), .Y(n_549) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_198), .A2(n_318), .B1(n_319), .B2(n_321), .Y(n_317) );
OAI21x1_ASAP7_75t_L g576 ( .A1(n_201), .A2(n_577), .B(n_579), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_209), .B(n_210), .Y(n_202) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g240 ( .A(n_206), .Y(n_240) );
INVx2_ASAP7_75t_L g272 ( .A(n_206), .Y(n_272) );
INVx2_ASAP7_75t_L g274 ( .A(n_206), .Y(n_274) );
INVx1_ASAP7_75t_L g525 ( .A(n_206), .Y(n_525) );
AO21x1_ASAP7_75t_L g316 ( .A1(n_209), .A2(n_317), .B(n_322), .Y(n_316) );
AOI21x1_ASAP7_75t_L g324 ( .A1(n_209), .A2(n_325), .B(n_327), .Y(n_324) );
OAI21xp33_ASAP7_75t_L g564 ( .A1(n_209), .A2(n_565), .B(n_567), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_209), .A2(n_593), .B(n_594), .Y(n_592) );
OAI21xp5_ASAP7_75t_L g468 ( .A1(n_213), .A2(n_469), .B(n_471), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_214), .B(n_229), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_214), .B(n_306), .Y(n_360) );
HB1xp67_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g286 ( .A(n_215), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_215), .B(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g341 ( .A(n_215), .Y(n_341) );
AND2x2_ASAP7_75t_L g353 ( .A(n_215), .B(n_287), .Y(n_353) );
INVx1_ASAP7_75t_L g369 ( .A(n_215), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_215), .B(n_339), .Y(n_446) );
INVx1_ASAP7_75t_L g462 ( .A(n_215), .Y(n_462) );
AND2x2_ASAP7_75t_L g479 ( .A(n_215), .B(n_313), .Y(n_479) );
AND2x4_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_222), .C(n_227), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_218), .A2(n_237), .B(n_239), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_218), .A2(n_537), .B(n_538), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_218), .A2(n_547), .B(n_548), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_218), .A2(n_607), .B(n_608), .Y(n_606) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_225), .C(n_226), .Y(n_222) );
AND2x2_ASAP7_75t_L g478 ( .A(n_229), .B(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_229), .B(n_498), .Y(n_497) );
AND2x4_ASAP7_75t_L g229 ( .A(n_230), .B(n_246), .Y(n_229) );
BUFx2_ASAP7_75t_L g288 ( .A(n_230), .Y(n_288) );
INVx1_ASAP7_75t_L g349 ( .A(n_230), .Y(n_349) );
AND2x4_ASAP7_75t_L g394 ( .A(n_230), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g414 ( .A(n_230), .B(n_341), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_230), .B(n_358), .Y(n_451) );
INVx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x4_ASAP7_75t_L g378 ( .A(n_231), .B(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g295 ( .A(n_232), .Y(n_295) );
OAI21x1_ASAP7_75t_SL g232 ( .A1(n_233), .A2(n_235), .B(n_245), .Y(n_232) );
OAI21x1_ASAP7_75t_L g590 ( .A1(n_233), .A2(n_591), .B(n_598), .Y(n_590) );
OAI21xp5_ASAP7_75t_L g618 ( .A1(n_233), .A2(n_619), .B(n_627), .Y(n_618) );
OAI21x1_ASAP7_75t_L g652 ( .A1(n_233), .A2(n_619), .B(n_627), .Y(n_652) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_241), .B(n_244), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_238), .B(n_566), .Y(n_565) );
OAI21x1_ASAP7_75t_SL g248 ( .A1(n_244), .A2(n_249), .B(n_254), .Y(n_248) );
AO31x2_ASAP7_75t_L g267 ( .A1(n_244), .A2(n_268), .A3(n_269), .B(n_276), .Y(n_267) );
OAI21x1_ASAP7_75t_L g521 ( .A1(n_244), .A2(n_522), .B(n_527), .Y(n_521) );
OAI21x1_ASAP7_75t_L g535 ( .A1(n_244), .A2(n_536), .B(n_539), .Y(n_535) );
OAI21x1_ASAP7_75t_L g545 ( .A1(n_244), .A2(n_546), .B(n_549), .Y(n_545) );
OAI21x1_ASAP7_75t_L g591 ( .A1(n_244), .A2(n_592), .B(n_595), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g601 ( .A1(n_244), .A2(n_602), .B(n_606), .Y(n_601) );
AND2x2_ASAP7_75t_L g311 ( .A(n_246), .B(n_295), .Y(n_311) );
AND2x2_ASAP7_75t_L g338 ( .A(n_246), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g350 ( .A(n_246), .B(n_341), .Y(n_350) );
BUFx2_ASAP7_75t_L g377 ( .A(n_246), .Y(n_377) );
INVx2_ASAP7_75t_L g395 ( .A(n_246), .Y(n_395) );
BUFx3_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g287 ( .A(n_247), .Y(n_287) );
AOI21x1_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_251), .B(n_253), .Y(n_249) );
O2A1O1Ixp5_ASAP7_75t_L g602 ( .A1(n_253), .A2(n_603), .B(n_604), .C(n_605), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_256), .B(n_257), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g595 ( .A1(n_257), .A2(n_596), .B(n_597), .Y(n_595) );
OAI21xp5_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_279), .B(n_284), .Y(n_259) );
AND2x4_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
AND2x2_ASAP7_75t_L g335 ( .A(n_261), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g302 ( .A(n_262), .B(n_267), .Y(n_302) );
INVx1_ASAP7_75t_L g409 ( .A(n_262), .Y(n_409) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_262), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_262), .B(n_264), .Y(n_509) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx2_ASAP7_75t_L g301 ( .A(n_264), .Y(n_301) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_265), .Y(n_371) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_SL g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g299 ( .A(n_267), .Y(n_299) );
AND2x2_ASAP7_75t_L g364 ( .A(n_267), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g400 ( .A(n_267), .Y(n_400) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g604 ( .A(n_274), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
INVx1_ASAP7_75t_L g428 ( .A(n_280), .Y(n_428) );
INVxp67_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
AND2x4_ASAP7_75t_L g336 ( .A(n_281), .B(n_299), .Y(n_336) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g427 ( .A(n_283), .B(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g470 ( .A(n_283), .Y(n_470) );
AND2x4_ASAP7_75t_L g284 ( .A(n_285), .B(n_288), .Y(n_284) );
AND2x4_ASAP7_75t_L g304 ( .A(n_285), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g433 ( .A(n_285), .B(n_403), .Y(n_433) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx1_ASAP7_75t_L g293 ( .A(n_287), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_287), .B(n_295), .Y(n_390) );
OR2x2_ASAP7_75t_L g385 ( .A(n_288), .B(n_340), .Y(n_385) );
INVx1_ASAP7_75t_L g444 ( .A(n_288), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_296), .B1(n_300), .B2(n_303), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_293), .B(n_388), .Y(n_463) );
BUFx2_ASAP7_75t_L g490 ( .A(n_293), .Y(n_490) );
OR2x2_ASAP7_75t_L g505 ( .A(n_294), .B(n_312), .Y(n_505) );
INVx2_ASAP7_75t_L g306 ( .A(n_295), .Y(n_306) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AOI221xp5_ASAP7_75t_L g495 ( .A1(n_297), .A2(n_380), .B1(n_445), .B2(n_496), .C(n_499), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_298), .B(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AOI322xp5_ASAP7_75t_L g502 ( .A1(n_301), .A2(n_364), .A3(n_475), .B1(n_503), .B2(n_504), .C1(n_506), .C2(n_507), .Y(n_502) );
INVx1_ASAP7_75t_L g420 ( .A(n_302), .Y(n_420) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_302), .A2(n_387), .B1(n_439), .B2(n_440), .Y(n_438) );
NAND3xp33_ASAP7_75t_L g471 ( .A(n_302), .B(n_334), .C(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g506 ( .A(n_302), .B(n_373), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_303), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g352 ( .A(n_306), .B(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g366 ( .A(n_306), .B(n_367), .Y(n_366) );
AND2x4_ASAP7_75t_L g480 ( .A(n_306), .B(n_368), .Y(n_480) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g507 ( .A(n_310), .B(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_311), .B(n_340), .Y(n_405) );
INVx2_ASAP7_75t_L g393 ( .A(n_312), .Y(n_393) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_314), .Y(n_358) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g339 ( .A(n_315), .Y(n_339) );
BUFx3_ASAP7_75t_L g379 ( .A(n_315), .Y(n_379) );
OAI21x1_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_324), .B(n_330), .Y(n_315) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g581 ( .A(n_320), .Y(n_581) );
INVxp67_ASAP7_75t_L g331 ( .A(n_322), .Y(n_331) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AOI21xp33_ASAP7_75t_L g354 ( .A1(n_332), .A2(n_355), .B(n_359), .Y(n_354) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_332), .A2(n_418), .B1(n_450), .B2(n_452), .Y(n_449) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g419 ( .A(n_333), .B(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_SL g501 ( .A(n_335), .Y(n_501) );
AND2x4_ASAP7_75t_L g407 ( .A(n_336), .B(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_336), .B(n_436), .Y(n_435) );
NOR2x1_ASAP7_75t_L g485 ( .A(n_337), .B(n_486), .Y(n_485) );
AND2x4_ASAP7_75t_SL g337 ( .A(n_338), .B(n_340), .Y(n_337) );
INVx1_ASAP7_75t_L g422 ( .A(n_338), .Y(n_422) );
AND2x2_ASAP7_75t_L g368 ( .A(n_339), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g388 ( .A(n_339), .Y(n_388) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x4_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
AND2x2_ASAP7_75t_L g396 ( .A(n_343), .B(n_372), .Y(n_396) );
INVx1_ASAP7_75t_L g417 ( .A(n_343), .Y(n_417) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_343), .Y(n_431) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g457 ( .A(n_345), .B(n_403), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_351), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x4_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
AND2x2_ASAP7_75t_L g402 ( .A(n_350), .B(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g454 ( .A(n_350), .Y(n_454) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_352), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g466 ( .A(n_357), .B(n_389), .Y(n_466) );
INVx1_ASAP7_75t_L g498 ( .A(n_357), .Y(n_498) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_361), .B1(n_366), .B2(n_370), .Y(n_359) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x4_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx1_ASAP7_75t_L g477 ( .A(n_364), .Y(n_477) );
AND2x2_ASAP7_75t_L g399 ( .A(n_365), .B(n_400), .Y(n_399) );
OAI21xp5_ASAP7_75t_L g429 ( .A1(n_366), .A2(n_430), .B(n_432), .Y(n_429) );
INVx1_ASAP7_75t_L g503 ( .A(n_366), .Y(n_503) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
BUFx3_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_373), .B(n_408), .Y(n_465) );
NAND3xp33_ASAP7_75t_L g374 ( .A(n_375), .B(n_410), .C(n_425), .Y(n_374) );
AOI221xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_380), .B1(n_384), .B2(n_396), .C(n_397), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_376), .A2(n_411), .B1(n_415), .B2(n_418), .C(n_421), .Y(n_410) );
AND2x4_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
AND2x4_ASAP7_75t_L g413 ( .A(n_377), .B(n_414), .Y(n_413) );
AOI211xp5_ASAP7_75t_L g425 ( .A1(n_378), .A2(n_426), .B(n_429), .C(n_437), .Y(n_425) );
INVx2_ASAP7_75t_L g404 ( .A(n_379), .Y(n_404) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g416 ( .A(n_382), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND3xp33_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .C(n_391), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_388), .B(n_414), .Y(n_500) );
INVx1_ASAP7_75t_L g487 ( .A(n_389), .Y(n_487) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
OR2x6_ASAP7_75t_L g453 ( .A(n_393), .B(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g441 ( .A(n_394), .Y(n_441) );
OAI22xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_401), .B1(n_405), .B2(n_406), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g459 ( .A(n_400), .Y(n_459) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI21xp33_ASAP7_75t_L g421 ( .A1(n_405), .A2(n_422), .B(n_423), .Y(n_421) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g469 ( .A(n_408), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_426), .A2(n_474), .B1(n_478), .B2(n_480), .Y(n_473) );
INVx2_ASAP7_75t_SL g442 ( .A(n_427), .Y(n_442) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_433), .B(n_434), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_441), .B1(n_442), .B2(n_443), .Y(n_437) );
BUFx2_ASAP7_75t_L g492 ( .A(n_440), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NOR2xp67_ASAP7_75t_L g447 ( .A(n_448), .B(n_481), .Y(n_447) );
NAND4xp25_ASAP7_75t_SL g448 ( .A(n_449), .B(n_455), .C(n_467), .D(n_473), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g472 ( .A(n_454), .Y(n_472) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx3_ASAP7_75t_L g483 ( .A(n_469), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_477), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g488 ( .A(n_479), .Y(n_488) );
NAND3xp33_ASAP7_75t_L g481 ( .A(n_482), .B(n_495), .C(n_502), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B1(n_489), .B2(n_491), .Y(n_482) );
INVxp67_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NOR2xp67_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NOR2xp67_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g857 ( .A(n_510), .Y(n_857) );
BUFx8_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
AND2x4_ASAP7_75t_L g512 ( .A(n_513), .B(n_765), .Y(n_512) );
NOR4xp25_ASAP7_75t_L g513 ( .A(n_514), .B(n_662), .C(n_706), .D(n_725), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_647), .Y(n_514) );
AOI222xp33_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_553), .B1(n_588), .B2(n_613), .C1(n_628), .C2(n_637), .Y(n_515) );
AOI221xp5_ASAP7_75t_L g844 ( .A1(n_516), .A2(n_670), .B1(n_790), .B2(n_845), .C(n_847), .Y(n_844) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_531), .Y(n_516) );
BUFx2_ASAP7_75t_L g781 ( .A(n_517), .Y(n_781) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x4_ASAP7_75t_L g681 ( .A(n_518), .B(n_666), .Y(n_681) );
AND2x4_ASAP7_75t_L g759 ( .A(n_518), .B(n_760), .Y(n_759) );
AND2x2_ASAP7_75t_L g816 ( .A(n_518), .B(n_756), .Y(n_816) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g642 ( .A(n_520), .Y(n_642) );
HB1xp67_ASAP7_75t_L g762 ( .A(n_520), .Y(n_762) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g721 ( .A(n_531), .B(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVxp67_ASAP7_75t_SL g784 ( .A(n_532), .Y(n_784) );
NAND2x1p5_ASAP7_75t_L g532 ( .A(n_533), .B(n_543), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
OR2x2_ASAP7_75t_L g732 ( .A(n_534), .B(n_644), .Y(n_732) );
AND2x2_ASAP7_75t_L g789 ( .A(n_534), .B(n_644), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_534), .B(n_697), .Y(n_798) );
INVx1_ASAP7_75t_L g614 ( .A(n_543), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_543), .B(n_642), .Y(n_685) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g673 ( .A(n_544), .B(n_650), .Y(n_673) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g763 ( .A(n_555), .B(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_L g808 ( .A(n_555), .B(n_809), .Y(n_808) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_571), .Y(n_555) );
AND2x2_ASAP7_75t_L g654 ( .A(n_556), .B(n_612), .Y(n_654) );
OR2x2_ASAP7_75t_L g661 ( .A(n_556), .B(n_590), .Y(n_661) );
AND2x2_ASAP7_75t_L g814 ( .A(n_556), .B(n_600), .Y(n_814) );
AO21x2_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_558), .B(n_570), .Y(n_556) );
INVx3_ASAP7_75t_L g574 ( .A(n_557), .Y(n_574) );
AO21x2_ASAP7_75t_L g635 ( .A1(n_557), .A2(n_558), .B(n_570), .Y(n_635) );
NOR2xp33_ASAP7_75t_SL g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_568), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g612 ( .A(n_571), .Y(n_612) );
AND2x2_ASAP7_75t_L g714 ( .A(n_571), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g793 ( .A(n_571), .Y(n_793) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g632 ( .A(n_572), .Y(n_632) );
AOI21x1_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_575), .B(n_587), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_582), .Y(n_575) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AOI221xp5_ASAP7_75t_L g726 ( .A1(n_588), .A2(n_727), .B1(n_729), .B2(n_733), .C(n_738), .Y(n_726) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_610), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_589), .B(n_744), .Y(n_743) );
NAND2xp67_ASAP7_75t_L g780 ( .A(n_589), .B(n_654), .Y(n_780) );
AND2x4_ASAP7_75t_L g835 ( .A(n_589), .B(n_714), .Y(n_835) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_599), .Y(n_589) );
INVx1_ASAP7_75t_L g636 ( .A(n_590), .Y(n_636) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_590), .Y(n_657) );
INVx1_ASAP7_75t_L g702 ( .A(n_590), .Y(n_702) );
INVx1_ASAP7_75t_L g751 ( .A(n_590), .Y(n_751) );
AND2x2_ASAP7_75t_L g792 ( .A(n_590), .B(n_793), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_599), .B(n_635), .Y(n_692) );
OR2x2_ASAP7_75t_L g750 ( .A(n_599), .B(n_751), .Y(n_750) );
BUFx3_ASAP7_75t_L g839 ( .A(n_599), .Y(n_839) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g633 ( .A(n_600), .Y(n_633) );
AOI22xp33_ASAP7_75t_SL g840 ( .A1(n_610), .A2(n_681), .B1(n_841), .B2(n_842), .Y(n_840) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g799 ( .A(n_611), .B(n_735), .Y(n_799) );
OR2x2_ASAP7_75t_L g843 ( .A(n_611), .B(n_661), .Y(n_843) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_613), .A2(n_648), .B1(n_653), .B2(n_658), .Y(n_647) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
OR2x2_ASAP7_75t_L g825 ( .A(n_614), .B(n_741), .Y(n_825) );
BUFx3_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g719 ( .A(n_616), .Y(n_719) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
INVx1_ASAP7_75t_L g697 ( .A(n_617), .Y(n_697) );
OR2x2_ASAP7_75t_L g710 ( .A(n_617), .B(n_651), .Y(n_710) );
AND2x2_ASAP7_75t_L g807 ( .A(n_617), .B(n_644), .Y(n_807) );
BUFx2_ASAP7_75t_L g742 ( .A(n_618), .Y(n_742) );
OAI21x1_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_623), .B(n_626), .Y(n_619) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_634), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_631), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g660 ( .A(n_632), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_632), .B(n_633), .Y(n_688) );
INVxp67_ASAP7_75t_SL g745 ( .A(n_632), .Y(n_745) );
OR2x2_ASAP7_75t_L g656 ( .A(n_633), .B(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g736 ( .A(n_633), .Y(n_736) );
AND2x2_ASAP7_75t_L g786 ( .A(n_633), .B(n_702), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_633), .B(n_737), .Y(n_811) );
OR2x2_ASAP7_75t_L g687 ( .A(n_634), .B(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g704 ( .A(n_635), .Y(n_704) );
INVx2_ASAP7_75t_SL g715 ( .A(n_635), .Y(n_715) );
INVx1_ASAP7_75t_L g771 ( .A(n_636), .Y(n_771) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .Y(n_638) );
OR2x2_ASAP7_75t_L g823 ( .A(n_639), .B(n_698), .Y(n_823) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx2_ASAP7_75t_SL g669 ( .A(n_640), .Y(n_669) );
INVx1_ASAP7_75t_SL g680 ( .A(n_640), .Y(n_680) );
BUFx2_ASAP7_75t_L g829 ( .A(n_640), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_641), .B(n_834), .Y(n_833) );
NAND2x1_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
AND2x4_ASAP7_75t_SL g665 ( .A(n_642), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g722 ( .A(n_642), .Y(n_722) );
BUFx2_ASAP7_75t_L g730 ( .A(n_642), .Y(n_730) );
INVx1_ASAP7_75t_L g778 ( .A(n_643), .Y(n_778) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_644), .B(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g668 ( .A(n_644), .B(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g760 ( .A(n_645), .B(n_651), .Y(n_760) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g756 ( .A(n_646), .B(n_651), .Y(n_756) );
AND2x2_ASAP7_75t_L g705 ( .A(n_648), .B(n_672), .Y(n_705) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g761 ( .A(n_649), .B(n_762), .Y(n_761) );
INVx2_ASAP7_75t_L g666 ( .A(n_650), .Y(n_666) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g767 ( .A1(n_653), .A2(n_671), .B1(n_768), .B2(n_773), .Y(n_767) );
AND2x4_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
INVx1_ASAP7_75t_L g723 ( .A(n_654), .Y(n_723) );
INVx1_ASAP7_75t_L g856 ( .A(n_654), .Y(n_856) );
INVx1_ASAP7_75t_L g802 ( .A(n_655), .Y(n_802) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OAI211xp5_ASAP7_75t_L g662 ( .A1(n_659), .A2(n_663), .B(n_674), .C(n_689), .Y(n_662) );
OR2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVx1_ASAP7_75t_L g820 ( .A(n_660), .Y(n_820) );
INVx2_ASAP7_75t_L g737 ( .A(n_661), .Y(n_737) );
INVxp67_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
AO21x1_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_667), .B(n_670), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_665), .B(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g728 ( .A(n_665), .Y(n_728) );
INVx1_ASAP7_75t_L g806 ( .A(n_666), .Y(n_806) );
BUFx2_ASAP7_75t_L g841 ( .A(n_666), .Y(n_841) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NOR2x1_ASAP7_75t_SL g718 ( .A(n_668), .B(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_669), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g749 ( .A(n_669), .Y(n_749) );
AND2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_673), .Y(n_670) );
OR2x6_ASAP7_75t_SL g709 ( .A(n_671), .B(n_710), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_671), .B(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g677 ( .A(n_672), .Y(n_677) );
INVx2_ASAP7_75t_L g698 ( .A(n_673), .Y(n_698) );
OAI31xp33_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_678), .A3(n_682), .B(n_686), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g838 ( .A(n_677), .B(n_839), .Y(n_838) );
AND2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_681), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NOR2x1p5_ASAP7_75t_L g803 ( .A(n_680), .B(n_758), .Y(n_803) );
INVx2_ASAP7_75t_L g772 ( .A(n_681), .Y(n_772) );
INVxp67_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g846 ( .A(n_688), .Y(n_846) );
AOI22xp33_ASAP7_75t_SL g689 ( .A1(n_690), .A2(n_693), .B1(n_699), .B2(n_705), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
OR2x2_ASAP7_75t_L g830 ( .A(n_691), .B(n_701), .Y(n_830) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AOI21xp5_ASAP7_75t_L g738 ( .A1(n_694), .A2(n_739), .B(n_743), .Y(n_738) );
OR2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_698), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_695), .B(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_SL g755 ( .A(n_696), .B(n_756), .Y(n_755) );
BUFx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_703), .Y(n_700) );
INVx1_ASAP7_75t_L g724 ( .A(n_701), .Y(n_724) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
BUFx2_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g791 ( .A(n_704), .B(n_792), .Y(n_791) );
O2A1O1Ixp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_711), .B(n_716), .C(n_724), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVxp67_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_709), .B(n_774), .Y(n_773) );
OR2x2_ASAP7_75t_L g848 ( .A(n_710), .B(n_749), .Y(n_848) );
OAI21xp5_ASAP7_75t_L g850 ( .A1(n_710), .A2(n_851), .B(n_853), .Y(n_850) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g770 ( .A(n_714), .B(n_771), .Y(n_770) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_715), .Y(n_754) );
AO21x1_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_720), .B(n_723), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_719), .A2(n_723), .B1(n_769), .B2(n_772), .Y(n_768) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
OAI21xp5_ASAP7_75t_L g795 ( .A1(n_721), .A2(n_796), .B(n_799), .Y(n_795) );
AND2x2_ASAP7_75t_L g788 ( .A(n_722), .B(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_746), .Y(n_725) );
AND2x2_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g832 ( .A(n_732), .Y(n_832) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx3_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AND2x4_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
AND2x4_ASAP7_75t_L g790 ( .A(n_736), .B(n_791), .Y(n_790) );
OR2x2_ASAP7_75t_L g855 ( .A(n_736), .B(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g834 ( .A(n_742), .Y(n_834) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AOI32xp33_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_752), .A3(n_755), .B1(n_757), .B2(n_763), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OR2x2_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
INVx1_ASAP7_75t_L g775 ( .A(n_749), .Y(n_775) );
INVx1_ASAP7_75t_L g764 ( .A(n_750), .Y(n_764) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_753), .B(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
OAI21xp33_ASAP7_75t_L g853 ( .A1(n_755), .A2(n_808), .B(n_854), .Y(n_853) );
AND2x2_ASAP7_75t_L g828 ( .A(n_756), .B(n_829), .Y(n_828) );
NAND2xp33_ASAP7_75t_SL g757 ( .A(n_758), .B(n_761), .Y(n_757) );
INVx3_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
NOR4xp75_ASAP7_75t_L g765 ( .A(n_766), .B(n_794), .C(n_836), .D(n_850), .Y(n_765) );
NAND3xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_776), .C(n_787), .Y(n_766) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g809 ( .A(n_771), .Y(n_809) );
A2O1A1Ixp33_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_779), .B(n_781), .C(n_782), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
OAI21xp5_ASAP7_75t_L g782 ( .A1(n_781), .A2(n_783), .B(n_785), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g821 ( .A(n_786), .Y(n_821) );
NAND2x1_ASAP7_75t_L g787 ( .A(n_788), .B(n_790), .Y(n_787) );
AND2x4_ASAP7_75t_L g813 ( .A(n_792), .B(n_814), .Y(n_813) );
NAND4xp75_ASAP7_75t_L g794 ( .A(n_795), .B(n_800), .C(n_817), .D(n_826), .Y(n_794) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
HB1xp67_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
AOI211x1_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_803), .B(n_804), .C(n_810), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g817 ( .A1(n_801), .A2(n_818), .B1(n_822), .B2(n_824), .Y(n_817) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
NOR3xp33_ASAP7_75t_L g847 ( .A(n_802), .B(n_848), .C(n_849), .Y(n_847) );
AND2x2_ASAP7_75t_L g804 ( .A(n_805), .B(n_808), .Y(n_804) );
AND2x4_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
AOI21xp5_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_812), .B(n_815), .Y(n_810) );
NOR2xp67_ASAP7_75t_L g852 ( .A(n_812), .B(n_829), .Y(n_852) );
INVx2_ASAP7_75t_SL g812 ( .A(n_813), .Y(n_812) );
INVx2_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
OR2x2_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
INVx1_ASAP7_75t_L g849 ( .A(n_820), .Y(n_849) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
OA21x2_ASAP7_75t_L g826 ( .A1(n_827), .A2(n_830), .B(n_831), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
OAI21xp5_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_833), .B(n_835), .Y(n_831) );
OAI21xp5_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_840), .B(n_844), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
HB1xp67_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVxp67_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx2_ASAP7_75t_SL g858 ( .A(n_859), .Y(n_858) );
AOI21xp5_ASAP7_75t_L g863 ( .A1(n_864), .A2(n_868), .B(n_875), .Y(n_863) );
CKINVDCx5p33_ASAP7_75t_R g864 ( .A(n_865), .Y(n_864) );
CKINVDCx5p33_ASAP7_75t_R g865 ( .A(n_866), .Y(n_865) );
CKINVDCx5p33_ASAP7_75t_R g866 ( .A(n_867), .Y(n_866) );
OAI21xp5_ASAP7_75t_L g868 ( .A1(n_869), .A2(n_870), .B(n_874), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g875 ( .A(n_876), .B(n_877), .Y(n_875) );
BUFx12f_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
CKINVDCx5p33_ASAP7_75t_R g880 ( .A(n_881), .Y(n_880) );
endmodule