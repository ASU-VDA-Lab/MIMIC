module fake_netlist_6_371_n_1690 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1690);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1690;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_12),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_21),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_73),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_129),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g169 ( 
.A(n_36),
.Y(n_169)
);

BUFx10_ASAP7_75t_L g170 ( 
.A(n_163),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_26),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_28),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_15),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_58),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_161),
.Y(n_176)
);

BUFx10_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_108),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_95),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_96),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_51),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_24),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_81),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_154),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_62),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_94),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_38),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_126),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_3),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_131),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_155),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_28),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_137),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_144),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_1),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_122),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_111),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_3),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_97),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_106),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_55),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_43),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_14),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_39),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_136),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_6),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_52),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_49),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_64),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_53),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_8),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_4),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_121),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_140),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_109),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_117),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_47),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_77),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_65),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_83),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_138),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_99),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_92),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_22),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_69),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_47),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_156),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_2),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_1),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_50),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_41),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_2),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_30),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_93),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_132),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_157),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_19),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_35),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_18),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_119),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_115),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_44),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_61),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_60),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_78),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_34),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_145),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_146),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_32),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_40),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_5),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_38),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_128),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_66),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_147),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_127),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_14),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_75),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_135),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_10),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_149),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_134),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_101),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_9),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_22),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_150),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_35),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_29),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_74),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_103),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_53),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_40),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_88),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_43),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_20),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_143),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_104),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_6),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_107),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_27),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_42),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_0),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_85),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_118),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_89),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_18),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_113),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_49),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_37),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_27),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_87),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_19),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_52),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_125),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_34),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_12),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_37),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_102),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_159),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_51),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_63),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_110),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_15),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_76),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_26),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_7),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_86),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_45),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_105),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_130),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g314 ( 
.A(n_91),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_45),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_13),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_39),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_114),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_71),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_98),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_141),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_124),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_10),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_31),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_152),
.Y(n_325)
);

BUFx10_ASAP7_75t_L g326 ( 
.A(n_57),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_123),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_220),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_255),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_255),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_166),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_315),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_315),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_289),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_289),
.Y(n_335)
);

INVxp33_ASAP7_75t_SL g336 ( 
.A(n_166),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_172),
.B(n_0),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_289),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_289),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_200),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_289),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_207),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_233),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_233),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_216),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_270),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_270),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_190),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_196),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_211),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_205),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_215),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_231),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_287),
.B(n_4),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_235),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_171),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_221),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_243),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_240),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_210),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_265),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_213),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_279),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_286),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_214),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_227),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_322),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_229),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_234),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_169),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_236),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_165),
.Y(n_372)
);

INVxp33_ASAP7_75t_SL g373 ( 
.A(n_171),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_245),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_199),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_208),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_241),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_249),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_173),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_254),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_179),
.B(n_5),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_252),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_253),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_204),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_263),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_173),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_260),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_274),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_275),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_283),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_179),
.B(n_7),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_285),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_291),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_298),
.Y(n_394)
);

CKINVDCx14_ASAP7_75t_R g395 ( 
.A(n_169),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_300),
.Y(n_396)
);

BUFx2_ASAP7_75t_SL g397 ( 
.A(n_247),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_267),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_316),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_323),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_299),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_299),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_217),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_247),
.B(n_314),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_169),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_314),
.B(n_8),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_223),
.Y(n_407)
);

NAND2xp33_ASAP7_75t_R g408 ( 
.A(n_168),
.B(n_9),
.Y(n_408)
);

NOR2xp67_ASAP7_75t_L g409 ( 
.A(n_311),
.B(n_11),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_363),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_363),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_331),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_363),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_404),
.B(n_168),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_363),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_375),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_338),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_376),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_372),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_363),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_397),
.B(n_222),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_403),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_338),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_407),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_339),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_339),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_340),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_328),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_R g429 ( 
.A(n_340),
.B(n_230),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_334),
.B(n_176),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_337),
.B(n_306),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_342),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_345),
.B(n_209),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_342),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_356),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_350),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_335),
.B(n_176),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_341),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_341),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_358),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_343),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_371),
.B(n_264),
.Y(n_442)
);

NAND2x1_ASAP7_75t_L g443 ( 
.A(n_381),
.B(n_279),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_371),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_348),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_350),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_343),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_348),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_349),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_352),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_349),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_352),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_391),
.B(n_178),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_351),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_344),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_351),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_400),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_361),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_344),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_400),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_353),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_R g462 ( 
.A(n_353),
.B(n_246),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_346),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_346),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_347),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_328),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_347),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_360),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_364),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_329),
.B(n_311),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_362),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_379),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_330),
.B(n_264),
.Y(n_473)
);

INVx4_ASAP7_75t_SL g474 ( 
.A(n_332),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_365),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_367),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_355),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_366),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_368),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_359),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_R g481 ( 
.A(n_359),
.B(n_374),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_369),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_417),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_417),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_419),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_411),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_423),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_423),
.Y(n_488)
);

AND2x2_ASAP7_75t_SL g489 ( 
.A(n_431),
.B(n_354),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_421),
.B(n_397),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_411),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_414),
.B(n_406),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_425),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_431),
.B(n_357),
.Y(n_494)
);

AND3x2_ASAP7_75t_L g495 ( 
.A(n_428),
.B(n_239),
.C(n_224),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_414),
.B(n_374),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_473),
.B(n_333),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_453),
.B(n_378),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_419),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_425),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_453),
.A2(n_409),
.B1(n_336),
.B2(n_373),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_443),
.A2(n_239),
.B1(n_224),
.B2(n_386),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_427),
.B(n_378),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_426),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_442),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_473),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_411),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_470),
.B(n_401),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_412),
.A2(n_387),
.B1(n_383),
.B2(n_398),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_470),
.B(n_401),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_426),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_443),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_438),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_430),
.B(n_382),
.Y(n_514)
);

AO22x2_ASAP7_75t_L g515 ( 
.A1(n_433),
.A2(n_181),
.B1(n_242),
.B2(n_384),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_438),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_429),
.B(n_382),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_462),
.B(n_383),
.Y(n_518)
);

NAND2xp33_ASAP7_75t_L g519 ( 
.A(n_430),
.B(n_279),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_437),
.B(n_387),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_432),
.B(n_398),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_481),
.B(n_370),
.Y(n_522)
);

NOR2x1p5_ASAP7_75t_L g523 ( 
.A(n_434),
.B(n_174),
.Y(n_523)
);

INVx4_ASAP7_75t_SL g524 ( 
.A(n_411),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_439),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_439),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_441),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_412),
.A2(n_408),
.B1(n_395),
.B2(n_405),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_441),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_435),
.Y(n_530)
);

AND2x2_ASAP7_75t_SL g531 ( 
.A(n_480),
.B(n_279),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_442),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g533 ( 
.A(n_435),
.B(n_377),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_436),
.B(n_402),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_441),
.Y(n_535)
);

BUFx10_ASAP7_75t_L g536 ( 
.A(n_446),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_450),
.B(n_402),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_452),
.B(n_170),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_437),
.B(n_410),
.Y(n_539)
);

NOR2x1p5_ASAP7_75t_L g540 ( 
.A(n_461),
.B(n_174),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_468),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_442),
.B(n_463),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_410),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_447),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_447),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_410),
.Y(n_546)
);

AND2x6_ASAP7_75t_L g547 ( 
.A(n_442),
.B(n_279),
.Y(n_547)
);

OR2x6_ASAP7_75t_L g548 ( 
.A(n_480),
.B(n_380),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_474),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_463),
.B(n_465),
.Y(n_550)
);

INVxp67_ASAP7_75t_SL g551 ( 
.A(n_413),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_447),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_413),
.B(n_226),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_468),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_474),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_474),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_455),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_413),
.B(n_248),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_474),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_455),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_477),
.B(n_183),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_455),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_428),
.B(n_170),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_466),
.B(n_170),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_465),
.B(n_385),
.Y(n_565)
);

BUFx4f_ASAP7_75t_L g566 ( 
.A(n_471),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_416),
.Y(n_567)
);

INVxp67_ASAP7_75t_SL g568 ( 
.A(n_415),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_466),
.B(n_177),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_415),
.B(n_250),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_472),
.B(n_177),
.Y(n_571)
);

AND2x6_ASAP7_75t_L g572 ( 
.A(n_471),
.B(n_167),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_472),
.Y(n_573)
);

AO22x2_ASAP7_75t_L g574 ( 
.A1(n_433),
.A2(n_219),
.B1(n_321),
.B2(n_305),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_415),
.B(n_251),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_420),
.B(n_257),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_445),
.B(n_183),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_445),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_448),
.Y(n_579)
);

BUFx10_ASAP7_75t_L g580 ( 
.A(n_418),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_448),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_475),
.A2(n_186),
.B1(n_327),
.B2(n_185),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_475),
.A2(n_399),
.B1(n_396),
.B2(n_394),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_449),
.Y(n_584)
);

INVx1_ASAP7_75t_SL g585 ( 
.A(n_440),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_449),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_451),
.B(n_388),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_422),
.B(n_177),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_458),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_451),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_454),
.B(n_185),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_454),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_478),
.B(n_262),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_SL g594 ( 
.A(n_424),
.B(n_232),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_456),
.B(n_186),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_456),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_457),
.Y(n_597)
);

INVxp67_ASAP7_75t_SL g598 ( 
.A(n_457),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_460),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_460),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_482),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_478),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_478),
.B(n_266),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_459),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_479),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_479),
.B(n_389),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_459),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_479),
.A2(n_302),
.B1(n_327),
.B2(n_195),
.Y(n_608)
);

AND2x6_ASAP7_75t_L g609 ( 
.A(n_482),
.B(n_175),
.Y(n_609)
);

AND2x2_ASAP7_75t_SL g610 ( 
.A(n_482),
.B(n_180),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_444),
.B(n_390),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_464),
.B(n_269),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_464),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_464),
.A2(n_393),
.B1(n_392),
.B2(n_201),
.Y(n_614)
);

OAI22xp33_ASAP7_75t_SL g615 ( 
.A1(n_467),
.A2(n_193),
.B1(n_188),
.B2(n_182),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_467),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_467),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_469),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_476),
.A2(n_302),
.B1(n_195),
.B2(n_294),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_R g620 ( 
.A(n_481),
.B(n_187),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_417),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_473),
.B(n_326),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_431),
.B(n_189),
.Y(n_623)
);

NAND2xp33_ASAP7_75t_SL g624 ( 
.A(n_453),
.B(n_182),
.Y(n_624)
);

OR2x6_ASAP7_75t_L g625 ( 
.A(n_485),
.B(n_184),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_498),
.B(n_189),
.Y(n_626)
);

NOR2x1p5_ASAP7_75t_L g627 ( 
.A(n_496),
.B(n_188),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_487),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_485),
.B(n_306),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_531),
.B(n_194),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_567),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_492),
.B(n_198),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_531),
.A2(n_206),
.B1(n_212),
.B2(n_225),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_505),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_499),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_499),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_506),
.B(n_191),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_505),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_506),
.B(n_202),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_602),
.B(n_203),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_487),
.Y(n_641)
);

A2O1A1Ixp33_ASAP7_75t_L g642 ( 
.A1(n_623),
.A2(n_218),
.B(n_280),
.C(n_228),
.Y(n_642)
);

OAI221xp5_ASAP7_75t_L g643 ( 
.A1(n_624),
.A2(n_304),
.B1(n_237),
.B2(n_261),
.C(n_238),
.Y(n_643)
);

NAND3xp33_ASAP7_75t_L g644 ( 
.A(n_534),
.B(n_268),
.C(n_271),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_566),
.B(n_191),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_537),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_489),
.A2(n_290),
.B1(n_325),
.B2(n_288),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_514),
.B(n_192),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_602),
.B(n_244),
.Y(n_649)
);

OAI22xp33_ASAP7_75t_L g650 ( 
.A1(n_520),
.A2(n_259),
.B1(n_258),
.B2(n_256),
.Y(n_650)
);

A2O1A1Ixp33_ASAP7_75t_L g651 ( 
.A1(n_539),
.A2(n_272),
.B(n_282),
.C(n_320),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_598),
.B(n_273),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_493),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_573),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_601),
.B(n_318),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_601),
.B(n_319),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_533),
.B(n_193),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_497),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_605),
.B(n_192),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_489),
.A2(n_293),
.B1(n_292),
.B2(n_295),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_605),
.B(n_197),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_493),
.Y(n_662)
);

INVx8_ASAP7_75t_L g663 ( 
.A(n_548),
.Y(n_663)
);

AO22x1_ASAP7_75t_L g664 ( 
.A1(n_494),
.A2(n_309),
.B1(n_295),
.B2(n_303),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_542),
.B(n_197),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_532),
.B(n_294),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_622),
.B(n_306),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_542),
.B(n_310),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_610),
.A2(n_309),
.B1(n_293),
.B2(n_303),
.Y(n_669)
);

NAND2x1_ASAP7_75t_L g670 ( 
.A(n_549),
.B(n_80),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_578),
.B(n_584),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_511),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_586),
.B(n_310),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_566),
.B(n_297),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_596),
.B(n_297),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_597),
.B(n_599),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_511),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_622),
.B(n_277),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_490),
.B(n_307),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_600),
.B(n_312),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_548),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_497),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_561),
.B(n_533),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_579),
.B(n_307),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_532),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_525),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_566),
.B(n_312),
.Y(n_687)
);

INVx8_ASAP7_75t_L g688 ( 
.A(n_548),
.Y(n_688)
);

NAND2xp33_ASAP7_75t_SL g689 ( 
.A(n_620),
.B(n_296),
.Y(n_689)
);

A2O1A1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_624),
.A2(n_313),
.B(n_324),
.C(n_317),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_567),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_512),
.B(n_313),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_512),
.B(n_326),
.Y(n_693)
);

BUFx5_ASAP7_75t_L g694 ( 
.A(n_572),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_551),
.A2(n_278),
.B(n_281),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_501),
.A2(n_502),
.B1(n_610),
.B2(n_528),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_581),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_581),
.Y(n_698)
);

NAND3xp33_ASAP7_75t_L g699 ( 
.A(n_582),
.B(n_284),
.C(n_308),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_525),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_590),
.B(n_326),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_590),
.B(n_301),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_530),
.B(n_308),
.Y(n_703)
);

NAND2xp33_ASAP7_75t_L g704 ( 
.A(n_572),
.B(n_296),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_592),
.B(n_301),
.Y(n_705)
);

NAND2x1_ASAP7_75t_L g706 ( 
.A(n_549),
.B(n_56),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_526),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_550),
.A2(n_292),
.B1(n_301),
.B2(n_276),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_526),
.Y(n_709)
);

AO221x1_ASAP7_75t_L g710 ( 
.A1(n_574),
.A2(n_276),
.B1(n_13),
.B2(n_16),
.C(n_17),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_592),
.B(n_483),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_571),
.B(n_563),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_594),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_565),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_483),
.B(n_276),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_SL g716 ( 
.A(n_536),
.B(n_11),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_565),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_564),
.B(n_16),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_527),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_527),
.Y(n_720)
);

INVx4_ASAP7_75t_L g721 ( 
.A(n_617),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_529),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_550),
.Y(n_723)
);

OAI22xp33_ASAP7_75t_L g724 ( 
.A1(n_548),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_529),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_569),
.B(n_23),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_541),
.B(n_67),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_554),
.B(n_23),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_484),
.B(n_68),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_617),
.B(n_59),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_538),
.B(n_24),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_484),
.B(n_70),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_488),
.B(n_72),
.Y(n_733)
);

NOR2xp67_ASAP7_75t_L g734 ( 
.A(n_503),
.B(n_164),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_L g735 ( 
.A(n_572),
.B(n_54),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_508),
.B(n_25),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_606),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_508),
.B(n_25),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_618),
.Y(n_739)
);

NAND2x1_ASAP7_75t_L g740 ( 
.A(n_549),
.B(n_79),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_488),
.B(n_162),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_535),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_486),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_535),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_544),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_500),
.B(n_153),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_617),
.B(n_148),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_509),
.B(n_577),
.Y(n_748)
);

AO221x1_ASAP7_75t_L g749 ( 
.A1(n_574),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.C(n_32),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_606),
.Y(n_750)
);

INVxp67_ASAP7_75t_SL g751 ( 
.A(n_617),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_500),
.B(n_82),
.Y(n_752)
);

AND2x2_ASAP7_75t_SL g753 ( 
.A(n_519),
.B(n_139),
.Y(n_753)
);

AND2x2_ASAP7_75t_SL g754 ( 
.A(n_519),
.B(n_133),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_510),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_504),
.B(n_116),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_504),
.B(n_112),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_611),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_513),
.B(n_100),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_513),
.B(n_90),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_618),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_521),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_516),
.B(n_84),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_544),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_516),
.B(n_33),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_517),
.B(n_33),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_611),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_621),
.B(n_50),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_545),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_518),
.B(n_36),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_545),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_552),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_591),
.B(n_48),
.Y(n_773)
);

NAND2xp33_ASAP7_75t_L g774 ( 
.A(n_572),
.B(n_41),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_552),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_587),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_613),
.B(n_42),
.Y(n_777)
);

OR2x2_ASAP7_75t_SL g778 ( 
.A(n_574),
.B(n_515),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_557),
.Y(n_779)
);

O2A1O1Ixp5_ASAP7_75t_L g780 ( 
.A1(n_568),
.A2(n_44),
.B(n_46),
.C(n_48),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_557),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_617),
.B(n_46),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_613),
.B(n_612),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_585),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_553),
.B(n_593),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_603),
.B(n_595),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_L g787 ( 
.A1(n_619),
.A2(n_608),
.B1(n_576),
.B2(n_570),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_560),
.Y(n_788)
);

INVxp33_ASAP7_75t_L g789 ( 
.A(n_510),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_523),
.A2(n_540),
.B1(n_522),
.B2(n_587),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_495),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_786),
.B(n_587),
.Y(n_792)
);

O2A1O1Ixp33_ASAP7_75t_SL g793 ( 
.A1(n_630),
.A2(n_575),
.B(n_558),
.C(n_588),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_751),
.A2(n_785),
.B(n_721),
.Y(n_794)
);

O2A1O1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_632),
.A2(n_615),
.B(n_616),
.C(n_607),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_L g796 ( 
.A(n_694),
.B(n_743),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_683),
.B(n_604),
.Y(n_797)
);

O2A1O1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_630),
.A2(n_616),
.B(n_560),
.C(n_607),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_628),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_683),
.B(n_536),
.Y(n_800)
);

CKINVDCx10_ASAP7_75t_R g801 ( 
.A(n_625),
.Y(n_801)
);

NOR2xp67_ASAP7_75t_L g802 ( 
.A(n_636),
.B(n_604),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_646),
.B(n_762),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_641),
.Y(n_804)
);

BUFx2_ASAP7_75t_L g805 ( 
.A(n_635),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_748),
.A2(n_574),
.B1(n_614),
.B2(n_546),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_711),
.A2(n_556),
.B(n_559),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_787),
.A2(n_572),
.B1(n_609),
.B2(n_547),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_638),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_789),
.B(n_536),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_654),
.Y(n_811)
);

AOI21x1_ASAP7_75t_L g812 ( 
.A1(n_640),
.A2(n_562),
.B(n_524),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_638),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_685),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_755),
.Y(n_815)
);

BUFx12f_ASAP7_75t_L g816 ( 
.A(n_631),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_629),
.B(n_580),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_743),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_655),
.A2(n_555),
.B(n_559),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_696),
.B(n_580),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_656),
.A2(n_555),
.B(n_559),
.Y(n_821)
);

OAI21xp5_ASAP7_75t_L g822 ( 
.A1(n_723),
.A2(n_562),
.B(n_507),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_685),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_712),
.A2(n_692),
.B1(n_750),
.B2(n_737),
.Y(n_824)
);

AOI21x1_ASAP7_75t_L g825 ( 
.A1(n_649),
.A2(n_524),
.B(n_507),
.Y(n_825)
);

O2A1O1Ixp5_ASAP7_75t_L g826 ( 
.A1(n_639),
.A2(n_546),
.B(n_543),
.C(n_507),
.Y(n_826)
);

O2A1O1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_782),
.A2(n_546),
.B(n_543),
.C(n_583),
.Y(n_827)
);

NOR2x1_ASAP7_75t_L g828 ( 
.A(n_734),
.B(n_589),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_743),
.A2(n_556),
.B(n_486),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_671),
.A2(n_486),
.B(n_491),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_679),
.B(n_543),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_653),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_712),
.A2(n_609),
.B1(n_547),
.B2(n_515),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_676),
.A2(n_486),
.B(n_491),
.Y(n_834)
);

NOR2xp67_ASAP7_75t_L g835 ( 
.A(n_691),
.B(n_580),
.Y(n_835)
);

AOI21x1_ASAP7_75t_L g836 ( 
.A1(n_729),
.A2(n_524),
.B(n_491),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_713),
.B(n_491),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_658),
.B(n_524),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_766),
.A2(n_491),
.B(n_515),
.C(n_609),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_735),
.A2(n_547),
.B(n_609),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_659),
.A2(n_547),
.B(n_609),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_761),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_661),
.A2(n_652),
.B(n_732),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_682),
.B(n_547),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_784),
.Y(n_845)
);

NOR2x1p5_ASAP7_75t_SL g846 ( 
.A(n_694),
.B(n_547),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_714),
.B(n_609),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_662),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_733),
.A2(n_515),
.B(n_741),
.Y(n_849)
);

AOI21x1_ASAP7_75t_L g850 ( 
.A1(n_746),
.A2(n_756),
.B(n_752),
.Y(n_850)
);

O2A1O1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_782),
.A2(n_774),
.B(n_780),
.C(n_773),
.Y(n_851)
);

O2A1O1Ixp5_ASAP7_75t_L g852 ( 
.A1(n_672),
.A2(n_707),
.B(n_700),
.C(n_709),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_672),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_692),
.A2(n_776),
.B1(n_634),
.B2(n_717),
.Y(n_854)
);

OAI21x1_ASAP7_75t_L g855 ( 
.A1(n_719),
.A2(n_781),
.B(n_769),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_758),
.B(n_767),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_667),
.B(n_678),
.Y(n_857)
);

OAI321xp33_ASAP7_75t_L g858 ( 
.A1(n_708),
.A2(n_724),
.A3(n_643),
.B1(n_731),
.B2(n_718),
.C(n_726),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_657),
.B(n_625),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_757),
.A2(n_760),
.B(n_759),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_749),
.A2(n_710),
.B1(n_754),
.B2(n_753),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_R g862 ( 
.A(n_689),
.B(n_761),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_763),
.A2(n_686),
.B(n_700),
.Y(n_863)
);

NAND2x1p5_ASAP7_75t_L g864 ( 
.A(n_670),
.B(n_706),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_739),
.Y(n_865)
);

O2A1O1Ixp33_ASAP7_75t_SL g866 ( 
.A1(n_642),
.A2(n_727),
.B(n_651),
.C(n_730),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_677),
.A2(n_709),
.B(n_686),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_753),
.A2(n_754),
.B1(n_697),
.B2(n_698),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_791),
.B(n_666),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_684),
.B(n_665),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_677),
.A2(n_707),
.B(n_788),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_684),
.B(n_668),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_766),
.A2(n_770),
.B1(n_693),
.B2(n_674),
.Y(n_873)
);

INVx4_ASAP7_75t_L g874 ( 
.A(n_663),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_736),
.B(n_738),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_765),
.B(n_768),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_740),
.Y(n_877)
);

CKINVDCx8_ASAP7_75t_R g878 ( 
.A(n_663),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_L g879 ( 
.A1(n_633),
.A2(n_790),
.B1(n_687),
.B2(n_674),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_687),
.A2(n_730),
.B(n_747),
.Y(n_880)
);

NAND2x1p5_ASAP7_75t_L g881 ( 
.A(n_747),
.B(n_727),
.Y(n_881)
);

O2A1O1Ixp5_ASAP7_75t_L g882 ( 
.A1(n_777),
.A2(n_788),
.B(n_781),
.C(n_742),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_L g883 ( 
.A1(n_770),
.A2(n_693),
.B1(n_731),
.B2(n_645),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_720),
.A2(n_764),
.B(n_775),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_722),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_663),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_728),
.B(n_779),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_722),
.A2(n_764),
.B(n_775),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_666),
.B(n_681),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_725),
.A2(n_779),
.B(n_772),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_725),
.A2(n_742),
.B(n_772),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_744),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_701),
.B(n_702),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_728),
.B(n_771),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_718),
.A2(n_726),
.B(n_647),
.C(n_708),
.Y(n_895)
);

BUFx12f_ASAP7_75t_L g896 ( 
.A(n_625),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_745),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_769),
.B(n_771),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_705),
.B(n_715),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_703),
.B(n_680),
.Y(n_900)
);

O2A1O1Ixp5_ASAP7_75t_L g901 ( 
.A1(n_673),
.A2(n_675),
.B(n_650),
.C(n_637),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_644),
.B(n_694),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_704),
.A2(n_695),
.B(n_694),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_664),
.B(n_627),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_690),
.Y(n_905)
);

NOR2x1_ASAP7_75t_L g906 ( 
.A(n_699),
.B(n_716),
.Y(n_906)
);

BUFx4f_ASAP7_75t_L g907 ( 
.A(n_688),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_778),
.B(n_660),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_688),
.A2(n_694),
.B1(n_660),
.B2(n_669),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_688),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_669),
.A2(n_623),
.B(n_626),
.C(n_648),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_694),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_638),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_786),
.B(n_785),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_628),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_783),
.A2(n_751),
.B(n_512),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_785),
.A2(n_630),
.B(n_786),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_628),
.Y(n_918)
);

OA22x2_ASAP7_75t_L g919 ( 
.A1(n_749),
.A2(n_710),
.B1(n_748),
.B2(n_790),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_628),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_683),
.B(n_485),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_632),
.A2(n_630),
.B(n_696),
.C(n_492),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_786),
.B(n_785),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_646),
.B(n_683),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_786),
.B(n_785),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_786),
.B(n_785),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_628),
.Y(n_927)
);

O2A1O1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_632),
.A2(n_630),
.B(n_696),
.C(n_492),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_761),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_786),
.B(n_785),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_631),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_786),
.B(n_785),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_628),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_628),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_786),
.B(n_785),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_786),
.B(n_785),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_632),
.A2(n_630),
.B(n_696),
.C(n_492),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_646),
.B(n_683),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_628),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_L g940 ( 
.A1(n_749),
.A2(n_710),
.B1(n_754),
.B2(n_753),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_626),
.A2(n_623),
.B(n_648),
.C(n_683),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_SL g942 ( 
.A(n_631),
.B(n_691),
.Y(n_942)
);

O2A1O1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_632),
.A2(n_630),
.B(n_696),
.C(n_492),
.Y(n_943)
);

NOR3xp33_ASAP7_75t_L g944 ( 
.A(n_683),
.B(n_623),
.C(n_646),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_638),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_683),
.B(n_485),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_786),
.B(n_785),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_628),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_786),
.B(n_785),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_924),
.B(n_938),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_845),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_914),
.B(n_923),
.Y(n_952)
);

AO31x2_ASAP7_75t_L g953 ( 
.A1(n_839),
.A2(n_911),
.A3(n_849),
.B(n_879),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_799),
.Y(n_954)
);

OA22x2_ASAP7_75t_L g955 ( 
.A1(n_873),
.A2(n_883),
.B1(n_921),
.B2(n_946),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_925),
.B(n_926),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_811),
.Y(n_957)
);

INVx6_ASAP7_75t_L g958 ( 
.A(n_816),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_930),
.B(n_932),
.Y(n_959)
);

INVxp67_ASAP7_75t_L g960 ( 
.A(n_811),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_941),
.A2(n_935),
.B(n_949),
.C(n_947),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_936),
.B(n_944),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_924),
.B(n_938),
.Y(n_963)
);

OR2x2_ASAP7_75t_L g964 ( 
.A(n_805),
.B(n_944),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_804),
.Y(n_965)
);

INVx4_ASAP7_75t_L g966 ( 
.A(n_818),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_794),
.A2(n_796),
.B(n_860),
.Y(n_967)
);

AOI21x1_ASAP7_75t_L g968 ( 
.A1(n_836),
.A2(n_812),
.B(n_825),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_817),
.B(n_803),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_892),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_880),
.A2(n_843),
.B(n_916),
.Y(n_971)
);

AOI21xp33_ASAP7_75t_L g972 ( 
.A1(n_922),
.A2(n_937),
.B(n_928),
.Y(n_972)
);

AO22x1_ASAP7_75t_L g973 ( 
.A1(n_906),
.A2(n_803),
.B1(n_908),
.B2(n_865),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_792),
.B(n_870),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_922),
.A2(n_937),
.B(n_928),
.Y(n_975)
);

OAI21x1_ASAP7_75t_L g976 ( 
.A1(n_855),
.A2(n_863),
.B(n_852),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_895),
.A2(n_943),
.B(n_858),
.C(n_917),
.Y(n_977)
);

BUFx6f_ASAP7_75t_SL g978 ( 
.A(n_929),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_861),
.A2(n_940),
.B1(n_908),
.B2(n_909),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_872),
.B(n_875),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_874),
.B(n_910),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_857),
.B(n_859),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_818),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_874),
.B(n_886),
.Y(n_984)
);

OAI21x1_ASAP7_75t_L g985 ( 
.A1(n_852),
.A2(n_882),
.B(n_903),
.Y(n_985)
);

INVx4_ASAP7_75t_L g986 ( 
.A(n_818),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_900),
.B(n_797),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_900),
.B(n_824),
.Y(n_988)
);

OAI22x1_ASAP7_75t_L g989 ( 
.A1(n_833),
.A2(n_800),
.B1(n_820),
.B2(n_889),
.Y(n_989)
);

NOR2xp67_ASAP7_75t_L g990 ( 
.A(n_931),
.B(n_835),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_882),
.A2(n_871),
.B(n_890),
.Y(n_991)
);

OAI21x1_ASAP7_75t_L g992 ( 
.A1(n_867),
.A2(n_884),
.B(n_888),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_832),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_818),
.Y(n_994)
);

OAI21x1_ASAP7_75t_L g995 ( 
.A1(n_891),
.A2(n_826),
.B(n_830),
.Y(n_995)
);

OAI21x1_ASAP7_75t_L g996 ( 
.A1(n_826),
.A2(n_834),
.B(n_798),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_876),
.B(n_887),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_851),
.A2(n_901),
.B(n_905),
.C(n_795),
.Y(n_998)
);

AOI21xp33_ASAP7_75t_L g999 ( 
.A1(n_919),
.A2(n_795),
.B(n_861),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_892),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_842),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_856),
.B(n_837),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_869),
.Y(n_1003)
);

OAI21x1_ASAP7_75t_L g1004 ( 
.A1(n_864),
.A2(n_898),
.B(n_829),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_901),
.A2(n_854),
.B(n_940),
.C(n_868),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_810),
.B(n_815),
.Y(n_1006)
);

AO31x2_ASAP7_75t_L g1007 ( 
.A1(n_806),
.A2(n_894),
.A3(n_840),
.B(n_831),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_810),
.B(n_815),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_896),
.Y(n_1009)
);

AOI21x1_ASAP7_75t_L g1010 ( 
.A1(n_850),
.A2(n_902),
.B(n_893),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_899),
.A2(n_837),
.B(n_827),
.C(n_847),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_919),
.A2(n_822),
.B(n_827),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_809),
.B(n_813),
.Y(n_1013)
);

OAI22x1_ASAP7_75t_L g1014 ( 
.A1(n_889),
.A2(n_904),
.B1(n_869),
.B2(n_881),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_841),
.A2(n_821),
.B(n_819),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_942),
.B(n_862),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_848),
.B(n_915),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_912),
.A2(n_807),
.B(n_881),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_838),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_809),
.B(n_945),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_793),
.A2(n_866),
.B(n_844),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_877),
.A2(n_808),
.B(n_814),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_862),
.B(n_945),
.Y(n_1023)
);

AO31x2_ASAP7_75t_L g1024 ( 
.A1(n_918),
.A2(n_927),
.A3(n_920),
.B(n_885),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_907),
.Y(n_1025)
);

NAND2x1p5_ASAP7_75t_L g1026 ( 
.A(n_907),
.B(n_913),
.Y(n_1026)
);

AOI21xp33_ASAP7_75t_L g1027 ( 
.A1(n_853),
.A2(n_948),
.B(n_933),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_828),
.A2(n_846),
.B(n_934),
.C(n_939),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_802),
.A2(n_823),
.B(n_813),
.C(n_897),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_823),
.B(n_838),
.Y(n_1030)
);

INVx1_ASAP7_75t_SL g1031 ( 
.A(n_801),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_877),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_SL g1033 ( 
.A1(n_878),
.A2(n_489),
.B1(n_594),
.B2(n_431),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_924),
.B(n_485),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_914),
.B(n_932),
.Y(n_1035)
);

AND2x6_ASAP7_75t_L g1036 ( 
.A(n_909),
.B(n_808),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_SL g1037 ( 
.A1(n_911),
.A2(n_941),
.B(n_873),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_944),
.A2(n_919),
.B1(n_489),
.B2(n_908),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_924),
.B(n_938),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_924),
.B(n_485),
.Y(n_1040)
);

AOI21xp33_ASAP7_75t_L g1041 ( 
.A1(n_911),
.A2(n_928),
.B(n_922),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_914),
.A2(n_936),
.B(n_932),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_911),
.A2(n_941),
.B(n_914),
.C(n_925),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_914),
.A2(n_936),
.B(n_932),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_874),
.B(n_910),
.Y(n_1045)
);

AOI21xp33_ASAP7_75t_L g1046 ( 
.A1(n_911),
.A2(n_928),
.B(n_922),
.Y(n_1046)
);

AOI21x1_ASAP7_75t_L g1047 ( 
.A1(n_836),
.A2(n_812),
.B(n_825),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_911),
.A2(n_928),
.B(n_922),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_914),
.A2(n_923),
.B1(n_926),
.B2(n_925),
.Y(n_1049)
);

OAI21xp33_ASAP7_75t_L g1050 ( 
.A1(n_911),
.A2(n_908),
.B(n_941),
.Y(n_1050)
);

OAI21xp33_ASAP7_75t_SL g1051 ( 
.A1(n_914),
.A2(n_925),
.B(n_923),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_924),
.B(n_938),
.Y(n_1052)
);

O2A1O1Ixp5_ASAP7_75t_L g1053 ( 
.A1(n_941),
.A2(n_911),
.B(n_849),
.C(n_899),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_914),
.A2(n_936),
.B(n_932),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_914),
.B(n_932),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_818),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_892),
.Y(n_1057)
);

BUFx2_ASAP7_75t_SL g1058 ( 
.A(n_845),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_914),
.B(n_923),
.Y(n_1059)
);

OR2x6_ASAP7_75t_SL g1060 ( 
.A(n_931),
.B(n_631),
.Y(n_1060)
);

AO21x1_ASAP7_75t_L g1061 ( 
.A1(n_922),
.A2(n_937),
.B(n_928),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_855),
.A2(n_836),
.B(n_863),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_818),
.Y(n_1063)
);

CKINVDCx20_ASAP7_75t_R g1064 ( 
.A(n_931),
.Y(n_1064)
);

CKINVDCx6p67_ASAP7_75t_R g1065 ( 
.A(n_816),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_855),
.A2(n_836),
.B(n_863),
.Y(n_1066)
);

OAI21xp33_ASAP7_75t_L g1067 ( 
.A1(n_911),
.A2(n_908),
.B(n_941),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_931),
.Y(n_1068)
);

NAND2x1p5_ASAP7_75t_L g1069 ( 
.A(n_874),
.B(n_818),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_914),
.A2(n_923),
.B1(n_926),
.B2(n_925),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_914),
.B(n_923),
.Y(n_1071)
);

NAND3xp33_ASAP7_75t_SL g1072 ( 
.A(n_911),
.B(n_941),
.C(n_419),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_799),
.Y(n_1073)
);

AO31x2_ASAP7_75t_L g1074 ( 
.A1(n_839),
.A2(n_911),
.A3(n_849),
.B(n_879),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_855),
.A2(n_836),
.B(n_863),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_931),
.Y(n_1076)
);

CKINVDCx20_ASAP7_75t_R g1077 ( 
.A(n_931),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_914),
.B(n_932),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_924),
.B(n_485),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_874),
.B(n_910),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_892),
.Y(n_1081)
);

OAI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_911),
.A2(n_928),
.B(n_922),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_914),
.A2(n_936),
.B(n_932),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_1034),
.B(n_1040),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_954),
.Y(n_1085)
);

OA21x2_ASAP7_75t_L g1086 ( 
.A1(n_985),
.A2(n_1053),
.B(n_975),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_1072),
.A2(n_1067),
.B1(n_1050),
.B2(n_979),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_965),
.Y(n_1088)
);

AND2x2_ASAP7_75t_SL g1089 ( 
.A(n_1038),
.B(n_988),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_952),
.B(n_956),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_959),
.B(n_1035),
.Y(n_1091)
);

OR2x6_ASAP7_75t_L g1092 ( 
.A(n_1025),
.B(n_1058),
.Y(n_1092)
);

BUFx2_ASAP7_75t_SL g1093 ( 
.A(n_1064),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_1068),
.Y(n_1094)
);

OAI21xp33_ASAP7_75t_L g1095 ( 
.A1(n_950),
.A2(n_1052),
.B(n_1039),
.Y(n_1095)
);

AO21x1_ASAP7_75t_L g1096 ( 
.A1(n_1037),
.A2(n_979),
.B(n_1041),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1024),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_984),
.B(n_1025),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1083),
.A2(n_967),
.B(n_1051),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1079),
.B(n_969),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_1077),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_968),
.A2(n_1047),
.B(n_1066),
.Y(n_1102)
);

CKINVDCx8_ASAP7_75t_R g1103 ( 
.A(n_1076),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1055),
.A2(n_1078),
.B(n_1071),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_1001),
.Y(n_1105)
);

OR2x6_ASAP7_75t_L g1106 ( 
.A(n_1026),
.B(n_958),
.Y(n_1106)
);

INVx1_ASAP7_75t_SL g1107 ( 
.A(n_957),
.Y(n_1107)
);

NOR2x1_ASAP7_75t_L g1108 ( 
.A(n_990),
.B(n_1059),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_993),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1059),
.B(n_1071),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1050),
.A2(n_1067),
.B1(n_1033),
.B2(n_955),
.Y(n_1111)
);

INVx5_ASAP7_75t_L g1112 ( 
.A(n_983),
.Y(n_1112)
);

AOI21xp33_ASAP7_75t_L g1113 ( 
.A1(n_1037),
.A2(n_1082),
.B(n_1048),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1073),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_961),
.A2(n_971),
.B(n_1070),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1049),
.B(n_1070),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_1049),
.A2(n_963),
.B1(n_977),
.B2(n_1043),
.Y(n_1117)
);

OA21x2_ASAP7_75t_L g1118 ( 
.A1(n_975),
.A2(n_998),
.B(n_972),
.Y(n_1118)
);

NAND2x1p5_ASAP7_75t_L g1119 ( 
.A(n_966),
.B(n_986),
.Y(n_1119)
);

BUFx12f_ASAP7_75t_L g1120 ( 
.A(n_958),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_980),
.B(n_962),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_1036),
.A2(n_964),
.B1(n_982),
.B2(n_1082),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1006),
.A2(n_974),
.B1(n_973),
.B2(n_1008),
.Y(n_1123)
);

AO21x2_ASAP7_75t_L g1124 ( 
.A1(n_1041),
.A2(n_1046),
.B(n_972),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_SL g1125 ( 
.A1(n_957),
.A2(n_1048),
.B1(n_960),
.B2(n_1031),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_1065),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_997),
.B(n_987),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1017),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_1016),
.B(n_997),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1005),
.A2(n_1002),
.B1(n_1046),
.B2(n_999),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_984),
.B(n_981),
.Y(n_1131)
);

NAND2xp33_ASAP7_75t_L g1132 ( 
.A(n_1026),
.B(n_1023),
.Y(n_1132)
);

OR2x2_ASAP7_75t_L g1133 ( 
.A(n_951),
.B(n_1003),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1011),
.A2(n_1012),
.B(n_1021),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_999),
.A2(n_1012),
.B1(n_1022),
.B2(n_1017),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1030),
.B(n_981),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_970),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_1045),
.B(n_1080),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1061),
.B(n_1036),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1030),
.B(n_1080),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1000),
.Y(n_1141)
);

AND2x4_ASAP7_75t_L g1142 ( 
.A(n_1045),
.B(n_1019),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1057),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_983),
.Y(n_1144)
);

OR2x2_ASAP7_75t_L g1145 ( 
.A(n_1013),
.B(n_1020),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_1019),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1015),
.A2(n_1004),
.B(n_1018),
.Y(n_1147)
);

OAI21xp33_ASAP7_75t_L g1148 ( 
.A1(n_989),
.A2(n_1014),
.B(n_1028),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_1009),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_991),
.A2(n_992),
.B(n_995),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_978),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_983),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1081),
.B(n_1060),
.Y(n_1153)
);

OAI21xp33_ASAP7_75t_L g1154 ( 
.A1(n_1029),
.A2(n_1027),
.B(n_1010),
.Y(n_1154)
);

INVx5_ASAP7_75t_L g1155 ( 
.A(n_1056),
.Y(n_1155)
);

AO21x2_ASAP7_75t_L g1156 ( 
.A1(n_996),
.A2(n_976),
.B(n_1075),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1036),
.B(n_953),
.Y(n_1157)
);

INVxp67_ASAP7_75t_SL g1158 ( 
.A(n_1056),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1032),
.A2(n_1069),
.B1(n_1063),
.B2(n_1056),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_994),
.Y(n_1160)
);

INVx4_ASAP7_75t_L g1161 ( 
.A(n_978),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_1069),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1074),
.B(n_1031),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1062),
.Y(n_1164)
);

BUFx12f_ASAP7_75t_L g1165 ( 
.A(n_1027),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1007),
.Y(n_1166)
);

CKINVDCx8_ASAP7_75t_R g1167 ( 
.A(n_1007),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_984),
.B(n_1025),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_952),
.B(n_956),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_1025),
.Y(n_1170)
);

INVx1_ASAP7_75t_SL g1171 ( 
.A(n_957),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_954),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_952),
.B(n_956),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1034),
.B(n_1040),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1072),
.A2(n_944),
.B1(n_489),
.B2(n_1050),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_952),
.A2(n_1078),
.B1(n_959),
.B2(n_1035),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_952),
.B(n_956),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1025),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_952),
.B(n_1055),
.Y(n_1179)
);

NAND2x1p5_ASAP7_75t_L g1180 ( 
.A(n_966),
.B(n_874),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1042),
.A2(n_1054),
.B(n_1044),
.Y(n_1181)
);

BUFx2_ASAP7_75t_L g1182 ( 
.A(n_1001),
.Y(n_1182)
);

INVxp67_ASAP7_75t_SL g1183 ( 
.A(n_952),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_950),
.B(n_1039),
.Y(n_1184)
);

OR2x2_ASAP7_75t_L g1185 ( 
.A(n_980),
.B(n_485),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1042),
.A2(n_1054),
.B(n_1044),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_954),
.Y(n_1187)
);

INVx2_ASAP7_75t_SL g1188 ( 
.A(n_951),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1072),
.A2(n_944),
.B1(n_489),
.B2(n_1050),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_954),
.Y(n_1190)
);

CKINVDCx6p67_ASAP7_75t_R g1191 ( 
.A(n_1064),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_1064),
.Y(n_1192)
);

BUFx10_ASAP7_75t_L g1193 ( 
.A(n_1068),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_954),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_950),
.B(n_1039),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_1072),
.A2(n_944),
.B1(n_489),
.B2(n_1050),
.Y(n_1196)
);

AOI21xp33_ASAP7_75t_SL g1197 ( 
.A1(n_973),
.A2(n_691),
.B(n_631),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_SL g1198 ( 
.A1(n_961),
.A2(n_1043),
.B(n_1049),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1034),
.B(n_1040),
.Y(n_1199)
);

NAND3xp33_ASAP7_75t_SL g1200 ( 
.A(n_1033),
.B(n_911),
.C(n_941),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_1064),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_984),
.B(n_1025),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_952),
.B(n_1055),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_1064),
.Y(n_1204)
);

OR2x6_ASAP7_75t_L g1205 ( 
.A(n_1025),
.B(n_663),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_957),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_950),
.B(n_1039),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1034),
.B(n_1040),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1034),
.B(n_1040),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_954),
.Y(n_1210)
);

NAND3xp33_ASAP7_75t_L g1211 ( 
.A(n_1037),
.B(n_941),
.C(n_911),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_1146),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1200),
.A2(n_1089),
.B1(n_1207),
.B2(n_1184),
.Y(n_1213)
);

INVx6_ASAP7_75t_L g1214 ( 
.A(n_1112),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1085),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_1115),
.A2(n_1099),
.B(n_1150),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1195),
.A2(n_1095),
.B1(n_1211),
.B2(n_1096),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1111),
.B(n_1183),
.Y(n_1218)
);

BUFx2_ASAP7_75t_SL g1219 ( 
.A(n_1112),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1175),
.B(n_1189),
.Y(n_1220)
);

CKINVDCx11_ASAP7_75t_R g1221 ( 
.A(n_1103),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1095),
.A2(n_1211),
.B1(n_1196),
.B2(n_1125),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_1105),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1088),
.Y(n_1224)
);

INVx2_ASAP7_75t_SL g1225 ( 
.A(n_1155),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1125),
.A2(n_1113),
.B1(n_1121),
.B2(n_1087),
.Y(n_1226)
);

CKINVDCx6p67_ASAP7_75t_R g1227 ( 
.A(n_1120),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1122),
.B(n_1129),
.Y(n_1228)
);

BUFx12f_ASAP7_75t_L g1229 ( 
.A(n_1094),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_1191),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1155),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1113),
.A2(n_1163),
.B1(n_1117),
.B2(n_1176),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1157),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1102),
.A2(n_1181),
.B(n_1186),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1139),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1139),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1146),
.Y(n_1237)
);

NOR2x1_ASAP7_75t_R g1238 ( 
.A(n_1126),
.B(n_1093),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1123),
.A2(n_1108),
.B1(n_1176),
.B2(n_1179),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1104),
.A2(n_1117),
.B(n_1203),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1100),
.A2(n_1165),
.B1(n_1209),
.B2(n_1084),
.Y(n_1241)
);

CKINVDCx11_ASAP7_75t_R g1242 ( 
.A(n_1193),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1174),
.A2(n_1208),
.B1(n_1199),
.B2(n_1091),
.Y(n_1243)
);

AO21x1_ASAP7_75t_L g1244 ( 
.A1(n_1130),
.A2(n_1116),
.B(n_1134),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1109),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1114),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1182),
.Y(n_1247)
);

INVx2_ASAP7_75t_SL g1248 ( 
.A(n_1092),
.Y(n_1248)
);

BUFx2_ASAP7_75t_R g1249 ( 
.A(n_1101),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1185),
.B(n_1090),
.Y(n_1250)
);

INVx1_ASAP7_75t_SL g1251 ( 
.A(n_1107),
.Y(n_1251)
);

BUFx2_ASAP7_75t_R g1252 ( 
.A(n_1192),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1138),
.B(n_1142),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1172),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1206),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1187),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_1131),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1148),
.A2(n_1169),
.B1(n_1090),
.B2(n_1177),
.Y(n_1258)
);

AO21x2_ASAP7_75t_L g1259 ( 
.A1(n_1148),
.A2(n_1154),
.B(n_1156),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1190),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1169),
.A2(n_1177),
.B1(n_1173),
.B2(n_1124),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1166),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1194),
.Y(n_1263)
);

INVx4_ASAP7_75t_SL g1264 ( 
.A(n_1106),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_SL g1265 ( 
.A1(n_1173),
.A2(n_1110),
.B1(n_1153),
.B2(n_1127),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1127),
.B(n_1128),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1118),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1132),
.A2(n_1140),
.B1(n_1136),
.B2(n_1151),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_1193),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1124),
.A2(n_1135),
.B1(n_1171),
.B2(n_1161),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1086),
.Y(n_1271)
);

AO21x1_ASAP7_75t_L g1272 ( 
.A1(n_1198),
.A2(n_1145),
.B(n_1159),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1154),
.A2(n_1210),
.B(n_1162),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1171),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1137),
.Y(n_1275)
);

CKINVDCx6p67_ASAP7_75t_R g1276 ( 
.A(n_1092),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1141),
.B(n_1143),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_SL g1278 ( 
.A1(n_1161),
.A2(n_1204),
.B1(n_1201),
.B2(n_1106),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1142),
.B(n_1160),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1156),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1158),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1144),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1138),
.A2(n_1106),
.B1(n_1197),
.B2(n_1167),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1164),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1119),
.Y(n_1285)
);

INVx3_ASAP7_75t_L g1286 ( 
.A(n_1119),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1131),
.A2(n_1133),
.B1(n_1149),
.B2(n_1092),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1205),
.A2(n_1188),
.B1(n_1098),
.B2(n_1202),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1180),
.A2(n_1205),
.B(n_1168),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1152),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_1202),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1152),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1152),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1170),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1178),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1178),
.A2(n_1200),
.B1(n_489),
.B2(n_1089),
.Y(n_1296)
);

INVx3_ASAP7_75t_L g1297 ( 
.A(n_1146),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1094),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1200),
.A2(n_489),
.B1(n_1089),
.B2(n_1072),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1200),
.A2(n_489),
.B1(n_1089),
.B2(n_1072),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1138),
.B(n_1142),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1094),
.Y(n_1302)
);

AOI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1184),
.A2(n_345),
.B1(n_361),
.B2(n_358),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1112),
.Y(n_1304)
);

AO21x2_ASAP7_75t_L g1305 ( 
.A1(n_1147),
.A2(n_1082),
.B(n_1048),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1097),
.Y(n_1306)
);

OAI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1184),
.A2(n_716),
.B1(n_431),
.B2(n_594),
.Y(n_1307)
);

NAND2x1p5_ASAP7_75t_L g1308 ( 
.A(n_1118),
.B(n_1097),
.Y(n_1308)
);

OA21x2_ASAP7_75t_L g1309 ( 
.A1(n_1115),
.A2(n_1082),
.B(n_1048),
.Y(n_1309)
);

BUFx12f_ASAP7_75t_L g1310 ( 
.A(n_1094),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1111),
.B(n_1089),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1200),
.A2(n_489),
.B1(n_1089),
.B2(n_1072),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_1105),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1274),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1306),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1250),
.B(n_1266),
.Y(n_1316)
);

AO31x2_ASAP7_75t_L g1317 ( 
.A1(n_1244),
.A2(n_1267),
.A3(n_1271),
.B(n_1280),
.Y(n_1317)
);

OR2x6_ASAP7_75t_L g1318 ( 
.A(n_1240),
.B(n_1234),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1213),
.B(n_1265),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1255),
.Y(n_1320)
);

INVxp33_ASAP7_75t_L g1321 ( 
.A(n_1303),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1266),
.B(n_1258),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1255),
.Y(n_1323)
);

BUFx4_ASAP7_75t_R g1324 ( 
.A(n_1257),
.Y(n_1324)
);

NAND2x1p5_ASAP7_75t_L g1325 ( 
.A(n_1309),
.B(n_1273),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1239),
.B(n_1307),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1262),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1273),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_1214),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_1251),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1217),
.B(n_1218),
.Y(n_1331)
);

BUFx2_ASAP7_75t_L g1332 ( 
.A(n_1233),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1233),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1235),
.B(n_1236),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_SL g1335 ( 
.A1(n_1309),
.A2(n_1304),
.B(n_1231),
.Y(n_1335)
);

INVx5_ASAP7_75t_SL g1336 ( 
.A(n_1276),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1284),
.B(n_1264),
.Y(n_1337)
);

OA21x2_ASAP7_75t_L g1338 ( 
.A1(n_1244),
.A2(n_1232),
.B(n_1261),
.Y(n_1338)
);

BUFx4f_ASAP7_75t_L g1339 ( 
.A(n_1276),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1281),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1254),
.Y(n_1341)
);

AO21x2_ASAP7_75t_L g1342 ( 
.A1(n_1305),
.A2(n_1259),
.B(n_1272),
.Y(n_1342)
);

AO21x2_ASAP7_75t_L g1343 ( 
.A1(n_1305),
.A2(n_1259),
.B(n_1272),
.Y(n_1343)
);

INVx2_ASAP7_75t_SL g1344 ( 
.A(n_1214),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1260),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1220),
.B(n_1228),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1263),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1308),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1309),
.B(n_1270),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1259),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1216),
.A2(n_1312),
.B(n_1299),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1263),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1214),
.Y(n_1353)
);

AO21x2_ASAP7_75t_L g1354 ( 
.A1(n_1220),
.A2(n_1256),
.B(n_1224),
.Y(n_1354)
);

INVxp67_ASAP7_75t_L g1355 ( 
.A(n_1223),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1264),
.B(n_1212),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1218),
.B(n_1228),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1222),
.B(n_1226),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1215),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1245),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1246),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1311),
.B(n_1300),
.Y(n_1362)
);

AOI21xp33_ASAP7_75t_L g1363 ( 
.A1(n_1296),
.A2(n_1311),
.B(n_1241),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1216),
.B(n_1243),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1275),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1277),
.Y(n_1366)
);

AO21x2_ASAP7_75t_L g1367 ( 
.A1(n_1268),
.A2(n_1285),
.B(n_1283),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1277),
.B(n_1279),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1237),
.B(n_1297),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_1221),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1317),
.B(n_1342),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1317),
.B(n_1292),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1317),
.B(n_1292),
.Y(n_1373)
);

BUFx3_ASAP7_75t_L g1374 ( 
.A(n_1337),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1354),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1315),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1317),
.B(n_1293),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1317),
.B(n_1293),
.Y(n_1378)
);

INVx4_ASAP7_75t_SL g1379 ( 
.A(n_1356),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1354),
.B(n_1313),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1342),
.B(n_1295),
.Y(n_1381)
);

INVx4_ASAP7_75t_L g1382 ( 
.A(n_1324),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1354),
.B(n_1313),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1343),
.B(n_1282),
.Y(n_1384)
);

NOR2x1_ASAP7_75t_L g1385 ( 
.A(n_1335),
.B(n_1219),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1343),
.B(n_1290),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1349),
.B(n_1294),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1349),
.B(n_1325),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1364),
.B(n_1247),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1334),
.B(n_1278),
.Y(n_1390)
);

INVx2_ASAP7_75t_R g1391 ( 
.A(n_1350),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1325),
.B(n_1294),
.Y(n_1392)
);

INVxp67_ASAP7_75t_L g1393 ( 
.A(n_1320),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1326),
.B(n_1286),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1364),
.B(n_1223),
.Y(n_1395)
);

INVx2_ASAP7_75t_SL g1396 ( 
.A(n_1328),
.Y(n_1396)
);

NAND2x1_ASAP7_75t_L g1397 ( 
.A(n_1335),
.B(n_1214),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_1319),
.B(n_1288),
.Y(n_1398)
);

INVxp67_ASAP7_75t_SL g1399 ( 
.A(n_1341),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1358),
.A2(n_1242),
.B1(n_1253),
.B2(n_1301),
.Y(n_1400)
);

OAI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1358),
.A2(n_1248),
.B1(n_1269),
.B2(n_1257),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1382),
.A2(n_1321),
.B1(n_1331),
.B2(n_1339),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1387),
.B(n_1348),
.Y(n_1403)
);

NAND3xp33_ASAP7_75t_L g1404 ( 
.A(n_1398),
.B(n_1351),
.C(n_1363),
.Y(n_1404)
);

AOI21xp33_ASAP7_75t_L g1405 ( 
.A1(n_1398),
.A2(n_1322),
.B(n_1367),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1393),
.B(n_1314),
.Y(n_1406)
);

OAI221xp5_ASAP7_75t_L g1407 ( 
.A1(n_1400),
.A2(n_1287),
.B1(n_1355),
.B2(n_1316),
.C(n_1339),
.Y(n_1407)
);

OAI21xp5_ASAP7_75t_SL g1408 ( 
.A1(n_1400),
.A2(n_1362),
.B(n_1346),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1382),
.A2(n_1362),
.B1(n_1367),
.B2(n_1338),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1389),
.B(n_1327),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_SL g1411 ( 
.A1(n_1382),
.A2(n_1338),
.B(n_1356),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1388),
.B(n_1327),
.Y(n_1412)
);

NOR2x1_ASAP7_75t_SL g1413 ( 
.A(n_1382),
.B(n_1328),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1389),
.B(n_1340),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1388),
.B(n_1392),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1376),
.Y(n_1416)
);

OAI221xp5_ASAP7_75t_L g1417 ( 
.A1(n_1394),
.A2(n_1339),
.B1(n_1330),
.B2(n_1357),
.C(n_1289),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1388),
.B(n_1368),
.Y(n_1418)
);

NAND3xp33_ASAP7_75t_L g1419 ( 
.A(n_1394),
.B(n_1338),
.C(n_1323),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1382),
.A2(n_1339),
.B1(n_1357),
.B2(n_1336),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1395),
.B(n_1345),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1392),
.B(n_1368),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1395),
.B(n_1347),
.Y(n_1423)
);

OAI21xp33_ASAP7_75t_L g1424 ( 
.A1(n_1390),
.A2(n_1318),
.B(n_1366),
.Y(n_1424)
);

NOR3xp33_ASAP7_75t_L g1425 ( 
.A(n_1401),
.B(n_1385),
.C(n_1397),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1390),
.A2(n_1336),
.B1(n_1269),
.B2(n_1338),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1376),
.Y(n_1427)
);

AOI221xp5_ASAP7_75t_L g1428 ( 
.A1(n_1401),
.A2(n_1366),
.B1(n_1361),
.B2(n_1359),
.C(n_1360),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1392),
.B(n_1372),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1372),
.B(n_1373),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1385),
.A2(n_1336),
.B1(n_1230),
.B2(n_1291),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1399),
.B(n_1352),
.Y(n_1432)
);

NAND3xp33_ASAP7_75t_L g1433 ( 
.A(n_1380),
.B(n_1318),
.C(n_1361),
.Y(n_1433)
);

NAND4xp25_ASAP7_75t_L g1434 ( 
.A(n_1380),
.B(n_1359),
.C(n_1360),
.D(n_1365),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1399),
.B(n_1365),
.Y(n_1435)
);

OAI221xp5_ASAP7_75t_L g1436 ( 
.A1(n_1397),
.A2(n_1318),
.B1(n_1329),
.B2(n_1344),
.C(n_1353),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1372),
.B(n_1332),
.Y(n_1437)
);

NAND3xp33_ASAP7_75t_L g1438 ( 
.A(n_1380),
.B(n_1318),
.C(n_1369),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1383),
.B(n_1332),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1383),
.B(n_1333),
.Y(n_1440)
);

NAND3xp33_ASAP7_75t_L g1441 ( 
.A(n_1383),
.B(n_1386),
.C(n_1384),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1430),
.B(n_1391),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1441),
.B(n_1371),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1416),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1430),
.B(n_1391),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1416),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1427),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1439),
.B(n_1384),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1427),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1435),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1440),
.B(n_1386),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1429),
.B(n_1391),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1429),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1403),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1415),
.B(n_1371),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1422),
.Y(n_1456)
);

NOR2xp67_ASAP7_75t_L g1457 ( 
.A(n_1419),
.B(n_1375),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1437),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1413),
.B(n_1396),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1421),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1414),
.B(n_1371),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1418),
.B(n_1373),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1418),
.B(n_1373),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1412),
.B(n_1377),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1423),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1424),
.B(n_1377),
.Y(n_1466)
);

INVxp67_ASAP7_75t_L g1467 ( 
.A(n_1410),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1411),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1432),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1434),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1419),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1424),
.B(n_1378),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1453),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1455),
.B(n_1413),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1461),
.B(n_1406),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1455),
.B(n_1462),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1453),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1453),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1446),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1455),
.B(n_1411),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1446),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1444),
.Y(n_1482)
);

NAND3xp33_ASAP7_75t_L g1483 ( 
.A(n_1471),
.B(n_1404),
.C(n_1405),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1467),
.B(n_1370),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1444),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1444),
.Y(n_1486)
);

INVxp67_ASAP7_75t_L g1487 ( 
.A(n_1470),
.Y(n_1487)
);

INVx2_ASAP7_75t_SL g1488 ( 
.A(n_1459),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1471),
.B(n_1378),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1447),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1468),
.B(n_1379),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1471),
.B(n_1378),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1447),
.Y(n_1493)
);

OR2x6_ASAP7_75t_L g1494 ( 
.A(n_1468),
.B(n_1397),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1467),
.B(n_1230),
.Y(n_1495)
);

INVxp67_ASAP7_75t_L g1496 ( 
.A(n_1470),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1447),
.Y(n_1497)
);

INVxp67_ASAP7_75t_L g1498 ( 
.A(n_1470),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1449),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1469),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1453),
.Y(n_1501)
);

NOR5xp2_ASAP7_75t_L g1502 ( 
.A(n_1450),
.B(n_1436),
.C(n_1433),
.D(n_1438),
.E(n_1417),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1462),
.B(n_1374),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1460),
.B(n_1229),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1449),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1449),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1468),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1454),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1462),
.B(n_1374),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1450),
.B(n_1381),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1482),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1505),
.Y(n_1512)
);

INVx1_ASAP7_75t_SL g1513 ( 
.A(n_1484),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1489),
.B(n_1443),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1480),
.B(n_1463),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1487),
.Y(n_1516)
);

NOR2x1_ASAP7_75t_L g1517 ( 
.A(n_1483),
.B(n_1457),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1482),
.Y(n_1518)
);

INVxp67_ASAP7_75t_L g1519 ( 
.A(n_1495),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1496),
.B(n_1469),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1485),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1483),
.A2(n_1425),
.B1(n_1402),
.B2(n_1426),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1504),
.B(n_1229),
.Y(n_1523)
);

NAND2x1p5_ASAP7_75t_L g1524 ( 
.A(n_1507),
.B(n_1457),
.Y(n_1524)
);

NAND2x1_ASAP7_75t_L g1525 ( 
.A(n_1480),
.B(n_1468),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1485),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1505),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1486),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1498),
.A2(n_1409),
.B1(n_1457),
.B2(n_1443),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1474),
.B(n_1463),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1486),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1474),
.B(n_1463),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1476),
.B(n_1442),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1475),
.B(n_1469),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1475),
.B(n_1469),
.Y(n_1535)
);

AOI322xp5_ASAP7_75t_L g1536 ( 
.A1(n_1489),
.A2(n_1472),
.A3(n_1466),
.B1(n_1442),
.B2(n_1445),
.C1(n_1458),
.C2(n_1464),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1507),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1491),
.Y(n_1538)
);

INVx2_ASAP7_75t_SL g1539 ( 
.A(n_1491),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1491),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1490),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1490),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1492),
.B(n_1443),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1492),
.B(n_1461),
.Y(n_1544)
);

NOR2x1p5_ASAP7_75t_L g1545 ( 
.A(n_1491),
.B(n_1227),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1510),
.B(n_1310),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_1503),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1510),
.B(n_1469),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1493),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1505),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1506),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1476),
.B(n_1503),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1473),
.B(n_1461),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1511),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1511),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1522),
.A2(n_1517),
.B1(n_1519),
.B2(n_1529),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1515),
.B(n_1488),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1515),
.B(n_1488),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1513),
.B(n_1310),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1545),
.B(n_1494),
.Y(n_1560)
);

INVx1_ASAP7_75t_SL g1561 ( 
.A(n_1516),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1546),
.A2(n_1431),
.B1(n_1420),
.B2(n_1494),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1526),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1526),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1541),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1514),
.B(n_1473),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1541),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1540),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1514),
.B(n_1473),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1523),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1540),
.B(n_1509),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1518),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1521),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1540),
.B(n_1552),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1538),
.B(n_1298),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1552),
.B(n_1509),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1537),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1528),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1520),
.B(n_1469),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1531),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1524),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1530),
.B(n_1532),
.Y(n_1582)
);

OR2x6_ASAP7_75t_L g1583 ( 
.A(n_1524),
.B(n_1494),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1543),
.B(n_1477),
.Y(n_1584)
);

NOR2x1_ASAP7_75t_L g1585 ( 
.A(n_1525),
.B(n_1479),
.Y(n_1585)
);

OR2x6_ASAP7_75t_L g1586 ( 
.A(n_1524),
.B(n_1494),
.Y(n_1586)
);

AOI222xp33_ASAP7_75t_L g1587 ( 
.A1(n_1547),
.A2(n_1472),
.B1(n_1466),
.B2(n_1408),
.C1(n_1502),
.C2(n_1428),
.Y(n_1587)
);

BUFx3_ASAP7_75t_L g1588 ( 
.A(n_1538),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1530),
.B(n_1532),
.Y(n_1589)
);

OAI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1587),
.A2(n_1525),
.B(n_1536),
.Y(n_1590)
);

NAND4xp25_ASAP7_75t_L g1591 ( 
.A(n_1556),
.B(n_1502),
.C(n_1543),
.D(n_1535),
.Y(n_1591)
);

AOI21xp33_ASAP7_75t_L g1592 ( 
.A1(n_1561),
.A2(n_1539),
.B(n_1494),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1588),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1555),
.Y(n_1594)
);

AOI21xp33_ASAP7_75t_SL g1595 ( 
.A1(n_1559),
.A2(n_1539),
.B(n_1302),
.Y(n_1595)
);

AOI222xp33_ASAP7_75t_L g1596 ( 
.A1(n_1577),
.A2(n_1570),
.B1(n_1574),
.B2(n_1568),
.C1(n_1562),
.C2(n_1588),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1555),
.Y(n_1597)
);

OAI221xp5_ASAP7_75t_SL g1598 ( 
.A1(n_1583),
.A2(n_1544),
.B1(n_1466),
.B2(n_1472),
.C(n_1407),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1563),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1563),
.Y(n_1600)
);

AOI322xp5_ASAP7_75t_L g1601 ( 
.A1(n_1585),
.A2(n_1442),
.A3(n_1445),
.B1(n_1533),
.B2(n_1534),
.C1(n_1548),
.C2(n_1458),
.Y(n_1601)
);

AOI221xp5_ASAP7_75t_L g1602 ( 
.A1(n_1572),
.A2(n_1549),
.B1(n_1542),
.B2(n_1450),
.C(n_1550),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1570),
.B(n_1298),
.Y(n_1603)
);

INVxp67_ASAP7_75t_L g1604 ( 
.A(n_1575),
.Y(n_1604)
);

OAI31xp33_ASAP7_75t_L g1605 ( 
.A1(n_1560),
.A2(n_1544),
.A3(n_1500),
.B(n_1533),
.Y(n_1605)
);

AOI32xp33_ASAP7_75t_L g1606 ( 
.A1(n_1574),
.A2(n_1445),
.A3(n_1452),
.B1(n_1481),
.B2(n_1479),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1579),
.B(n_1553),
.Y(n_1607)
);

AOI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1560),
.A2(n_1459),
.B1(n_1465),
.B2(n_1460),
.Y(n_1608)
);

AND3x2_ASAP7_75t_L g1609 ( 
.A(n_1581),
.B(n_1227),
.C(n_1238),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1564),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_SL g1611 ( 
.A(n_1560),
.B(n_1581),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1576),
.B(n_1460),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1576),
.B(n_1456),
.Y(n_1613)
);

OAI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1583),
.A2(n_1458),
.B1(n_1451),
.B2(n_1448),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1582),
.B(n_1456),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1593),
.B(n_1582),
.Y(n_1616)
);

INVxp67_ASAP7_75t_L g1617 ( 
.A(n_1603),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1596),
.B(n_1589),
.Y(n_1618)
);

NAND2xp33_ASAP7_75t_L g1619 ( 
.A(n_1590),
.B(n_1302),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1594),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1597),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1599),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1604),
.B(n_1589),
.Y(n_1623)
);

INVxp67_ASAP7_75t_L g1624 ( 
.A(n_1611),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1604),
.B(n_1571),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1612),
.B(n_1573),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1600),
.Y(n_1627)
);

AND2x4_ASAP7_75t_L g1628 ( 
.A(n_1609),
.B(n_1583),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1609),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1595),
.B(n_1571),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1610),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1607),
.Y(n_1632)
);

AND2x4_ASAP7_75t_L g1633 ( 
.A(n_1615),
.B(n_1583),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1613),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1605),
.B(n_1578),
.Y(n_1635)
);

AOI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1619),
.A2(n_1591),
.B1(n_1598),
.B2(n_1606),
.C(n_1592),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_L g1637 ( 
.A(n_1617),
.B(n_1598),
.Y(n_1637)
);

AOI21xp33_ASAP7_75t_L g1638 ( 
.A1(n_1619),
.A2(n_1586),
.B(n_1580),
.Y(n_1638)
);

AOI221xp5_ASAP7_75t_L g1639 ( 
.A1(n_1624),
.A2(n_1602),
.B1(n_1614),
.B2(n_1580),
.C(n_1565),
.Y(n_1639)
);

AOI211xp5_ASAP7_75t_L g1640 ( 
.A1(n_1618),
.A2(n_1635),
.B(n_1629),
.C(n_1628),
.Y(n_1640)
);

AOI211xp5_ASAP7_75t_SL g1641 ( 
.A1(n_1628),
.A2(n_1608),
.B(n_1565),
.C(n_1567),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1616),
.B(n_1601),
.Y(n_1642)
);

XNOR2xp5_ASAP7_75t_L g1643 ( 
.A(n_1616),
.B(n_1586),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1623),
.B(n_1557),
.Y(n_1644)
);

AOI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1630),
.A2(n_1586),
.B(n_1554),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1625),
.B(n_1557),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1630),
.A2(n_1586),
.B(n_1567),
.Y(n_1647)
);

AOI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1632),
.A2(n_1564),
.B(n_1558),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1643),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1646),
.Y(n_1650)
);

AOI211xp5_ASAP7_75t_L g1651 ( 
.A1(n_1636),
.A2(n_1628),
.B(n_1625),
.C(n_1621),
.Y(n_1651)
);

AOI22x1_ASAP7_75t_L g1652 ( 
.A1(n_1641),
.A2(n_1633),
.B1(n_1627),
.B2(n_1620),
.Y(n_1652)
);

NOR2x1_ASAP7_75t_L g1653 ( 
.A(n_1637),
.B(n_1627),
.Y(n_1653)
);

NOR3xp33_ASAP7_75t_L g1654 ( 
.A(n_1640),
.B(n_1631),
.C(n_1622),
.Y(n_1654)
);

NOR3x1_ASAP7_75t_L g1655 ( 
.A(n_1642),
.B(n_1626),
.C(n_1634),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1648),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_SL g1657 ( 
.A1(n_1647),
.A2(n_1633),
.B(n_1626),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1644),
.Y(n_1658)
);

NOR3xp33_ASAP7_75t_L g1659 ( 
.A(n_1638),
.B(n_1633),
.C(n_1569),
.Y(n_1659)
);

NOR4xp25_ASAP7_75t_L g1660 ( 
.A(n_1656),
.B(n_1639),
.C(n_1645),
.D(n_1566),
.Y(n_1660)
);

OAI211xp5_ASAP7_75t_SL g1661 ( 
.A1(n_1651),
.A2(n_1657),
.B(n_1653),
.C(n_1658),
.Y(n_1661)
);

NAND3xp33_ASAP7_75t_L g1662 ( 
.A(n_1652),
.B(n_1569),
.C(n_1566),
.Y(n_1662)
);

NOR2x1p5_ASAP7_75t_L g1663 ( 
.A(n_1650),
.B(n_1584),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1654),
.B(n_1558),
.Y(n_1664)
);

AOI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1661),
.A2(n_1659),
.B1(n_1654),
.B2(n_1649),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1663),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1664),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1662),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1660),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1663),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1666),
.B(n_1655),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1665),
.B(n_1584),
.Y(n_1672)
);

NOR3xp33_ASAP7_75t_L g1673 ( 
.A(n_1670),
.B(n_1252),
.C(n_1249),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1668),
.Y(n_1674)
);

NOR2x1_ASAP7_75t_L g1675 ( 
.A(n_1669),
.B(n_1512),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1671),
.A2(n_1667),
.B1(n_1551),
.B2(n_1512),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1672),
.Y(n_1677)
);

NAND4xp75_ASAP7_75t_L g1678 ( 
.A(n_1674),
.B(n_1675),
.C(n_1673),
.D(n_1225),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1677),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1679),
.A2(n_1676),
.B1(n_1678),
.B2(n_1550),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1680),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1680),
.Y(n_1682)
);

OR2x4_ASAP7_75t_L g1683 ( 
.A(n_1682),
.B(n_1231),
.Y(n_1683)
);

OAI21x1_ASAP7_75t_L g1684 ( 
.A1(n_1682),
.A2(n_1551),
.B(n_1527),
.Y(n_1684)
);

AOI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1683),
.A2(n_1681),
.B1(n_1527),
.B2(n_1481),
.Y(n_1685)
);

AOI221xp5_ASAP7_75t_L g1686 ( 
.A1(n_1684),
.A2(n_1553),
.B1(n_1499),
.B2(n_1497),
.C(n_1493),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1685),
.A2(n_1478),
.B1(n_1477),
.B2(n_1501),
.Y(n_1687)
);

AOI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1687),
.A2(n_1686),
.B1(n_1477),
.B2(n_1478),
.Y(n_1688)
);

AOI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1688),
.A2(n_1497),
.B1(n_1499),
.B2(n_1506),
.C(n_1508),
.Y(n_1689)
);

AOI211xp5_ASAP7_75t_L g1690 ( 
.A1(n_1689),
.A2(n_1231),
.B(n_1304),
.C(n_1225),
.Y(n_1690)
);


endmodule