module real_aes_7998_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_725;
wire n_504;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g108 ( .A(n_0), .Y(n_108) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_1), .A2(n_144), .B(n_147), .C(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g210 ( .A(n_2), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_3), .A2(n_139), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_4), .B(n_220), .Y(n_533) );
AOI21xp33_ASAP7_75t_L g221 ( .A1(n_5), .A2(n_139), .B(n_222), .Y(n_221) );
AND2x6_ASAP7_75t_L g144 ( .A(n_6), .B(n_145), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_7), .A2(n_190), .B(n_191), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_8), .B(n_41), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_8), .B(n_41), .Y(n_124) );
OAI22xp5_ASAP7_75t_L g127 ( .A1(n_9), .A2(n_31), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_9), .Y(n_129) );
INVx1_ASAP7_75t_L g468 ( .A(n_10), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_11), .B(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g227 ( .A(n_12), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_13), .B(n_180), .Y(n_489) );
INVx1_ASAP7_75t_L g165 ( .A(n_14), .Y(n_165) );
INVx1_ASAP7_75t_L g198 ( .A(n_15), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_16), .A2(n_153), .B(n_199), .C(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_17), .B(n_220), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_18), .B(n_155), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_19), .B(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_20), .B(n_569), .Y(n_568) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_21), .A2(n_179), .B(n_213), .C(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_22), .B(n_220), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_23), .B(n_180), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_24), .A2(n_195), .B(n_197), .C(n_199), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_25), .B(n_180), .Y(n_508) );
CKINVDCx16_ASAP7_75t_R g518 ( .A(n_26), .Y(n_518) );
INVx1_ASAP7_75t_L g507 ( .A(n_27), .Y(n_507) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_28), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_29), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_30), .B(n_180), .Y(n_211) );
INVx1_ASAP7_75t_L g128 ( .A(n_31), .Y(n_128) );
INVx1_ASAP7_75t_L g565 ( .A(n_32), .Y(n_565) );
INVx1_ASAP7_75t_L g237 ( .A(n_33), .Y(n_237) );
INVx2_ASAP7_75t_L g142 ( .A(n_34), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_35), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_36), .A2(n_179), .B(n_228), .C(n_531), .Y(n_530) );
INVxp67_ASAP7_75t_L g566 ( .A(n_37), .Y(n_566) );
A2O1A1Ixp33_ASAP7_75t_L g146 ( .A1(n_38), .A2(n_144), .B(n_147), .C(n_150), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_39), .A2(n_147), .B(n_506), .C(n_511), .Y(n_505) );
CKINVDCx14_ASAP7_75t_R g529 ( .A(n_40), .Y(n_529) );
INVx1_ASAP7_75t_L g235 ( .A(n_42), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g466 ( .A1(n_43), .A2(n_157), .B(n_225), .C(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_44), .B(n_180), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_45), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_46), .Y(n_562) );
INVx1_ASAP7_75t_L g496 ( .A(n_47), .Y(n_496) );
CKINVDCx16_ASAP7_75t_R g238 ( .A(n_48), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_49), .B(n_139), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_50), .Y(n_125) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_51), .A2(n_147), .B1(n_213), .B2(n_234), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_52), .Y(n_167) );
CKINVDCx16_ASAP7_75t_R g206 ( .A(n_53), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_54), .A2(n_225), .B(n_226), .C(n_228), .Y(n_224) );
CKINVDCx14_ASAP7_75t_R g465 ( .A(n_55), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_56), .Y(n_275) );
INVx1_ASAP7_75t_L g223 ( .A(n_57), .Y(n_223) );
INVx1_ASAP7_75t_L g145 ( .A(n_58), .Y(n_145) );
INVx1_ASAP7_75t_L g164 ( .A(n_59), .Y(n_164) );
INVx1_ASAP7_75t_SL g532 ( .A(n_60), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_61), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_62), .B(n_220), .Y(n_500) );
INVx1_ASAP7_75t_L g521 ( .A(n_63), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_SL g245 ( .A1(n_64), .A2(n_155), .B(n_228), .C(n_246), .Y(n_245) );
INVxp67_ASAP7_75t_L g247 ( .A(n_65), .Y(n_247) );
INVx1_ASAP7_75t_L g112 ( .A(n_66), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_67), .A2(n_139), .B(n_464), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_68), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_69), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_70), .A2(n_139), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g268 ( .A(n_71), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_72), .A2(n_190), .B(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g475 ( .A(n_73), .Y(n_475) );
CKINVDCx16_ASAP7_75t_R g504 ( .A(n_74), .Y(n_504) );
OAI22xp5_ASAP7_75t_SL g737 ( .A1(n_75), .A2(n_76), .B1(n_738), .B2(n_739), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_75), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_76), .Y(n_738) );
A2O1A1Ixp33_ASAP7_75t_L g269 ( .A1(n_77), .A2(n_144), .B(n_147), .C(n_270), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_78), .A2(n_139), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g478 ( .A(n_79), .Y(n_478) );
AOI222xp33_ASAP7_75t_SL g126 ( .A1(n_80), .A2(n_127), .B1(n_130), .B2(n_726), .C1(n_727), .C2(n_731), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_81), .B(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g162 ( .A(n_82), .Y(n_162) );
INVx1_ASAP7_75t_L g487 ( .A(n_83), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_84), .B(n_155), .Y(n_154) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_85), .A2(n_102), .B1(n_113), .B2(n_741), .Y(n_101) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_86), .A2(n_144), .B(n_147), .C(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g109 ( .A(n_87), .Y(n_109) );
OR2x2_ASAP7_75t_L g121 ( .A(n_87), .B(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g725 ( .A(n_87), .B(n_123), .Y(n_725) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_88), .A2(n_147), .B(n_520), .C(n_523), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_89), .B(n_173), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_90), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g175 ( .A1(n_91), .A2(n_144), .B(n_147), .C(n_176), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_92), .Y(n_185) );
INVx1_ASAP7_75t_L g244 ( .A(n_93), .Y(n_244) );
CKINVDCx16_ASAP7_75t_R g192 ( .A(n_94), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_95), .B(n_152), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_96), .B(n_169), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_97), .B(n_169), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_98), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_99), .A2(n_139), .B(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g499 ( .A(n_100), .Y(n_499) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
CKINVDCx9p33_ASAP7_75t_R g742 ( .A(n_103), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx14_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_109), .C(n_110), .Y(n_107) );
AND2x2_ASAP7_75t_L g123 ( .A(n_108), .B(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g455 ( .A(n_109), .B(n_123), .Y(n_455) );
NOR2x2_ASAP7_75t_L g733 ( .A(n_109), .B(n_122), .Y(n_733) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AOI22x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_126), .B1(n_734), .B2(n_735), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_119), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_SL g734 ( .A(n_116), .Y(n_734) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_119), .A2(n_736), .B(n_740), .Y(n_735) );
NOR2xp33_ASAP7_75t_SL g119 ( .A(n_120), .B(n_125), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_121), .Y(n_740) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g726 ( .A(n_127), .Y(n_726) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_455), .B1(n_456), .B2(n_725), .Y(n_130) );
INVx2_ASAP7_75t_L g728 ( .A(n_131), .Y(n_728) );
AND2x2_ASAP7_75t_SL g131 ( .A(n_132), .B(n_424), .Y(n_131) );
NOR3xp33_ASAP7_75t_L g132 ( .A(n_133), .B(n_317), .C(n_390), .Y(n_132) );
OAI211xp5_ASAP7_75t_SL g133 ( .A1(n_134), .A2(n_202), .B(n_249), .C(n_301), .Y(n_133) );
INVxp67_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_170), .Y(n_135) );
AND2x2_ASAP7_75t_L g265 ( .A(n_136), .B(n_266), .Y(n_265) );
INVx3_ASAP7_75t_L g284 ( .A(n_136), .Y(n_284) );
INVx2_ASAP7_75t_L g299 ( .A(n_136), .Y(n_299) );
INVx1_ASAP7_75t_L g329 ( .A(n_136), .Y(n_329) );
AND2x2_ASAP7_75t_L g379 ( .A(n_136), .B(n_300), .Y(n_379) );
AOI32xp33_ASAP7_75t_L g406 ( .A1(n_136), .A2(n_334), .A3(n_407), .B1(n_409), .B2(n_410), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_136), .B(n_255), .Y(n_412) );
AND2x2_ASAP7_75t_L g439 ( .A(n_136), .B(n_282), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_136), .B(n_448), .Y(n_447) );
OR2x6_ASAP7_75t_L g136 ( .A(n_137), .B(n_166), .Y(n_136) );
AOI21xp5_ASAP7_75t_SL g137 ( .A1(n_138), .A2(n_146), .B(n_159), .Y(n_137) );
BUFx2_ASAP7_75t_L g190 ( .A(n_139), .Y(n_190) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_144), .Y(n_139) );
NAND2x1p5_ASAP7_75t_L g207 ( .A(n_140), .B(n_144), .Y(n_207) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
INVx1_ASAP7_75t_L g510 ( .A(n_141), .Y(n_510) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g148 ( .A(n_142), .Y(n_148) );
INVx1_ASAP7_75t_L g214 ( .A(n_142), .Y(n_214) );
INVx1_ASAP7_75t_L g149 ( .A(n_143), .Y(n_149) );
INVx3_ASAP7_75t_L g153 ( .A(n_143), .Y(n_153) );
INVx1_ASAP7_75t_L g155 ( .A(n_143), .Y(n_155) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_143), .Y(n_180) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_143), .Y(n_196) );
INVx4_ASAP7_75t_SL g200 ( .A(n_144), .Y(n_200) );
BUFx3_ASAP7_75t_L g511 ( .A(n_144), .Y(n_511) );
INVx5_ASAP7_75t_L g193 ( .A(n_147), .Y(n_193) );
AND2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
BUFx3_ASAP7_75t_L g158 ( .A(n_148), .Y(n_158) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_148), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_154), .B(n_156), .Y(n_150) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_152), .A2(n_210), .B(n_211), .C(n_212), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_L g506 ( .A1(n_152), .A2(n_507), .B(n_508), .C(n_509), .Y(n_506) );
OAI22xp33_ASAP7_75t_L g564 ( .A1(n_152), .A2(n_195), .B1(n_565), .B2(n_566), .Y(n_564) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_153), .B(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_153), .B(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_153), .B(n_468), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_156), .A2(n_271), .B(n_272), .Y(n_270) );
O2A1O1Ixp5_ASAP7_75t_L g486 ( .A1(n_156), .A2(n_487), .B(n_488), .C(n_489), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_L g520 ( .A1(n_156), .A2(n_488), .B(n_521), .C(n_522), .Y(n_520) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g199 ( .A(n_158), .Y(n_199) );
INVx1_ASAP7_75t_L g273 ( .A(n_159), .Y(n_273) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_160), .A2(n_205), .B(n_215), .Y(n_204) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_160), .A2(n_232), .B(n_239), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_160), .B(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_161), .Y(n_169) );
AND2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
AND2x2_ASAP7_75t_SL g173 ( .A(n_162), .B(n_163), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
NOR2xp33_ASAP7_75t_SL g166 ( .A(n_167), .B(n_168), .Y(n_166) );
INVx3_ASAP7_75t_L g220 ( .A(n_168), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_168), .B(n_491), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_168), .B(n_513), .Y(n_512) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_168), .A2(n_517), .B(n_524), .Y(n_516) );
INVx4_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_169), .A2(n_242), .B(n_248), .Y(n_241) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_169), .Y(n_472) );
AND2x2_ASAP7_75t_L g328 ( .A(n_170), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g350 ( .A(n_170), .Y(n_350) );
AND2x2_ASAP7_75t_L g435 ( .A(n_170), .B(n_265), .Y(n_435) );
AND2x2_ASAP7_75t_L g438 ( .A(n_170), .B(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_187), .Y(n_170) );
INVx2_ASAP7_75t_L g257 ( .A(n_171), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_171), .B(n_282), .Y(n_288) );
AND2x2_ASAP7_75t_L g298 ( .A(n_171), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g334 ( .A(n_171), .Y(n_334) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_174), .B(n_184), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_172), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g569 ( .A(n_172), .Y(n_569) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g186 ( .A(n_173), .Y(n_186) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_173), .A2(n_189), .B(n_201), .Y(n_188) );
OA21x2_ASAP7_75t_L g462 ( .A1(n_173), .A2(n_463), .B(n_469), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_L g503 ( .A1(n_173), .A2(n_207), .B(n_504), .C(n_505), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_175), .B(n_183), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_181), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_179), .B(n_532), .Y(n_531) );
INVx4_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g225 ( .A(n_180), .Y(n_225) );
HB1xp67_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx3_ASAP7_75t_L g228 ( .A(n_182), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_186), .B(n_216), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_186), .B(n_275), .Y(n_274) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_186), .A2(n_483), .B(n_490), .Y(n_482) );
AND2x2_ASAP7_75t_L g276 ( .A(n_187), .B(n_257), .Y(n_276) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g258 ( .A(n_188), .Y(n_258) );
AND2x2_ASAP7_75t_L g300 ( .A(n_188), .B(n_282), .Y(n_300) );
AND2x2_ASAP7_75t_L g369 ( .A(n_188), .B(n_266), .Y(n_369) );
O2A1O1Ixp33_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_194), .C(n_200), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_193), .A2(n_200), .B(n_223), .C(n_224), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_193), .A2(n_200), .B(n_244), .C(n_245), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_SL g464 ( .A1(n_193), .A2(n_200), .B(n_465), .C(n_466), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_SL g474 ( .A1(n_193), .A2(n_200), .B(n_475), .C(n_476), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_SL g495 ( .A1(n_193), .A2(n_200), .B(n_496), .C(n_497), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_193), .A2(n_200), .B(n_529), .C(n_530), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_SL g561 ( .A1(n_193), .A2(n_200), .B(n_562), .C(n_563), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_195), .B(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_195), .B(n_478), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_195), .B(n_499), .Y(n_498) );
INVx4_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
OAI22xp5_ASAP7_75t_SL g234 ( .A1(n_196), .A2(n_235), .B1(n_236), .B2(n_237), .Y(n_234) );
INVx2_ASAP7_75t_L g236 ( .A(n_196), .Y(n_236) );
OAI22xp33_ASAP7_75t_L g232 ( .A1(n_200), .A2(n_207), .B1(n_233), .B2(n_238), .Y(n_232) );
INVx1_ASAP7_75t_L g523 ( .A(n_200), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_203), .B(n_217), .Y(n_202) );
OR2x2_ASAP7_75t_L g263 ( .A(n_203), .B(n_231), .Y(n_263) );
INVx1_ASAP7_75t_L g342 ( .A(n_203), .Y(n_342) );
AND2x2_ASAP7_75t_L g356 ( .A(n_203), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_203), .B(n_230), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_203), .B(n_354), .Y(n_408) );
AND2x2_ASAP7_75t_L g416 ( .A(n_203), .B(n_417), .Y(n_416) );
INVx3_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx3_ASAP7_75t_L g253 ( .A(n_204), .Y(n_253) );
AND2x2_ASAP7_75t_L g323 ( .A(n_204), .B(n_231), .Y(n_323) );
OAI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_208), .Y(n_205) );
OAI21xp5_ASAP7_75t_L g267 ( .A1(n_207), .A2(n_268), .B(n_269), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g483 ( .A1(n_207), .A2(n_484), .B(n_485), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g517 ( .A1(n_207), .A2(n_518), .B(n_519), .Y(n_517) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx3_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_217), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g450 ( .A(n_217), .Y(n_450) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_230), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_218), .B(n_294), .Y(n_316) );
OR2x2_ASAP7_75t_L g345 ( .A(n_218), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g377 ( .A(n_218), .B(n_357), .Y(n_377) );
INVx1_ASAP7_75t_SL g397 ( .A(n_218), .Y(n_397) );
AND2x2_ASAP7_75t_L g401 ( .A(n_218), .B(n_262), .Y(n_401) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_SL g254 ( .A(n_219), .B(n_230), .Y(n_254) );
AND2x2_ASAP7_75t_L g261 ( .A(n_219), .B(n_241), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_219), .B(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g304 ( .A(n_219), .B(n_286), .Y(n_304) );
INVx1_ASAP7_75t_SL g311 ( .A(n_219), .Y(n_311) );
BUFx2_ASAP7_75t_L g322 ( .A(n_219), .Y(n_322) );
AND2x2_ASAP7_75t_L g338 ( .A(n_219), .B(n_253), .Y(n_338) );
AND2x2_ASAP7_75t_L g353 ( .A(n_219), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g417 ( .A(n_219), .B(n_231), .Y(n_417) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_229), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_230), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g341 ( .A(n_230), .B(n_342), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g358 ( .A1(n_230), .A2(n_359), .B1(n_362), .B2(n_365), .C(n_370), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_230), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_241), .Y(n_230) );
INVx3_ASAP7_75t_L g286 ( .A(n_231), .Y(n_286) );
INVx2_ASAP7_75t_L g488 ( .A(n_236), .Y(n_488) );
BUFx2_ASAP7_75t_L g296 ( .A(n_241), .Y(n_296) );
AND2x2_ASAP7_75t_L g310 ( .A(n_241), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g327 ( .A(n_241), .Y(n_327) );
OR2x2_ASAP7_75t_L g346 ( .A(n_241), .B(n_286), .Y(n_346) );
INVx3_ASAP7_75t_L g354 ( .A(n_241), .Y(n_354) );
AND2x2_ASAP7_75t_L g357 ( .A(n_241), .B(n_286), .Y(n_357) );
AOI221xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_255), .B1(n_259), .B2(n_264), .C(n_277), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_252), .B(n_326), .Y(n_451) );
OR2x2_ASAP7_75t_L g454 ( .A(n_252), .B(n_285), .Y(n_454) );
INVx1_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
OAI221xp5_ASAP7_75t_SL g277 ( .A1(n_253), .A2(n_278), .B1(n_285), .B2(n_287), .C(n_290), .Y(n_277) );
AND2x2_ASAP7_75t_L g294 ( .A(n_253), .B(n_286), .Y(n_294) );
AND2x2_ASAP7_75t_L g302 ( .A(n_253), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_253), .B(n_310), .Y(n_309) );
NAND2x1_ASAP7_75t_L g352 ( .A(n_253), .B(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g404 ( .A(n_253), .B(n_346), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g392 ( .A1(n_255), .A2(n_364), .B1(n_393), .B2(n_395), .Y(n_392) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AOI322xp5_ASAP7_75t_L g301 ( .A1(n_256), .A2(n_265), .A3(n_302), .B1(n_305), .B2(n_308), .C1(n_312), .C2(n_315), .Y(n_301) );
OR2x2_ASAP7_75t_L g313 ( .A(n_256), .B(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_257), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g292 ( .A(n_257), .B(n_266), .Y(n_292) );
INVx1_ASAP7_75t_L g307 ( .A(n_257), .Y(n_307) );
AND2x2_ASAP7_75t_L g373 ( .A(n_257), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g283 ( .A(n_258), .B(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g374 ( .A(n_258), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_258), .B(n_282), .Y(n_448) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_262), .B(n_397), .Y(n_396) );
INVx3_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g348 ( .A(n_263), .B(n_295), .Y(n_348) );
OR2x2_ASAP7_75t_L g445 ( .A(n_263), .B(n_296), .Y(n_445) );
INVx1_ASAP7_75t_L g426 ( .A(n_264), .Y(n_426) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_276), .Y(n_264) );
INVx4_ASAP7_75t_L g314 ( .A(n_265), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_265), .B(n_333), .Y(n_339) );
INVx2_ASAP7_75t_L g282 ( .A(n_266), .Y(n_282) );
AO21x2_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_273), .B(n_274), .Y(n_266) );
AO21x2_ASAP7_75t_L g558 ( .A1(n_273), .A2(n_559), .B(n_567), .Y(n_558) );
INVx1_ASAP7_75t_L g576 ( .A(n_273), .Y(n_576) );
INVx1_ASAP7_75t_L g364 ( .A(n_276), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_276), .B(n_336), .Y(n_405) );
AOI21xp33_ASAP7_75t_L g351 ( .A1(n_278), .A2(n_352), .B(n_355), .Y(n_351) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g336 ( .A(n_282), .Y(n_336) );
INVx1_ASAP7_75t_L g363 ( .A(n_282), .Y(n_363) );
INVx1_ASAP7_75t_L g289 ( .A(n_283), .Y(n_289) );
AND2x2_ASAP7_75t_L g291 ( .A(n_283), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g387 ( .A(n_284), .B(n_373), .Y(n_387) );
AND2x2_ASAP7_75t_L g409 ( .A(n_284), .B(n_369), .Y(n_409) );
BUFx2_ASAP7_75t_L g361 ( .A(n_286), .Y(n_361) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
AOI32xp33_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_293), .A3(n_294), .B1(n_295), .B2(n_297), .Y(n_290) );
INVx1_ASAP7_75t_L g371 ( .A(n_291), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_291), .A2(n_419), .B1(n_420), .B2(n_422), .Y(n_418) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_294), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_294), .B(n_353), .Y(n_394) );
AND2x2_ASAP7_75t_L g441 ( .A(n_294), .B(n_326), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_295), .B(n_342), .Y(n_389) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g442 ( .A(n_297), .Y(n_442) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
INVx1_ASAP7_75t_L g367 ( .A(n_298), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_300), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g414 ( .A(n_300), .B(n_334), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_300), .B(n_329), .Y(n_421) );
INVx1_ASAP7_75t_SL g403 ( .A(n_302), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_303), .B(n_354), .Y(n_381) );
NOR4xp25_ASAP7_75t_L g427 ( .A(n_303), .B(n_326), .C(n_428), .D(n_431), .Y(n_427) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_304), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVxp67_ASAP7_75t_L g384 ( .A(n_307), .Y(n_384) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OAI21xp33_ASAP7_75t_L g434 ( .A1(n_310), .A2(n_401), .B(n_435), .Y(n_434) );
AND2x4_ASAP7_75t_L g326 ( .A(n_311), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g375 ( .A(n_314), .Y(n_375) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND4xp25_ASAP7_75t_SL g317 ( .A(n_318), .B(n_343), .C(n_358), .D(n_378), .Y(n_317) );
O2A1O1Ixp33_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_324), .B(n_328), .C(n_330), .Y(n_318) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
INVx1_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g410 ( .A(n_323), .B(n_353), .Y(n_410) );
AND2x2_ASAP7_75t_L g419 ( .A(n_323), .B(n_397), .Y(n_419) );
INVx3_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_326), .B(n_361), .Y(n_423) );
AND2x2_ASAP7_75t_L g335 ( .A(n_329), .B(n_336), .Y(n_335) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_337), .B1(n_339), .B2(n_340), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
AND2x2_ASAP7_75t_L g433 ( .A(n_333), .B(n_379), .Y(n_433) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_335), .B(n_384), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_336), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
O2A1O1Ixp33_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_347), .B(n_349), .C(n_351), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g378 ( .A1(n_344), .A2(n_379), .B1(n_380), .B2(n_382), .C(n_385), .Y(n_378) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OAI221xp5_ASAP7_75t_L g436 ( .A1(n_352), .A2(n_437), .B1(n_440), .B2(n_442), .C(n_443), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_353), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_361), .B(n_430), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx1_ASAP7_75t_L g391 ( .A(n_363), .Y(n_391) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_366), .A2(n_386), .B1(n_388), .B2(n_389), .Y(n_385) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AOI21xp33_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_372), .B(n_376), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_375), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI221xp5_ASAP7_75t_L g449 ( .A1(n_386), .A2(n_412), .B1(n_450), .B2(n_451), .C(n_452), .Y(n_449) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g431 ( .A(n_388), .Y(n_431) );
OAI211xp5_ASAP7_75t_SL g390 ( .A1(n_391), .A2(n_392), .B(n_398), .C(n_418), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AOI211xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_401), .B(n_402), .C(n_411), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
A2O1A1Ixp33_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_404), .B(n_405), .C(n_406), .Y(n_402) );
INVx1_ASAP7_75t_L g430 ( .A(n_408), .Y(n_430) );
OAI21xp5_ASAP7_75t_SL g452 ( .A1(n_409), .A2(n_435), .B(n_453), .Y(n_452) );
AOI21xp33_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_413), .B(n_415), .Y(n_411) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVxp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OAI21xp5_ASAP7_75t_SL g444 ( .A1(n_421), .A2(n_445), .B(n_446), .Y(n_444) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NOR3xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_436), .C(n_449), .Y(n_424) );
OAI211xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .B(n_432), .C(n_434), .Y(n_425) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
CKINVDCx14_ASAP7_75t_R g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g730 ( .A(n_455), .Y(n_730) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OAI22xp5_ASAP7_75t_SL g727 ( .A1(n_457), .A2(n_725), .B1(n_728), .B2(n_729), .Y(n_727) );
XOR2xp5_ASAP7_75t_L g736 ( .A(n_457), .B(n_737), .Y(n_736) );
OR2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_655), .Y(n_457) );
NAND5xp2_ASAP7_75t_L g458 ( .A(n_459), .B(n_570), .C(n_602), .D(n_619), .E(n_642), .Y(n_458) );
AOI221xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_501), .B1(n_534), .B2(n_538), .C(n_542), .Y(n_459) );
INVx1_ASAP7_75t_L g682 ( .A(n_460), .Y(n_682) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_480), .Y(n_460) );
AND3x2_ASAP7_75t_L g657 ( .A(n_461), .B(n_482), .C(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_470), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_462), .B(n_540), .Y(n_539) );
BUFx3_ASAP7_75t_L g549 ( .A(n_462), .Y(n_549) );
AND2x2_ASAP7_75t_L g553 ( .A(n_462), .B(n_492), .Y(n_553) );
INVx2_ASAP7_75t_L g579 ( .A(n_462), .Y(n_579) );
OR2x2_ASAP7_75t_L g590 ( .A(n_462), .B(n_493), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_462), .B(n_481), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_462), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g669 ( .A(n_462), .B(n_493), .Y(n_669) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_470), .Y(n_552) );
AND2x2_ASAP7_75t_L g610 ( .A(n_470), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_470), .B(n_481), .Y(n_629) );
INVx1_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
OR2x2_ASAP7_75t_L g541 ( .A(n_471), .B(n_481), .Y(n_541) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_471), .Y(n_548) );
AND2x2_ASAP7_75t_L g596 ( .A(n_471), .B(n_493), .Y(n_596) );
NAND3xp33_ASAP7_75t_L g621 ( .A(n_471), .B(n_480), .C(n_579), .Y(n_621) );
AND2x2_ASAP7_75t_L g686 ( .A(n_471), .B(n_482), .Y(n_686) );
AND2x2_ASAP7_75t_L g720 ( .A(n_471), .B(n_481), .Y(n_720) );
OA21x2_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B(n_479), .Y(n_471) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_472), .A2(n_494), .B(n_500), .Y(n_493) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_472), .A2(n_527), .B(n_533), .Y(n_526) );
INVxp67_ASAP7_75t_L g550 ( .A(n_480), .Y(n_550) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_492), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_481), .B(n_579), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_481), .B(n_610), .Y(n_618) );
AND2x2_ASAP7_75t_L g668 ( .A(n_481), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g696 ( .A(n_481), .Y(n_696) );
INVx4_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g603 ( .A(n_482), .B(n_596), .Y(n_603) );
BUFx3_ASAP7_75t_L g635 ( .A(n_482), .Y(n_635) );
INVx2_ASAP7_75t_L g611 ( .A(n_492), .Y(n_611) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_493), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_501), .A2(n_671), .B1(n_673), .B2(n_674), .Y(n_670) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_514), .Y(n_501) );
AND2x2_ASAP7_75t_L g534 ( .A(n_502), .B(n_535), .Y(n_534) );
INVx3_ASAP7_75t_SL g545 ( .A(n_502), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_502), .B(n_574), .Y(n_606) );
OR2x2_ASAP7_75t_L g625 ( .A(n_502), .B(n_515), .Y(n_625) );
AND2x2_ASAP7_75t_L g630 ( .A(n_502), .B(n_582), .Y(n_630) );
AND2x2_ASAP7_75t_L g633 ( .A(n_502), .B(n_575), .Y(n_633) );
AND2x2_ASAP7_75t_L g645 ( .A(n_502), .B(n_526), .Y(n_645) );
AND2x2_ASAP7_75t_L g661 ( .A(n_502), .B(n_516), .Y(n_661) );
AND2x4_ASAP7_75t_L g664 ( .A(n_502), .B(n_536), .Y(n_664) );
OR2x2_ASAP7_75t_L g681 ( .A(n_502), .B(n_617), .Y(n_681) );
OR2x2_ASAP7_75t_L g712 ( .A(n_502), .B(n_558), .Y(n_712) );
NAND2xp5_ASAP7_75t_SL g714 ( .A(n_502), .B(n_640), .Y(n_714) );
OR2x6_ASAP7_75t_L g502 ( .A(n_503), .B(n_512), .Y(n_502) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_510), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g588 ( .A(n_514), .B(n_556), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_514), .B(n_575), .Y(n_707) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_526), .Y(n_514) );
AND2x2_ASAP7_75t_L g544 ( .A(n_515), .B(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g574 ( .A(n_515), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g582 ( .A(n_515), .B(n_558), .Y(n_582) );
AND2x2_ASAP7_75t_L g600 ( .A(n_515), .B(n_536), .Y(n_600) );
OR2x2_ASAP7_75t_L g617 ( .A(n_515), .B(n_575), .Y(n_617) );
INVx2_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
BUFx2_ASAP7_75t_L g537 ( .A(n_516), .Y(n_537) );
AND2x2_ASAP7_75t_L g640 ( .A(n_516), .B(n_526), .Y(n_640) );
INVx2_ASAP7_75t_L g536 ( .A(n_526), .Y(n_536) );
INVx1_ASAP7_75t_L g652 ( .A(n_526), .Y(n_652) );
AND2x2_ASAP7_75t_L g702 ( .A(n_526), .B(n_545), .Y(n_702) );
AND2x2_ASAP7_75t_L g555 ( .A(n_535), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g586 ( .A(n_535), .B(n_545), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_535), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
AND2x2_ASAP7_75t_L g573 ( .A(n_536), .B(n_545), .Y(n_573) );
OR2x2_ASAP7_75t_L g689 ( .A(n_537), .B(n_663), .Y(n_689) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_540), .B(n_669), .Y(n_675) );
INVx2_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
OAI32xp33_ASAP7_75t_L g631 ( .A1(n_541), .A2(n_632), .A3(n_634), .B1(n_636), .B2(n_637), .Y(n_631) );
OR2x2_ASAP7_75t_L g648 ( .A(n_541), .B(n_590), .Y(n_648) );
OAI21xp33_ASAP7_75t_SL g673 ( .A1(n_541), .A2(n_551), .B(n_578), .Y(n_673) );
OAI22xp33_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_546), .B1(n_551), .B2(n_554), .Y(n_542) );
INVxp33_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_544), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_545), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g599 ( .A(n_545), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g699 ( .A(n_545), .B(n_640), .Y(n_699) );
OR2x2_ASAP7_75t_L g723 ( .A(n_545), .B(n_617), .Y(n_723) );
AOI21xp33_ASAP7_75t_L g706 ( .A1(n_546), .A2(n_605), .B(n_707), .Y(n_706) );
OR2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_550), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
INVx1_ASAP7_75t_L g583 ( .A(n_548), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_548), .B(n_553), .Y(n_601) );
AND2x2_ASAP7_75t_L g623 ( .A(n_549), .B(n_596), .Y(n_623) );
INVx1_ASAP7_75t_L g636 ( .A(n_549), .Y(n_636) );
OR2x2_ASAP7_75t_L g641 ( .A(n_549), .B(n_575), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_552), .B(n_590), .Y(n_589) );
OAI22xp33_ASAP7_75t_L g571 ( .A1(n_553), .A2(n_572), .B1(n_577), .B2(n_581), .Y(n_571) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_556), .A2(n_614), .B1(n_621), .B2(n_622), .Y(n_620) );
AND2x2_ASAP7_75t_L g698 ( .A(n_556), .B(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_558), .B(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g717 ( .A(n_558), .B(n_600), .Y(n_717) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OA21x2_ASAP7_75t_L g575 ( .A1(n_560), .A2(n_568), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AOI221xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_583), .B1(n_584), .B2(n_589), .C(n_591), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_573), .B(n_575), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_573), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g592 ( .A(n_574), .Y(n_592) );
O2A1O1Ixp33_ASAP7_75t_L g679 ( .A1(n_574), .A2(n_680), .B(n_681), .C(n_682), .Y(n_679) );
AND2x2_ASAP7_75t_L g684 ( .A(n_574), .B(n_664), .Y(n_684) );
O2A1O1Ixp33_ASAP7_75t_SL g722 ( .A1(n_574), .A2(n_663), .B(n_723), .C(n_724), .Y(n_722) );
BUFx3_ASAP7_75t_L g614 ( .A(n_575), .Y(n_614) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_578), .B(n_635), .Y(n_678) );
AOI211xp5_ASAP7_75t_L g697 ( .A1(n_578), .A2(n_698), .B(n_700), .C(n_706), .Y(n_697) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
INVxp67_ASAP7_75t_L g658 ( .A(n_580), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_582), .B(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_585), .B(n_587), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
AOI211xp5_ASAP7_75t_L g602 ( .A1(n_586), .A2(n_603), .B(n_604), .C(n_612), .Y(n_602) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g687 ( .A(n_590), .Y(n_687) );
OR2x2_ASAP7_75t_L g704 ( .A(n_590), .B(n_634), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_593), .B1(n_598), .B2(n_601), .Y(n_591) );
OAI22xp33_ASAP7_75t_L g604 ( .A1(n_593), .A2(n_605), .B1(n_606), .B2(n_607), .Y(n_604) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
OR2x2_ASAP7_75t_L g691 ( .A(n_595), .B(n_635), .Y(n_691) );
INVx1_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g646 ( .A(n_596), .B(n_636), .Y(n_646) );
INVx1_ASAP7_75t_L g654 ( .A(n_597), .Y(n_654) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_600), .B(n_614), .Y(n_662) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_610), .B(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g719 ( .A(n_611), .Y(n_719) );
AOI21xp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_615), .B(n_618), .Y(n_612) );
INVx1_ASAP7_75t_L g649 ( .A(n_613), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_614), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_614), .B(n_645), .Y(n_644) );
NAND2x1p5_ASAP7_75t_L g665 ( .A(n_614), .B(n_640), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_614), .B(n_661), .Y(n_672) );
OAI211xp5_ASAP7_75t_L g676 ( .A1(n_614), .A2(n_624), .B(n_664), .C(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
AOI221xp5_ASAP7_75t_SL g619 ( .A1(n_620), .A2(n_624), .B1(n_626), .B2(n_630), .C(n_631), .Y(n_619) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVxp67_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_628), .B(n_636), .Y(n_710) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
O2A1O1Ixp33_ASAP7_75t_L g721 ( .A1(n_630), .A2(n_645), .B(n_647), .C(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_633), .B(n_640), .Y(n_705) );
NAND2xp5_ASAP7_75t_SL g724 ( .A(n_634), .B(n_687), .Y(n_724) );
CKINVDCx16_ASAP7_75t_R g634 ( .A(n_635), .Y(n_634) );
INVxp33_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .Y(n_638) );
AOI21xp33_ASAP7_75t_SL g650 ( .A1(n_639), .A2(n_651), .B(n_653), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_639), .B(n_712), .Y(n_711) );
INVx2_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_640), .B(n_694), .Y(n_693) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_646), .B1(n_647), .B2(n_649), .C(n_650), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_646), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g680 ( .A(n_652), .Y(n_680) );
NAND5xp2_ASAP7_75t_L g655 ( .A(n_656), .B(n_683), .C(n_697), .D(n_708), .E(n_721), .Y(n_655) );
AOI211xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_659), .B(n_666), .C(n_679), .Y(n_656) );
INVx2_ASAP7_75t_SL g703 ( .A(n_657), .Y(n_703) );
NAND4xp25_ASAP7_75t_SL g659 ( .A(n_660), .B(n_662), .C(n_663), .D(n_665), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx3_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OAI211xp5_ASAP7_75t_SL g666 ( .A1(n_665), .A2(n_667), .B(n_670), .C(n_676), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g667 ( .A(n_668), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_668), .A2(n_709), .B1(n_711), .B2(n_713), .C(n_715), .Y(n_708) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AOI221xp5_ASAP7_75t_SL g683 ( .A1(n_684), .A2(n_685), .B1(n_688), .B2(n_690), .C(n_692), .Y(n_683) );
AND2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_691), .A2(n_714), .B1(n_716), .B2(n_718), .Y(n_715) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_703), .B1(n_704), .B2(n_705), .Y(n_700) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx3_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
endmodule