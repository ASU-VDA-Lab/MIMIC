module fake_netlist_6_2009_n_178 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_17, n_23, n_12, n_20, n_7, n_2, n_5, n_19, n_25, n_178);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;
input n_25;

output n_178;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_28;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_47;
wire n_62;
wire n_29;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_108;
wire n_94;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_35;
wire n_115;
wire n_69;
wire n_128;
wire n_30;
wire n_79;
wire n_43;
wire n_171;
wire n_31;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_22),
.Y(n_31)
);

INVxp33_ASAP7_75t_SL g32 ( 
.A(n_24),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

INVxp33_ASAP7_75t_SL g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVxp33_ASAP7_75t_SL g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

INVxp33_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_0),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_29),
.B(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_48),
.B(n_3),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_32),
.B(n_3),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_34),
.B(n_4),
.Y(n_70)
);

OR2x6_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_43),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

AND2x6_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_66),
.Y(n_75)
);

AO22x2_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_76)
);

NAND2x1p5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_42),
.Y(n_77)
);

NAND2x1p5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_52),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_49),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_39),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

AO22x2_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_31),
.B1(n_38),
.B2(n_33),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_R g86 ( 
.A(n_79),
.B(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_74),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_59),
.Y(n_89)
);

OR2x6_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_52),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_80),
.Y(n_96)
);

OR2x6_ASAP7_75t_SL g97 ( 
.A(n_76),
.B(n_58),
.Y(n_97)
);

NAND2x1p5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_80),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_72),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_81),
.B(n_60),
.C(n_57),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_53),
.B(n_71),
.C(n_77),
.Y(n_103)
);

BUFx2_ASAP7_75t_R g104 ( 
.A(n_97),
.Y(n_104)
);

OAI21x1_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_77),
.B(n_84),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_96),
.B1(n_89),
.B2(n_93),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_96),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_90),
.B(n_71),
.C(n_91),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_90),
.Y(n_109)
);

AND2x4_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_90),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_88),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_74),
.B(n_90),
.Y(n_112)
);

OAI21x1_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_98),
.B(n_99),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_110),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_103),
.B(n_93),
.C(n_101),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_71),
.B1(n_109),
.B2(n_76),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_111),
.Y(n_123)
);

OA21x2_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_106),
.B(n_107),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

AOI31xp33_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_100),
.A3(n_112),
.B(n_97),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_115),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_71),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_125),
.A2(n_83),
.B1(n_74),
.B2(n_47),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_83),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

NAND3xp33_ASAP7_75t_SL g136 ( 
.A(n_122),
.B(n_64),
.C(n_62),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_135),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_104),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_123),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_126),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_127),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_126),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_118),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_142),
.B(n_127),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g146 ( 
.A1(n_142),
.A2(n_83),
.B(n_104),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_R g150 ( 
.A(n_138),
.B(n_144),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_124),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_124),
.B(n_119),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_130),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_124),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_130),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

NOR2x1_ASAP7_75t_SL g157 ( 
.A(n_145),
.B(n_153),
.Y(n_157)
);

NAND2xp33_ASAP7_75t_SL g158 ( 
.A(n_150),
.B(n_146),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_68),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_54),
.B(n_68),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_129),
.Y(n_162)
);

OAI221xp5_ASAP7_75t_SL g163 ( 
.A1(n_158),
.A2(n_69),
.B1(n_9),
.B2(n_10),
.C(n_128),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_121),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_14),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_160),
.A2(n_121),
.B(n_128),
.Y(n_167)
);

AOI221xp5_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_154),
.B1(n_155),
.B2(n_63),
.C(n_82),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

AND3x4_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_121),
.C(n_99),
.Y(n_170)
);

OA21x2_ASAP7_75t_L g171 ( 
.A1(n_162),
.A2(n_164),
.B(n_167),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_170),
.A2(n_128),
.B1(n_63),
.B2(n_98),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_168),
.A2(n_63),
.B1(n_91),
.B2(n_86),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_171),
.A2(n_63),
.B1(n_94),
.B2(n_95),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_172),
.A2(n_169),
.B1(n_25),
.B2(n_26),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_174),
.A2(n_94),
.B1(n_95),
.B2(n_173),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_176),
.B1(n_94),
.B2(n_95),
.Y(n_178)
);


endmodule