module fake_jpeg_16680_n_207 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_207);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_207;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_40),
.Y(n_49)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_0),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_28),
.B1(n_29),
.B2(n_22),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_44),
.B1(n_31),
.B2(n_19),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_28),
.B1(n_29),
.B2(n_22),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_45),
.B(n_57),
.Y(n_77)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_19),
.B(n_2),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_59),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_35),
.A2(n_19),
.B1(n_15),
.B2(n_21),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_21),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_21),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_61),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_25),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_25),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_63),
.B(n_67),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_51),
.A2(n_48),
.B1(n_59),
.B2(n_57),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_66),
.B1(n_82),
.B2(n_61),
.Y(n_83)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_70),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_36),
.B1(n_31),
.B2(n_27),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_27),
.Y(n_67)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_26),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_16),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_72),
.B(n_54),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_24),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_58),
.B(n_54),
.Y(n_89)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_45),
.A2(n_36),
.B1(n_33),
.B2(n_18),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_83),
.A2(n_68),
.B1(n_73),
.B2(n_18),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_77),
.B(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_84),
.B(n_92),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_49),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_104),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

AO21x1_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_93),
.B(n_26),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_74),
.A2(n_60),
.B(n_33),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_96),
.B(n_76),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_50),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_79),
.Y(n_109)
);

NOR2x1_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_50),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_74),
.A2(n_78),
.B1(n_47),
.B2(n_82),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_100),
.B1(n_103),
.B2(n_30),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_75),
.A2(n_47),
.B(n_53),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_71),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_70),
.A2(n_62),
.B1(n_33),
.B2(n_18),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_102),
.B1(n_73),
.B2(n_69),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_75),
.A2(n_62),
.B1(n_33),
.B2(n_4),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_77),
.A2(n_30),
.B1(n_24),
.B2(n_26),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_68),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_76),
.B(n_26),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_105),
.A2(n_104),
.B(n_91),
.Y(n_129)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_1),
.Y(n_106)
);

A2O1A1O1Ixp25_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_103),
.B(n_86),
.C(n_84),
.D(n_11),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_88),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_108),
.Y(n_128)
);

NAND3xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_65),
.C(n_13),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_120),
.C(n_104),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_115),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_111),
.A2(n_99),
.B1(n_87),
.B2(n_90),
.Y(n_127)
);

AO21x1_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_121),
.B(n_122),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_69),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_88),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_117),
.B(n_123),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_99),
.B1(n_87),
.B2(n_98),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_96),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_124),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_30),
.Y(n_120)
);

NOR2x1_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_26),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_102),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_100),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_126),
.B(n_134),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_141),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_133),
.Y(n_156)
);

AOI221xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_135),
.B1(n_11),
.B2(n_24),
.C(n_20),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_101),
.Y(n_139)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_101),
.Y(n_140)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_122),
.A2(n_94),
.B1(n_91),
.B2(n_83),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_106),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_142),
.B(n_113),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_118),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_109),
.C(n_112),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_149),
.C(n_141),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_120),
.C(n_123),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_SL g167 ( 
.A(n_150),
.B(n_158),
.C(n_159),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_98),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_153),
.B(n_125),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_98),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_157),
.Y(n_172)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

NOR3xp33_ASAP7_75t_SL g159 ( 
.A(n_132),
.B(n_20),
.C(n_16),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_144),
.C(n_149),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_162),
.C(n_163),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_126),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_136),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_165),
.C(n_168),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_148),
.B(n_131),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_166),
.B(n_125),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_134),
.C(n_127),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_152),
.B(n_137),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_171),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_135),
.C(n_128),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_169),
.A2(n_157),
.B1(n_155),
.B2(n_145),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_173),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_175),
.B(n_3),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_145),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_179),
.Y(n_184)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_167),
.A2(n_125),
.B(n_159),
.C(n_6),
.Y(n_180)
);

NOR3xp33_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_181),
.C(n_8),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_1),
.B(n_3),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_162),
.C(n_167),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_186),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_176),
.B(n_6),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_187),
.B(n_8),
.Y(n_193)
);

NAND4xp25_ASAP7_75t_SL g188 ( 
.A(n_182),
.B(n_20),
.C(n_16),
.D(n_18),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_18),
.Y(n_196)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_174),
.Y(n_194)
);

AOI31xp33_ASAP7_75t_SL g195 ( 
.A1(n_190),
.A2(n_8),
.A3(n_9),
.B(n_10),
.Y(n_195)
);

AOI31xp33_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_180),
.A3(n_184),
.B(n_181),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_193),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_195),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_26),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_183),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_200),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_199),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_201),
.A2(n_203),
.B(n_9),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_198),
.A2(n_195),
.B(n_189),
.Y(n_203)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_174),
.C(n_10),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_204),
.A2(n_205),
.B(n_9),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_16),
.Y(n_207)
);


endmodule