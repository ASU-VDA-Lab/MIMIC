module fake_aes_2422_n_705 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_705);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_705;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_695;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_L g80 ( .A(n_25), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_54), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_63), .Y(n_82) );
INVx1_ASAP7_75t_SL g83 ( .A(n_64), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_70), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_60), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_24), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_51), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_62), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_59), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_78), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_2), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_3), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_8), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_2), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_22), .Y(n_95) );
HB1xp67_ASAP7_75t_L g96 ( .A(n_65), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_44), .Y(n_97) );
INVxp33_ASAP7_75t_SL g98 ( .A(n_16), .Y(n_98) );
INVxp33_ASAP7_75t_L g99 ( .A(n_50), .Y(n_99) );
INVx1_ASAP7_75t_SL g100 ( .A(n_23), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_27), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_30), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_41), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_13), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_73), .Y(n_105) );
INVxp33_ASAP7_75t_SL g106 ( .A(n_20), .Y(n_106) );
INVxp67_ASAP7_75t_L g107 ( .A(n_75), .Y(n_107) );
OR2x2_ASAP7_75t_L g108 ( .A(n_58), .B(n_69), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_17), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_4), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_53), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_31), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_3), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_40), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_38), .Y(n_115) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_11), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_14), .Y(n_117) );
BUFx2_ASAP7_75t_SL g118 ( .A(n_17), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_26), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_5), .Y(n_120) );
INVxp67_ASAP7_75t_L g121 ( .A(n_68), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_61), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_6), .Y(n_123) );
BUFx3_ASAP7_75t_L g124 ( .A(n_1), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_4), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_48), .Y(n_126) );
INVxp33_ASAP7_75t_L g127 ( .A(n_8), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_82), .Y(n_128) );
AND2x4_ASAP7_75t_L g129 ( .A(n_124), .B(n_0), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_82), .Y(n_130) );
BUFx2_ASAP7_75t_L g131 ( .A(n_124), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_127), .B(n_0), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_101), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_84), .Y(n_134) );
BUFx12f_ASAP7_75t_L g135 ( .A(n_86), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_84), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_116), .B(n_1), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_85), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_85), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_96), .B(n_5), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_89), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_89), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_99), .B(n_6), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_126), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_101), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_90), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_111), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_90), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_123), .B(n_7), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_97), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_126), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_97), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_111), .Y(n_153) );
BUFx2_ASAP7_75t_L g154 ( .A(n_123), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_112), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_91), .B(n_7), .Y(n_156) );
BUFx2_ASAP7_75t_L g157 ( .A(n_86), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_115), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_112), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_114), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_115), .Y(n_161) );
BUFx2_ASAP7_75t_L g162 ( .A(n_102), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_114), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_122), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_104), .B(n_110), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_122), .Y(n_166) );
INVx5_ASAP7_75t_L g167 ( .A(n_108), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_117), .B(n_9), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_81), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_103), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_105), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_147), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_147), .Y(n_173) );
OAI221xp5_ASAP7_75t_L g174 ( .A1(n_165), .A2(n_125), .B1(n_91), .B2(n_120), .C(n_92), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_147), .Y(n_175) );
AND2x4_ASAP7_75t_SL g176 ( .A(n_137), .B(n_95), .Y(n_176) );
INVxp67_ASAP7_75t_L g177 ( .A(n_154), .Y(n_177) );
BUFx2_ASAP7_75t_L g178 ( .A(n_154), .Y(n_178) );
INVx4_ASAP7_75t_L g179 ( .A(n_167), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_147), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_147), .Y(n_181) );
INVx4_ASAP7_75t_L g182 ( .A(n_167), .Y(n_182) );
NAND2x1p5_ASAP7_75t_L g183 ( .A(n_167), .B(n_156), .Y(n_183) );
INVx2_ASAP7_75t_SL g184 ( .A(n_167), .Y(n_184) );
BUFx2_ASAP7_75t_L g185 ( .A(n_157), .Y(n_185) );
BUFx3_ASAP7_75t_L g186 ( .A(n_157), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_147), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_167), .B(n_102), .Y(n_188) );
INVx2_ASAP7_75t_SL g189 ( .A(n_167), .Y(n_189) );
BUFx3_ASAP7_75t_L g190 ( .A(n_162), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_166), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_131), .B(n_125), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_162), .B(n_92), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_133), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_166), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_133), .Y(n_196) );
INVx4_ASAP7_75t_L g197 ( .A(n_129), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_131), .B(n_93), .Y(n_198) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_133), .Y(n_199) );
AND2x6_ASAP7_75t_L g200 ( .A(n_129), .B(n_119), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_166), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_144), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_144), .Y(n_203) );
AND2x2_ASAP7_75t_SL g204 ( .A(n_129), .B(n_108), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_144), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_145), .Y(n_206) );
AND2x6_ASAP7_75t_L g207 ( .A(n_129), .B(n_93), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_143), .B(n_94), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_144), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_145), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_151), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_170), .B(n_121), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_128), .B(n_80), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_145), .Y(n_214) );
INVxp67_ASAP7_75t_L g215 ( .A(n_132), .Y(n_215) );
INVx3_ASAP7_75t_L g216 ( .A(n_156), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_151), .Y(n_217) );
AO22x2_ASAP7_75t_L g218 ( .A1(n_156), .A2(n_118), .B1(n_120), .B2(n_109), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_143), .B(n_109), .Y(n_219) );
NAND2x1p5_ASAP7_75t_L g220 ( .A(n_156), .B(n_94), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_153), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_170), .B(n_107), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_151), .Y(n_223) );
INVx1_ASAP7_75t_SL g224 ( .A(n_135), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_153), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_153), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_158), .Y(n_227) );
BUFx3_ASAP7_75t_L g228 ( .A(n_135), .Y(n_228) );
INVx3_ASAP7_75t_L g229 ( .A(n_151), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_132), .B(n_118), .Y(n_230) );
INVx1_ASAP7_75t_SL g231 ( .A(n_137), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_128), .B(n_113), .Y(n_232) );
BUFx4f_ASAP7_75t_L g233 ( .A(n_130), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_204), .A2(n_149), .B1(n_140), .B2(n_98), .Y(n_234) );
INVx2_ASAP7_75t_SL g235 ( .A(n_186), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_229), .Y(n_236) );
BUFx2_ASAP7_75t_L g237 ( .A(n_178), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_229), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_229), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_186), .B(n_171), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_220), .Y(n_241) );
INVxp67_ASAP7_75t_SL g242 ( .A(n_220), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_220), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_178), .B(n_171), .Y(n_244) );
HAxp5_ASAP7_75t_L g245 ( .A(n_231), .B(n_168), .CON(n_245), .SN(n_245) );
BUFx3_ASAP7_75t_L g246 ( .A(n_190), .Y(n_246) );
INVx2_ASAP7_75t_SL g247 ( .A(n_190), .Y(n_247) );
OR2x2_ASAP7_75t_L g248 ( .A(n_185), .B(n_150), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_204), .A2(n_142), .B1(n_164), .B2(n_163), .Y(n_249) );
INVxp67_ASAP7_75t_L g250 ( .A(n_185), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_215), .B(n_142), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_204), .B(n_146), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_191), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_191), .Y(n_254) );
AND2x4_ASAP7_75t_L g255 ( .A(n_192), .B(n_146), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_177), .B(n_141), .Y(n_256) );
OR2x6_ASAP7_75t_L g257 ( .A(n_228), .B(n_150), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_195), .Y(n_258) );
INVx1_ASAP7_75t_SL g259 ( .A(n_207), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_213), .B(n_141), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_195), .Y(n_261) );
AOI211xp5_ASAP7_75t_L g262 ( .A1(n_174), .A2(n_139), .B(n_164), .C(n_163), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_233), .B(n_106), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_201), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_208), .B(n_139), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_233), .B(n_138), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_201), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_228), .Y(n_268) );
INVxp67_ASAP7_75t_L g269 ( .A(n_232), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_233), .B(n_138), .Y(n_270) );
INVx5_ASAP7_75t_L g271 ( .A(n_207), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_207), .B(n_148), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_202), .Y(n_273) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_207), .Y(n_274) );
INVx3_ASAP7_75t_L g275 ( .A(n_197), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_202), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_203), .Y(n_277) );
INVx2_ASAP7_75t_SL g278 ( .A(n_192), .Y(n_278) );
OR2x2_ASAP7_75t_L g279 ( .A(n_224), .B(n_155), .Y(n_279) );
INVx2_ASAP7_75t_SL g280 ( .A(n_192), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_203), .Y(n_281) );
INVx3_ASAP7_75t_L g282 ( .A(n_197), .Y(n_282) );
INVx5_ASAP7_75t_L g283 ( .A(n_207), .Y(n_283) );
INVx5_ASAP7_75t_L g284 ( .A(n_207), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_205), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_207), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_192), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_208), .B(n_148), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_205), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_194), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_209), .Y(n_291) );
BUFx3_ASAP7_75t_L g292 ( .A(n_196), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_209), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_219), .B(n_136), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_211), .Y(n_295) );
INVx5_ASAP7_75t_L g296 ( .A(n_179), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_218), .A2(n_216), .B(n_211), .Y(n_297) );
AOI22x1_ASAP7_75t_L g298 ( .A1(n_218), .A2(n_169), .B1(n_158), .B2(n_160), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_194), .Y(n_299) );
CKINVDCx20_ASAP7_75t_R g300 ( .A(n_176), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_273), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_269), .B(n_176), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g303 ( .A(n_269), .B(n_230), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_274), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_276), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_277), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_255), .B(n_232), .Y(n_307) );
OAI22xp5_ASAP7_75t_SL g308 ( .A1(n_300), .A2(n_197), .B1(n_183), .B2(n_222), .Y(n_308) );
CKINVDCx6p67_ASAP7_75t_R g309 ( .A(n_257), .Y(n_309) );
INVxp67_ASAP7_75t_L g310 ( .A(n_237), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_242), .B(n_230), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_281), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_242), .A2(n_218), .B1(n_216), .B2(n_183), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_285), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_289), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_291), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_257), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_257), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_287), .A2(n_218), .B1(n_200), .B2(n_219), .Y(n_319) );
NOR2x1p5_ASAP7_75t_L g320 ( .A(n_268), .B(n_193), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g321 ( .A1(n_249), .A2(n_216), .B1(n_183), .B2(n_212), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_250), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_241), .B(n_193), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_274), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_293), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_287), .A2(n_200), .B1(n_198), .B2(n_223), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_255), .B(n_198), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_274), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_286), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_295), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_243), .A2(n_217), .B1(n_223), .B2(n_182), .Y(n_331) );
INVx3_ASAP7_75t_L g332 ( .A(n_286), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_278), .A2(n_200), .B1(n_217), .B2(n_188), .Y(n_333) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_250), .Y(n_334) );
NOR2x1_ASAP7_75t_R g335 ( .A(n_246), .B(n_179), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_292), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_253), .Y(n_337) );
AO22x1_ASAP7_75t_L g338 ( .A1(n_286), .A2(n_200), .B1(n_130), .B2(n_160), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_254), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_271), .B(n_200), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_258), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_235), .Y(n_342) );
CKINVDCx11_ASAP7_75t_R g343 ( .A(n_240), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_261), .Y(n_344) );
INVx4_ASAP7_75t_L g345 ( .A(n_271), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_271), .B(n_200), .Y(n_346) );
INVx4_ASAP7_75t_L g347 ( .A(n_271), .Y(n_347) );
AND2x4_ASAP7_75t_L g348 ( .A(n_283), .B(n_200), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_240), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_264), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_267), .Y(n_351) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_283), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_252), .A2(n_179), .B1(n_182), .B2(n_189), .Y(n_353) );
INVxp67_ASAP7_75t_L g354 ( .A(n_322), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_311), .A2(n_280), .B1(n_234), .B2(n_244), .Y(n_355) );
OAI22xp33_ASAP7_75t_L g356 ( .A1(n_309), .A2(n_279), .B1(n_248), .B2(n_252), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_319), .A2(n_294), .B1(n_297), .B2(n_288), .Y(n_357) );
OAI21xp5_ASAP7_75t_L g358 ( .A1(n_301), .A2(n_297), .B(n_298), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_311), .A2(n_294), .B1(n_265), .B2(n_259), .Y(n_359) );
AOI21xp33_ASAP7_75t_L g360 ( .A1(n_302), .A2(n_247), .B(n_256), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_311), .B(n_245), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_311), .B(n_251), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_301), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_313), .A2(n_262), .B1(n_259), .B2(n_152), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_323), .A2(n_251), .B1(n_282), .B2(n_275), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_306), .Y(n_366) );
NAND2xp5_ASAP7_75t_SL g367 ( .A(n_317), .B(n_283), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_306), .Y(n_368) );
O2A1O1Ixp33_ASAP7_75t_L g369 ( .A1(n_321), .A2(n_263), .B(n_266), .C(n_270), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_323), .B(n_260), .Y(n_370) );
INVx3_ASAP7_75t_L g371 ( .A(n_352), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_305), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_323), .A2(n_275), .B1(n_282), .B2(n_272), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_312), .Y(n_374) );
OAI221xp5_ASAP7_75t_L g375 ( .A1(n_303), .A2(n_260), .B1(n_272), .B2(n_236), .C(n_238), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_323), .A2(n_239), .B1(n_283), .B2(n_284), .Y(n_376) );
INVx6_ASAP7_75t_L g377 ( .A(n_345), .Y(n_377) );
O2A1O1Ixp33_ASAP7_75t_SL g378 ( .A1(n_305), .A2(n_184), .B(n_189), .C(n_134), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_327), .B(n_239), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_330), .Y(n_380) );
INVxp33_ASAP7_75t_SL g381 ( .A(n_317), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_327), .B(n_284), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_312), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_340), .B(n_284), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_308), .A2(n_159), .B1(n_155), .B2(n_152), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_334), .A2(n_284), .B1(n_296), .B2(n_159), .Y(n_386) );
A2O1A1Ixp33_ASAP7_75t_L g387 ( .A1(n_385), .A2(n_330), .B(n_339), .C(n_341), .Y(n_387) );
CKINVDCx11_ASAP7_75t_R g388 ( .A(n_366), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_356), .A2(n_307), .B1(n_310), .B2(n_349), .C(n_350), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_366), .Y(n_390) );
AOI21xp33_ASAP7_75t_L g391 ( .A1(n_357), .A2(n_335), .B(n_342), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_366), .Y(n_392) );
OAI22xp33_ASAP7_75t_L g393 ( .A1(n_385), .A2(n_309), .B1(n_318), .B2(n_349), .Y(n_393) );
OAI221xp5_ASAP7_75t_L g394 ( .A1(n_355), .A2(n_326), .B1(n_318), .B2(n_342), .C(n_341), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_368), .B(n_337), .Y(n_395) );
BUFx2_ASAP7_75t_L g396 ( .A(n_368), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_368), .B(n_339), .Y(n_397) );
OAI22xp33_ASAP7_75t_L g398 ( .A1(n_362), .A2(n_350), .B1(n_344), .B2(n_351), .Y(n_398) );
INVx3_ASAP7_75t_L g399 ( .A(n_384), .Y(n_399) );
CKINVDCx6p67_ASAP7_75t_R g400 ( .A(n_384), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g401 ( .A1(n_358), .A2(n_338), .B(n_314), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_374), .Y(n_402) );
BUFx2_ASAP7_75t_L g403 ( .A(n_374), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_361), .A2(n_320), .B1(n_343), .B2(n_351), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_361), .A2(n_320), .B1(n_344), .B2(n_337), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_374), .Y(n_406) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_383), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_383), .Y(n_408) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_383), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_363), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_363), .B(n_314), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_372), .B(n_315), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_354), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_372), .Y(n_414) );
BUFx2_ASAP7_75t_L g415 ( .A(n_380), .Y(n_415) );
AOI22xp33_ASAP7_75t_SL g416 ( .A1(n_394), .A2(n_381), .B1(n_364), .B2(n_380), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_392), .Y(n_417) );
OAI31xp33_ASAP7_75t_L g418 ( .A1(n_393), .A2(n_364), .A3(n_359), .B(n_360), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_389), .A2(n_370), .B1(n_375), .B2(n_382), .Y(n_419) );
AOI22xp33_ASAP7_75t_SL g420 ( .A1(n_415), .A2(n_377), .B1(n_358), .B2(n_382), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_404), .A2(n_379), .B1(n_134), .B2(n_136), .C(n_365), .Y(n_421) );
INVx1_ASAP7_75t_SL g422 ( .A(n_388), .Y(n_422) );
OAI31xp33_ASAP7_75t_L g423 ( .A1(n_398), .A2(n_369), .A3(n_378), .B(n_315), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g424 ( .A1(n_405), .A2(n_169), .B1(n_161), .B2(n_158), .C(n_386), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_397), .B(n_411), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_413), .A2(n_169), .B1(n_161), .B2(n_373), .C(n_325), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_410), .Y(n_427) );
OAI211xp5_ASAP7_75t_SL g428 ( .A1(n_391), .A2(n_83), .B(n_100), .C(n_87), .Y(n_428) );
AOI221xp5_ASAP7_75t_L g429 ( .A1(n_387), .A2(n_325), .B1(n_316), .B2(n_194), .C(n_199), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_415), .A2(n_316), .B1(n_377), .B2(n_336), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_411), .A2(n_331), .B1(n_336), .B2(n_377), .Y(n_431) );
OAI33xp33_ASAP7_75t_L g432 ( .A1(n_414), .A2(n_173), .A3(n_180), .B1(n_181), .B2(n_175), .B3(n_225), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_410), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g434 ( .A1(n_414), .A2(n_210), .B1(n_194), .B2(n_226), .C(n_199), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_399), .A2(n_377), .B1(n_367), .B2(n_384), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_392), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_392), .Y(n_437) );
AO21x2_ASAP7_75t_L g438 ( .A1(n_401), .A2(n_180), .B(n_173), .Y(n_438) );
OAI21xp5_ASAP7_75t_L g439 ( .A1(n_397), .A2(n_353), .B(n_206), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g440 ( .A1(n_412), .A2(n_210), .B1(n_226), .B2(n_199), .C(n_221), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_390), .Y(n_441) );
INVx3_ASAP7_75t_L g442 ( .A(n_395), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_390), .B(n_371), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_406), .Y(n_444) );
INVx3_ASAP7_75t_SL g445 ( .A(n_400), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_395), .Y(n_446) );
AOI221xp5_ASAP7_75t_L g447 ( .A1(n_406), .A2(n_210), .B1(n_226), .B2(n_199), .C(n_221), .Y(n_447) );
OAI21x1_ASAP7_75t_L g448 ( .A1(n_408), .A2(n_371), .B(n_328), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_408), .B(n_196), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_408), .B(n_371), .Y(n_450) );
INVx5_ASAP7_75t_L g451 ( .A(n_442), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_427), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_423), .B(n_407), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_427), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_425), .B(n_396), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_433), .Y(n_456) );
NOR3xp33_ASAP7_75t_SL g457 ( .A(n_428), .B(n_88), .C(n_400), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_425), .B(n_396), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_442), .B(n_402), .Y(n_459) );
OAI221xp5_ASAP7_75t_L g460 ( .A1(n_416), .A2(n_399), .B1(n_403), .B2(n_402), .C(n_376), .Y(n_460) );
NAND3xp33_ASAP7_75t_L g461 ( .A(n_418), .B(n_221), .C(n_199), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_433), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_442), .B(n_403), .Y(n_463) );
INVxp67_ASAP7_75t_L g464 ( .A(n_446), .Y(n_464) );
AO21x2_ASAP7_75t_L g465 ( .A1(n_438), .A2(n_181), .B(n_175), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_419), .A2(n_399), .B1(n_407), .B2(n_409), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_441), .B(n_399), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_441), .B(n_407), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_444), .Y(n_469) );
AOI33xp33_ASAP7_75t_L g470 ( .A1(n_422), .A2(n_227), .A3(n_225), .B1(n_214), .B2(n_206), .B3(n_13), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_417), .Y(n_471) );
INVx3_ASAP7_75t_L g472 ( .A(n_417), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_444), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_436), .B(n_407), .Y(n_474) );
NAND3xp33_ASAP7_75t_L g475 ( .A(n_418), .B(n_194), .C(n_210), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_436), .Y(n_476) );
AOI221xp5_ASAP7_75t_L g477 ( .A1(n_421), .A2(n_221), .B1(n_210), .B2(n_226), .C(n_214), .Y(n_477) );
NAND3xp33_ASAP7_75t_SL g478 ( .A(n_422), .B(n_227), .C(n_10), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_443), .Y(n_479) );
AND2x2_ASAP7_75t_SL g480 ( .A(n_445), .B(n_407), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_445), .A2(n_409), .B1(n_407), .B2(n_371), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_443), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_437), .B(n_409), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_437), .Y(n_484) );
OAI31xp33_ASAP7_75t_L g485 ( .A1(n_423), .A2(n_340), .A3(n_346), .B(n_348), .Y(n_485) );
AOI221xp5_ASAP7_75t_L g486 ( .A1(n_426), .A2(n_221), .B1(n_226), .B2(n_409), .C(n_338), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_450), .B(n_409), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_450), .Y(n_488) );
OAI33xp33_ASAP7_75t_L g489 ( .A1(n_449), .A2(n_9), .A3(n_10), .B1(n_11), .B2(n_12), .B3(n_14), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_431), .Y(n_490) );
NAND3xp33_ASAP7_75t_L g491 ( .A(n_424), .B(n_172), .C(n_409), .Y(n_491) );
NOR3xp33_ASAP7_75t_L g492 ( .A(n_432), .B(n_335), .C(n_187), .Y(n_492) );
INVx4_ASAP7_75t_L g493 ( .A(n_445), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_430), .B(n_12), .Y(n_494) );
BUFx2_ASAP7_75t_L g495 ( .A(n_448), .Y(n_495) );
INVx2_ASAP7_75t_SL g496 ( .A(n_448), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_420), .B(n_15), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_438), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_438), .B(n_15), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_431), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_487), .B(n_439), .Y(n_501) );
AOI31xp33_ASAP7_75t_L g502 ( .A1(n_478), .A2(n_429), .A3(n_435), .B(n_439), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_469), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_464), .B(n_16), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_469), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_473), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_487), .B(n_18), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_473), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_455), .B(n_18), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_455), .B(n_434), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_452), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_454), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_456), .Y(n_513) );
OAI33xp33_ASAP7_75t_L g514 ( .A1(n_462), .A2(n_187), .A3(n_299), .B1(n_290), .B2(n_29), .B3(n_32), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_479), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_472), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_459), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_482), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_468), .B(n_440), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_458), .B(n_447), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_472), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_472), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_488), .B(n_19), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_500), .B(n_172), .Y(n_524) );
AOI21x1_ASAP7_75t_L g525 ( .A1(n_499), .A2(n_384), .B(n_348), .Y(n_525) );
NAND3xp33_ASAP7_75t_L g526 ( .A(n_457), .B(n_172), .C(n_333), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_490), .B(n_172), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_459), .B(n_21), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_500), .B(n_28), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_467), .Y(n_530) );
NOR3xp33_ASAP7_75t_L g531 ( .A(n_489), .B(n_347), .C(n_345), .Y(n_531) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_463), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_483), .B(n_33), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_471), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_463), .B(n_34), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_491), .A2(n_329), .B(n_324), .Y(n_536) );
NOR2x1p5_ASAP7_75t_L g537 ( .A(n_493), .B(n_345), .Y(n_537) );
AOI21xp33_ASAP7_75t_L g538 ( .A1(n_494), .A2(n_332), .B(n_328), .Y(n_538) );
AOI221xp5_ASAP7_75t_L g539 ( .A1(n_497), .A2(n_182), .B1(n_184), .B2(n_340), .C(n_346), .Y(n_539) );
NOR2x1_ASAP7_75t_L g540 ( .A(n_493), .B(n_347), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g541 ( .A(n_493), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_471), .B(n_476), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_476), .Y(n_543) );
OAI21xp5_ASAP7_75t_L g544 ( .A1(n_470), .A2(n_348), .B(n_340), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_484), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_474), .B(n_35), .Y(n_546) );
NOR3xp33_ASAP7_75t_L g547 ( .A(n_470), .B(n_347), .C(n_332), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_499), .Y(n_548) );
NOR2x1_ASAP7_75t_L g549 ( .A(n_497), .B(n_348), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_461), .A2(n_329), .B(n_324), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_474), .B(n_36), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_451), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_483), .B(n_37), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_451), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_498), .B(n_39), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_494), .B(n_42), .Y(n_556) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_451), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_451), .B(n_43), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_548), .B(n_451), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_515), .B(n_480), .Y(n_560) );
OAI22xp33_ASAP7_75t_L g561 ( .A1(n_541), .A2(n_460), .B1(n_466), .B2(n_475), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_511), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_501), .B(n_498), .Y(n_563) );
INVx1_ASAP7_75t_SL g564 ( .A(n_541), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_517), .B(n_495), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_532), .B(n_480), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_512), .Y(n_567) );
INVxp67_ASAP7_75t_SL g568 ( .A(n_557), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_513), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_542), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_516), .B(n_496), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_516), .B(n_521), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_518), .B(n_453), .Y(n_573) );
AND2x4_ASAP7_75t_SL g574 ( .A(n_507), .B(n_481), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_504), .B(n_453), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_507), .B(n_496), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_549), .B(n_465), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_502), .B(n_465), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_503), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_505), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_530), .B(n_465), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_506), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_509), .B(n_485), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_508), .Y(n_584) );
AND4x1_ASAP7_75t_L g585 ( .A(n_540), .B(n_486), .C(n_477), .D(n_492), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_545), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_509), .B(n_45), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_542), .B(n_46), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_519), .B(n_47), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_527), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_519), .B(n_49), .Y(n_591) );
INVx3_ASAP7_75t_L g592 ( .A(n_552), .Y(n_592) );
XNOR2xp5_ASAP7_75t_L g593 ( .A(n_537), .B(n_346), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_527), .Y(n_594) );
NAND2x1p5_ASAP7_75t_L g595 ( .A(n_546), .B(n_324), .Y(n_595) );
INVx1_ASAP7_75t_SL g596 ( .A(n_533), .Y(n_596) );
NAND2xp33_ASAP7_75t_L g597 ( .A(n_523), .B(n_329), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_521), .B(n_52), .Y(n_598) );
INVx4_ASAP7_75t_L g599 ( .A(n_554), .Y(n_599) );
INVx3_ASAP7_75t_L g600 ( .A(n_534), .Y(n_600) );
BUFx2_ASAP7_75t_L g601 ( .A(n_533), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_534), .Y(n_602) );
OAI21xp33_ASAP7_75t_L g603 ( .A1(n_556), .A2(n_332), .B(n_328), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_543), .B(n_55), .Y(n_604) );
AOI31xp33_ASAP7_75t_L g605 ( .A1(n_556), .A2(n_346), .A3(n_57), .B(n_66), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_543), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_522), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_510), .B(n_56), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_522), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_524), .Y(n_610) );
OR2x2_ASAP7_75t_L g611 ( .A(n_563), .B(n_546), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_563), .B(n_551), .Y(n_612) );
AOI221x1_ASAP7_75t_L g613 ( .A1(n_578), .A2(n_558), .B1(n_531), .B2(n_538), .C(n_547), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_562), .Y(n_614) );
AOI21xp33_ASAP7_75t_L g615 ( .A1(n_578), .A2(n_575), .B(n_561), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_564), .Y(n_616) );
AND2x4_ASAP7_75t_L g617 ( .A(n_592), .B(n_525), .Y(n_617) );
AND2x4_ASAP7_75t_SL g618 ( .A(n_599), .B(n_566), .Y(n_618) );
BUFx3_ASAP7_75t_L g619 ( .A(n_592), .Y(n_619) );
INVxp67_ASAP7_75t_SL g620 ( .A(n_568), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_600), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_576), .B(n_555), .Y(n_622) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_592), .Y(n_623) );
INVxp67_ASAP7_75t_SL g624 ( .A(n_600), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_600), .Y(n_625) );
CKINVDCx14_ASAP7_75t_R g626 ( .A(n_601), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_567), .Y(n_627) );
XOR2x2_ASAP7_75t_L g628 ( .A(n_593), .B(n_539), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_570), .B(n_551), .Y(n_629) );
NOR3xp33_ASAP7_75t_SL g630 ( .A(n_561), .B(n_526), .C(n_514), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_569), .B(n_520), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_575), .B(n_535), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_572), .B(n_553), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_572), .B(n_553), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_586), .Y(n_635) );
NAND4xp25_ASAP7_75t_L g636 ( .A(n_583), .B(n_544), .C(n_528), .D(n_529), .Y(n_636) );
XOR2x2_ASAP7_75t_L g637 ( .A(n_596), .B(n_529), .Y(n_637) );
OAI22x1_ASAP7_75t_L g638 ( .A1(n_599), .A2(n_524), .B1(n_536), .B2(n_550), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_590), .B(n_67), .Y(n_639) );
OAI221xp5_ASAP7_75t_SL g640 ( .A1(n_587), .A2(n_304), .B1(n_72), .B2(n_74), .C(n_76), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_594), .B(n_71), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_599), .B(n_324), .Y(n_642) );
AOI21xp33_ASAP7_75t_L g643 ( .A1(n_577), .A2(n_77), .B(n_79), .Y(n_643) );
OAI221xp5_ASAP7_75t_SL g644 ( .A1(n_589), .A2(n_304), .B1(n_352), .B2(n_324), .C(n_329), .Y(n_644) );
NAND2xp33_ASAP7_75t_R g645 ( .A(n_577), .B(n_565), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_579), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_580), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_574), .A2(n_304), .B1(n_329), .B2(n_352), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_582), .Y(n_649) );
AOI211xp5_ASAP7_75t_SL g650 ( .A1(n_605), .A2(n_296), .B(n_352), .C(n_597), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_584), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_560), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_606), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_607), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_573), .B(n_296), .Y(n_655) );
INVxp67_ASAP7_75t_L g656 ( .A(n_581), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_602), .Y(n_657) );
NOR2x1_ASAP7_75t_L g658 ( .A(n_597), .B(n_352), .Y(n_658) );
OAI21xp33_ASAP7_75t_SL g659 ( .A1(n_559), .A2(n_296), .B(n_588), .Y(n_659) );
XNOR2x1_ASAP7_75t_L g660 ( .A(n_595), .B(n_591), .Y(n_660) );
NAND2xp33_ASAP7_75t_SL g661 ( .A(n_610), .B(n_598), .Y(n_661) );
AOI211xp5_ASAP7_75t_L g662 ( .A1(n_603), .A2(n_608), .B(n_571), .C(n_610), .Y(n_662) );
NOR3xp33_ASAP7_75t_L g663 ( .A(n_598), .B(n_604), .C(n_571), .Y(n_663) );
AOI211xp5_ASAP7_75t_SL g664 ( .A1(n_574), .A2(n_609), .B(n_602), .C(n_585), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_609), .Y(n_665) );
INVx2_ASAP7_75t_SL g666 ( .A(n_595), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_564), .B(n_422), .Y(n_667) );
AOI21xp5_ASAP7_75t_L g668 ( .A1(n_605), .A2(n_597), .B(n_561), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_562), .Y(n_669) );
INVxp33_ASAP7_75t_SL g670 ( .A(n_667), .Y(n_670) );
AO22x2_ASAP7_75t_L g671 ( .A1(n_616), .A2(n_620), .B1(n_668), .B2(n_617), .Y(n_671) );
BUFx2_ASAP7_75t_L g672 ( .A(n_626), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g673 ( .A1(n_615), .A2(n_645), .B1(n_630), .B2(n_664), .C(n_659), .Y(n_673) );
AOI221xp5_ASAP7_75t_SL g674 ( .A1(n_626), .A2(n_631), .B1(n_652), .B2(n_656), .C(n_632), .Y(n_674) );
OAI221xp5_ASAP7_75t_L g675 ( .A1(n_645), .A2(n_650), .B1(n_662), .B2(n_656), .C(n_661), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_669), .B(n_635), .Y(n_676) );
AOI21xp33_ASAP7_75t_L g677 ( .A1(n_632), .A2(n_638), .B(n_617), .Y(n_677) );
A2O1A1Ixp33_ASAP7_75t_L g678 ( .A1(n_618), .A2(n_617), .B(n_619), .C(n_623), .Y(n_678) );
AO221x1_ASAP7_75t_L g679 ( .A1(n_638), .A2(n_618), .B1(n_637), .B2(n_614), .C(n_627), .Y(n_679) );
OAI31xp33_ASAP7_75t_L g680 ( .A1(n_619), .A2(n_660), .A3(n_636), .B(n_663), .Y(n_680) );
NAND3xp33_ASAP7_75t_L g681 ( .A(n_613), .B(n_648), .C(n_655), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_621), .Y(n_682) );
NAND4xp25_ASAP7_75t_L g683 ( .A(n_648), .B(n_663), .C(n_640), .D(n_658), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_673), .A2(n_642), .B(n_637), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_676), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_672), .Y(n_686) );
A2O1A1Ixp33_ASAP7_75t_SL g687 ( .A1(n_680), .A2(n_643), .B(n_639), .C(n_641), .Y(n_687) );
AOI321xp33_ASAP7_75t_L g688 ( .A1(n_675), .A2(n_624), .A3(n_622), .B1(n_646), .B2(n_647), .C(n_649), .Y(n_688) );
INVxp67_ASAP7_75t_L g689 ( .A(n_671), .Y(n_689) );
XNOR2x1_ASAP7_75t_L g690 ( .A(n_671), .B(n_628), .Y(n_690) );
O2A1O1Ixp33_ASAP7_75t_L g691 ( .A1(n_677), .A2(n_681), .B(n_678), .C(n_670), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_686), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_690), .A2(n_674), .B1(n_679), .B2(n_683), .Y(n_693) );
AND5x1_ASAP7_75t_L g694 ( .A(n_684), .B(n_628), .C(n_644), .D(n_666), .E(n_642), .Y(n_694) );
NOR4xp25_ASAP7_75t_L g695 ( .A(n_689), .B(n_682), .C(n_651), .D(n_653), .Y(n_695) );
OAI211xp5_ASAP7_75t_SL g696 ( .A1(n_691), .A2(n_684), .B(n_687), .C(n_688), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_692), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_693), .A2(n_685), .B1(n_612), .B2(n_611), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_696), .A2(n_629), .B1(n_654), .B2(n_634), .Y(n_699) );
OAI22x1_ASAP7_75t_L g700 ( .A1(n_697), .A2(n_694), .B1(n_695), .B2(n_621), .Y(n_700) );
A2O1A1Ixp33_ASAP7_75t_SL g701 ( .A1(n_699), .A2(n_625), .B(n_657), .C(n_665), .Y(n_701) );
INVxp67_ASAP7_75t_L g702 ( .A(n_700), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_702), .Y(n_703) );
OAI22xp33_ASAP7_75t_L g704 ( .A1(n_703), .A2(n_698), .B1(n_701), .B2(n_625), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g705 ( .A1(n_704), .A2(n_633), .B(n_634), .Y(n_705) );
endmodule