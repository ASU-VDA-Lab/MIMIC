module fake_jpeg_29914_n_157 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_157);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_157;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_11),
.B(n_45),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_31),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_48),
.B(n_0),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_72),
.Y(n_79)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_74),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_69),
.A2(n_49),
.B1(n_62),
.B2(n_58),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_76),
.A2(n_85),
.B1(n_22),
.B2(n_41),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_74),
.B(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_2),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_47),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_53),
.B(n_52),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_0),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_51),
.B1(n_58),
.B2(n_62),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_51),
.B1(n_49),
.B2(n_60),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_66),
.A2(n_49),
.B1(n_53),
.B2(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_46),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_88),
.B(n_57),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_87),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_91),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_90),
.A2(n_84),
.B1(n_75),
.B2(n_7),
.Y(n_114)
);

AND2x6_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_61),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_94),
.Y(n_124)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_56),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_86),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_95),
.B(n_96),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_20),
.C(n_43),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_99),
.A2(n_3),
.B(n_6),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_100),
.A2(n_99),
.B(n_5),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_1),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_101),
.B(n_3),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_81),
.B(n_1),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_104),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_81),
.B(n_2),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_105),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_8),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_84),
.B(n_75),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_110),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_115),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_123),
.B1(n_10),
.B2(n_12),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_26),
.B(n_40),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_111),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_102),
.A2(n_6),
.B(n_8),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_119),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_9),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_127),
.C(n_19),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_90),
.A2(n_28),
.B1(n_38),
.B2(n_35),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_10),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_131),
.Y(n_142)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_138),
.B1(n_139),
.B2(n_112),
.Y(n_144)
);

AO21x1_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_137),
.B(n_140),
.Y(n_146)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_44),
.A3(n_23),
.B1(n_15),
.B2(n_16),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_120),
.A2(n_12),
.B1(n_13),
.B2(n_18),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_13),
.B1(n_33),
.B2(n_30),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_141),
.A2(n_136),
.B1(n_129),
.B2(n_134),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_144),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_133),
.A2(n_108),
.B(n_125),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_147),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_143),
.A2(n_130),
.B1(n_114),
.B2(n_145),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_118),
.C(n_138),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_150),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_148),
.B1(n_150),
.B2(n_137),
.Y(n_153)
);

AO21x1_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_146),
.B(n_142),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_154),
.A2(n_146),
.B(n_124),
.Y(n_155)
);

AOI221xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_140),
.B1(n_123),
.B2(n_109),
.C(n_112),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_32),
.Y(n_157)
);


endmodule