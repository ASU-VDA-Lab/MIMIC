module fake_jpeg_26761_n_200 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_200);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_200;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx2_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_33),
.Y(n_61)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_31),
.Y(n_40)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_43),
.Y(n_47)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_25),
.B1(n_18),
.B2(n_32),
.Y(n_48)
);

AOI22x1_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_60),
.B1(n_19),
.B2(n_38),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_49),
.B(n_53),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_25),
.B1(n_32),
.B2(n_18),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_59),
.C(n_20),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_25),
.B1(n_18),
.B2(n_32),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_54),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_26),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_26),
.Y(n_55)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_35),
.B(n_21),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_35),
.B(n_23),
.C(n_19),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_57),
.A2(n_38),
.B1(n_43),
.B2(n_30),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_28),
.B1(n_21),
.B2(n_29),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_38),
.B1(n_42),
.B2(n_34),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_50),
.A2(n_43),
.B1(n_16),
.B2(n_17),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_77),
.B1(n_44),
.B2(n_34),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_68),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_81),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_71),
.Y(n_89)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_16),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_76),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_67),
.B1(n_62),
.B2(n_42),
.Y(n_90)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_80),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_50),
.A2(n_17),
.B1(n_23),
.B2(n_19),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_79),
.Y(n_103)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_63),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_49),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_86),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_56),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_88),
.B1(n_92),
.B2(n_93),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_51),
.B1(n_59),
.B2(n_54),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_94),
.B1(n_71),
.B2(n_75),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_67),
.A2(n_73),
.B1(n_78),
.B2(n_66),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_62),
.B1(n_42),
.B2(n_34),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_66),
.A2(n_62),
.B1(n_44),
.B2(n_52),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_55),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_98),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_81),
.B(n_47),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_33),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_61),
.B(n_46),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_47),
.B(n_61),
.C(n_35),
.Y(n_100)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_33),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_61),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_84),
.B(n_20),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_105),
.B(n_110),
.Y(n_123)
);

A2O1A1O1Ixp25_ASAP7_75t_L g106 ( 
.A1(n_96),
.A2(n_35),
.B(n_33),
.C(n_36),
.D(n_39),
.Y(n_106)
);

A2O1A1O1Ixp25_ASAP7_75t_L g130 ( 
.A1(n_106),
.A2(n_100),
.B(n_99),
.C(n_98),
.D(n_89),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_39),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_109),
.A2(n_122),
.B(n_100),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_84),
.B(n_20),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_85),
.B1(n_93),
.B2(n_94),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_20),
.Y(n_113)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_119),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_68),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_115),
.B(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_61),
.Y(n_118)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_121),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_95),
.B(n_22),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_129),
.B(n_130),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_126),
.A2(n_36),
.B1(n_19),
.B2(n_22),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_117),
.Y(n_128)
);

NOR3xp33_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_110),
.C(n_105),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_118),
.A2(n_96),
.B(n_91),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_86),
.C(n_88),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_132),
.C(n_137),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_99),
.C(n_85),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_111),
.B(n_103),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_108),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_103),
.C(n_39),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_83),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_27),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_108),
.A2(n_19),
.B1(n_22),
.B2(n_68),
.Y(n_140)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_104),
.Y(n_141)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

AO221x1_ASAP7_75t_L g142 ( 
.A1(n_133),
.A2(n_114),
.B1(n_120),
.B2(n_46),
.C(n_122),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_155),
.B(n_125),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_143),
.A2(n_146),
.B1(n_148),
.B2(n_0),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_145),
.B(n_149),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_129),
.A2(n_107),
.B(n_106),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_109),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_153),
.C(n_27),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_134),
.A2(n_109),
.B1(n_107),
.B2(n_112),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_36),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_145),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_151),
.A2(n_127),
.B1(n_124),
.B2(n_134),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_27),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_154),
.A2(n_126),
.B1(n_14),
.B2(n_13),
.Y(n_160)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_157),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_136),
.C(n_132),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_159),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_130),
.C(n_123),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_160),
.A2(n_13),
.B(n_12),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_163),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_165),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_22),
.C(n_14),
.Y(n_165)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_166),
.Y(n_176)
);

OAI321xp33_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_146),
.A3(n_148),
.B1(n_152),
.B2(n_144),
.C(n_151),
.Y(n_167)
);

AOI31xp67_ASAP7_75t_L g172 ( 
.A1(n_167),
.A2(n_159),
.A3(n_165),
.B(n_161),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_1),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_10),
.C(n_5),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_162),
.A2(n_1),
.B(n_2),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_173),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_R g184 ( 
.A(n_172),
.B(n_175),
.C(n_4),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_158),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_178),
.B(n_181),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_169),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_10),
.C(n_6),
.Y(n_181)
);

NOR2xp67_ASAP7_75t_SL g182 ( 
.A(n_172),
.B(n_174),
.Y(n_182)
);

AOI21xp33_ASAP7_75t_L g187 ( 
.A1(n_182),
.A2(n_184),
.B(n_4),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_4),
.C(n_6),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_168),
.C(n_7),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_179),
.A2(n_176),
.B(n_173),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_189),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_190),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_187),
.A2(n_7),
.B(n_9),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_7),
.Y(n_189)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_191),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_168),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_188),
.C(n_9),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_192),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_194),
.C(n_196),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_198),
.Y(n_200)
);


endmodule