module fake_ariane_1977_n_156 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_41, n_38, n_2, n_18, n_32, n_28, n_37, n_9, n_11, n_34, n_26, n_3, n_14, n_0, n_36, n_33, n_19, n_30, n_39, n_40, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_156);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_41;
input n_38;
input n_2;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_11;
input n_34;
input n_26;
input n_3;
input n_14;
input n_0;
input n_36;
input n_33;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_156;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_124;
wire n_119;
wire n_90;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_149;
wire n_69;
wire n_95;
wire n_92;
wire n_143;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_152;
wire n_120;
wire n_106;
wire n_53;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_49;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_82;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_52;
wire n_135;
wire n_73;
wire n_77;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_125;
wire n_43;
wire n_81;
wire n_87;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_54;

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_22),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_33),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_13),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_4),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_29),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_6),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_10),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_37),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_46),
.B(n_0),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_0),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_3),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_3),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

AND2x4_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_45),
.B(n_5),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_9),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_45),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_11),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_85),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_67),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_59),
.B(n_50),
.Y(n_93)
);

AOI21x1_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_12),
.B(n_15),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_66),
.B(n_63),
.C(n_53),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_59),
.B(n_48),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_69),
.B(n_75),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_17),
.Y(n_101)
);

CKINVDCx5p33_ASAP7_75t_R g102 ( 
.A(n_90),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_80),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_73),
.B(n_71),
.C(n_82),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_80),
.B(n_69),
.Y(n_106)
);

AND2x4_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_71),
.Y(n_107)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_94),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_82),
.B1(n_88),
.B2(n_85),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_79),
.Y(n_110)
);

NOR2xp67_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_77),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_89),
.A2(n_78),
.B(n_20),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_78),
.B(n_21),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_78),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_19),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_101),
.B1(n_95),
.B2(n_99),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

OAI21x1_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_25),
.B(n_28),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_30),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_105),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_118),
.A2(n_109),
.B1(n_104),
.B2(n_114),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_121),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_105),
.Y(n_131)
);

NAND3xp33_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_106),
.C(n_103),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_115),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_122),
.Y(n_134)
);

OAI221xp5_ASAP7_75t_SL g135 ( 
.A1(n_124),
.A2(n_104),
.B1(n_113),
.B2(n_35),
.C(n_36),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_116),
.A2(n_31),
.B1(n_34),
.B2(n_38),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_119),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

AND2x4_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_119),
.Y(n_142)
);

INVxp67_ASAP7_75t_SL g143 ( 
.A(n_139),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_140),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_135),
.C(n_136),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_133),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_144),
.Y(n_148)
);

NAND4xp75_ASAP7_75t_L g149 ( 
.A(n_147),
.B(n_146),
.C(n_138),
.D(n_145),
.Y(n_149)
);

NAND3xp33_ASAP7_75t_L g150 ( 
.A(n_148),
.B(n_138),
.C(n_142),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_149),
.A2(n_142),
.B1(n_148),
.B2(n_127),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

OAI21x1_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_150),
.B(n_152),
.Y(n_155)
);

OAI221xp5_ASAP7_75t_R g156 ( 
.A1(n_155),
.A2(n_152),
.B1(n_39),
.B2(n_125),
.C(n_127),
.Y(n_156)
);


endmodule