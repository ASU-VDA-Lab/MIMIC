module fake_jpeg_22533_n_333 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_L g42 ( 
.A1(n_19),
.A2(n_9),
.B(n_15),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_35),
.B1(n_18),
.B2(n_29),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_45),
.Y(n_76)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_25),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx5_ASAP7_75t_SL g56 ( 
.A(n_48),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_49),
.B(n_35),
.Y(n_55)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_31),
.Y(n_57)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_20),
.B1(n_37),
.B2(n_36),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_58),
.A2(n_61),
.B1(n_63),
.B2(n_65),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_46),
.A2(n_17),
.B1(n_20),
.B2(n_32),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_17),
.B1(n_32),
.B2(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_37),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_64),
.B(n_81),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_17),
.B1(n_32),
.B2(n_21),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_68),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_49),
.Y(n_99)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_27),
.B1(n_35),
.B2(n_33),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_51),
.B1(n_29),
.B2(n_40),
.Y(n_88)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_80),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_26),
.B1(n_24),
.B2(n_27),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_71),
.A2(n_28),
.B1(n_36),
.B2(n_30),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_27),
.B1(n_18),
.B2(n_33),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_78),
.A2(n_30),
.B1(n_28),
.B2(n_44),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_31),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_40),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_83),
.Y(n_122)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_51),
.A2(n_27),
.B1(n_48),
.B2(n_40),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_23),
.B1(n_38),
.B2(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_87),
.B(n_93),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_88),
.A2(n_95),
.B1(n_60),
.B2(n_66),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_89),
.B(n_99),
.Y(n_127)
);

OR2x2_ASAP7_75t_SL g90 ( 
.A(n_67),
.B(n_26),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_90),
.A2(n_98),
.B(n_114),
.Y(n_153)
);

AO22x2_ASAP7_75t_SL g91 ( 
.A1(n_85),
.A2(n_47),
.B1(n_48),
.B2(n_39),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_91),
.A2(n_116),
.B1(n_117),
.B2(n_119),
.Y(n_124)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

HAxp5_ASAP7_75t_SL g98 ( 
.A(n_76),
.B(n_39),
.CON(n_98),
.SN(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_78),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_100),
.Y(n_150)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_104),
.Y(n_140)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_49),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_105),
.B(n_115),
.Y(n_142)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_109),
.Y(n_143)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_60),
.A2(n_26),
.B1(n_48),
.B2(n_47),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_113),
.A2(n_59),
.B1(n_44),
.B2(n_54),
.Y(n_149)
);

AO22x1_ASAP7_75t_L g114 ( 
.A1(n_71),
.A2(n_47),
.B1(n_23),
.B2(n_38),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_82),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_49),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_13),
.Y(n_120)
);

OR2x6_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_34),
.Y(n_145)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_108),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_132),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_83),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_155),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_39),
.C(n_74),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_39),
.C(n_80),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_103),
.A2(n_59),
.B1(n_68),
.B2(n_70),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_129),
.A2(n_106),
.B1(n_109),
.B2(n_94),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_86),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_96),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_139),
.Y(n_168)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_136),
.B(n_137),
.Y(n_177)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_149),
.B1(n_94),
.B2(n_97),
.Y(n_171)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_144),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_145),
.A2(n_104),
.B(n_54),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_146),
.B(n_151),
.Y(n_179)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g148 ( 
.A(n_90),
.B(n_39),
.C(n_44),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_38),
.C(n_34),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_113),
.Y(n_152)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_120),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_154),
.Y(n_180)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_158),
.Y(n_164)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_93),
.Y(n_157)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_62),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_186),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_173),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_165),
.A2(n_174),
.B1(n_149),
.B2(n_157),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_166),
.A2(n_169),
.B(n_182),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_116),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_170),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_153),
.A2(n_107),
.B(n_110),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_77),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_171),
.A2(n_175),
.B1(n_178),
.B2(n_191),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_62),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_181),
.Y(n_202)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_151),
.A2(n_92),
.B1(n_97),
.B2(n_73),
.Y(n_174)
);

AO21x2_ASAP7_75t_L g175 ( 
.A1(n_141),
.A2(n_77),
.B(n_102),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_SL g221 ( 
.A1(n_176),
.A2(n_190),
.B(n_0),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_158),
.A2(n_38),
.B1(n_102),
.B2(n_34),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_126),
.B(n_34),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_0),
.B(n_1),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_188),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_137),
.A2(n_0),
.B(n_1),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_148),
.A2(n_34),
.B(n_22),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_123),
.B(n_22),
.C(n_1),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_134),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_145),
.A2(n_22),
.B(n_1),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_144),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_145),
.A2(n_7),
.B(n_15),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

OAI21x1_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_145),
.B(n_176),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_195),
.A2(n_221),
.B(n_192),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_199),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_187),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_200),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_129),
.B1(n_146),
.B2(n_124),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_201),
.A2(n_218),
.B1(n_223),
.B2(n_174),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_182),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_203),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_167),
.A2(n_145),
.B1(n_142),
.B2(n_132),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_210),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_175),
.A2(n_145),
.B1(n_133),
.B2(n_136),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_175),
.A2(n_156),
.B1(n_131),
.B2(n_135),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_159),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_209),
.Y(n_236)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_177),
.Y(n_211)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_161),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_212),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_160),
.C(n_181),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_175),
.A2(n_131),
.B1(n_155),
.B2(n_135),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_214),
.A2(n_215),
.B1(n_191),
.B2(n_190),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_184),
.A2(n_147),
.B1(n_139),
.B2(n_130),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_216),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_217),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_183),
.A2(n_6),
.B1(n_14),
.B2(n_3),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_161),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_164),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_165),
.Y(n_222)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_222),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_179),
.A2(n_2),
.B(n_4),
.C(n_10),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_227),
.A2(n_199),
.B1(n_208),
.B2(n_197),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_228),
.A2(n_242),
.B(n_197),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_166),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_229),
.A2(n_194),
.B(n_223),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_244),
.C(n_213),
.Y(n_249)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_207),
.A2(n_164),
.B1(n_170),
.B2(n_178),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_235),
.A2(n_247),
.B1(n_200),
.B2(n_216),
.Y(n_263)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_193),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_239),
.Y(n_261)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_162),
.Y(n_240)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_198),
.B(n_185),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_243),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_203),
.A2(n_188),
.B(n_186),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_202),
.B(n_169),
.C(n_180),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_245),
.A2(n_220),
.B1(n_196),
.B2(n_211),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_214),
.A2(n_173),
.B1(n_189),
.B2(n_2),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_250),
.C(n_254),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_202),
.C(n_198),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_236),
.B(n_210),
.Y(n_251)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_252),
.A2(n_232),
.B(n_229),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_204),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_262),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_204),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_256),
.A2(n_265),
.B1(n_245),
.B2(n_224),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_220),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_264),
.C(n_248),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_259),
.A2(n_267),
.B(n_232),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_260),
.A2(n_266),
.B1(n_227),
.B2(n_243),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_205),
.Y(n_262)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_234),
.C(n_240),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_233),
.A2(n_2),
.B1(n_4),
.B2(n_10),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_233),
.A2(n_12),
.B1(n_14),
.B2(n_16),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_12),
.Y(n_268)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_268),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_273),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_279),
.C(n_254),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_274),
.A2(n_226),
.B(n_263),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_275),
.A2(n_282),
.B(n_259),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_246),
.C(n_225),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_261),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_281),
.Y(n_289)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

FAx1_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_229),
.CI(n_224),
.CON(n_282),
.SN(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_246),
.Y(n_283)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_283),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_250),
.B(n_237),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_226),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_225),
.Y(n_285)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_285),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_247),
.Y(n_286)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_286),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_288),
.A2(n_293),
.B1(n_283),
.B2(n_275),
.Y(n_307)
);

XOR2x2_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_262),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_271),
.B1(n_286),
.B2(n_273),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_296),
.C(n_270),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_299),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_276),
.A2(n_239),
.B1(n_266),
.B2(n_238),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_295),
.A2(n_269),
.B1(n_282),
.B2(n_265),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_230),
.C(n_238),
.Y(n_296)
);

INVx13_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_277),
.B(n_253),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_277),
.Y(n_306)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_301),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_230),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_302),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_296),
.B(n_272),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_305),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_304),
.A2(n_308),
.B(n_309),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_278),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_307),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_270),
.C(n_274),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_298),
.B1(n_290),
.B2(n_287),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_311),
.B(n_313),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_297),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_300),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_306),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_319),
.A2(n_321),
.B(n_323),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_317),
.A2(n_289),
.B(n_288),
.Y(n_320)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_320),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_314),
.A2(n_289),
.B(n_298),
.Y(n_321)
);

OAI21xp33_ASAP7_75t_L g322 ( 
.A1(n_315),
.A2(n_291),
.B(n_293),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_316),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_324),
.A2(n_325),
.B(n_304),
.Y(n_328)
);

NAND4xp25_ASAP7_75t_SL g327 ( 
.A(n_326),
.B(n_312),
.C(n_295),
.D(n_316),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_328),
.C(n_287),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_290),
.B(n_311),
.Y(n_330)
);

AOI21x1_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_286),
.B(n_318),
.Y(n_331)
);

O2A1O1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_235),
.B(n_12),
.C(n_16),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_16),
.Y(n_333)
);


endmodule