module fake_netlist_1_8186_n_667 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_667);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_667;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_482;
wire n_394;
wire n_243;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_L g78 ( .A(n_66), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_21), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_33), .Y(n_80) );
INVxp33_ASAP7_75t_SL g81 ( .A(n_34), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_61), .Y(n_82) );
INVxp67_ASAP7_75t_SL g83 ( .A(n_32), .Y(n_83) );
BUFx6f_ASAP7_75t_L g84 ( .A(n_77), .Y(n_84) );
BUFx3_ASAP7_75t_L g85 ( .A(n_73), .Y(n_85) );
INVxp33_ASAP7_75t_SL g86 ( .A(n_46), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_45), .Y(n_87) );
BUFx2_ASAP7_75t_L g88 ( .A(n_8), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_65), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_13), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_42), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_7), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_28), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_43), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_19), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_3), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_6), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_29), .Y(n_98) );
HB1xp67_ASAP7_75t_L g99 ( .A(n_20), .Y(n_99) );
INVxp33_ASAP7_75t_L g100 ( .A(n_44), .Y(n_100) );
INVxp33_ASAP7_75t_SL g101 ( .A(n_41), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_21), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_52), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_38), .Y(n_104) );
INVxp33_ASAP7_75t_SL g105 ( .A(n_53), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_67), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_18), .Y(n_107) );
INVxp67_ASAP7_75t_SL g108 ( .A(n_72), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_17), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_39), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_22), .Y(n_111) );
INVx1_ASAP7_75t_SL g112 ( .A(n_62), .Y(n_112) );
INVxp67_ASAP7_75t_L g113 ( .A(n_37), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_74), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_4), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_68), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_49), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_71), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_5), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_27), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_4), .Y(n_121) );
HB1xp67_ASAP7_75t_L g122 ( .A(n_57), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_76), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_70), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_50), .Y(n_125) );
INVxp33_ASAP7_75t_L g126 ( .A(n_19), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_84), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_102), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_122), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_106), .Y(n_130) );
NOR2xp33_ASAP7_75t_R g131 ( .A(n_106), .B(n_25), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_120), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_122), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_120), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_109), .Y(n_135) );
INVx4_ASAP7_75t_L g136 ( .A(n_85), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_88), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_109), .Y(n_138) );
NOR2xp33_ASAP7_75t_R g139 ( .A(n_87), .B(n_75), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_88), .Y(n_140) );
INVxp67_ASAP7_75t_L g141 ( .A(n_99), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_118), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_119), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_99), .B(n_0), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_103), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_84), .B(n_0), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_81), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_85), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_126), .B(n_113), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_109), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_113), .B(n_1), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_84), .Y(n_152) );
BUFx8_ASAP7_75t_L g153 ( .A(n_103), .Y(n_153) );
CKINVDCx6p67_ASAP7_75t_R g154 ( .A(n_85), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_86), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_101), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_121), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_84), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_84), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_125), .B(n_1), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_105), .Y(n_161) );
INVx1_ASAP7_75t_SL g162 ( .A(n_78), .Y(n_162) );
BUFx3_ASAP7_75t_L g163 ( .A(n_125), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_121), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_121), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_80), .B(n_2), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_103), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_79), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_79), .Y(n_169) );
AND2x2_ASAP7_75t_L g170 ( .A(n_100), .B(n_2), .Y(n_170) );
INVxp67_ASAP7_75t_L g171 ( .A(n_92), .Y(n_171) );
NOR2xp67_ASAP7_75t_L g172 ( .A(n_92), .B(n_3), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_169), .Y(n_173) );
AOI22xp33_ASAP7_75t_L g174 ( .A1(n_169), .A2(n_95), .B1(n_96), .B2(n_97), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_163), .B(n_124), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_169), .Y(n_176) );
AND2x6_ASAP7_75t_L g177 ( .A(n_144), .B(n_124), .Y(n_177) );
AOI22x1_ASAP7_75t_L g178 ( .A1(n_136), .A2(n_83), .B1(n_108), .B2(n_116), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_163), .Y(n_179) );
NAND2x1p5_ASAP7_75t_L g180 ( .A(n_144), .B(n_97), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_145), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_129), .B(n_123), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_136), .B(n_123), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_162), .B(n_111), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_145), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_149), .B(n_117), .Y(n_186) );
INVx2_ASAP7_75t_SL g187 ( .A(n_154), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_136), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_167), .Y(n_189) );
INVxp67_ASAP7_75t_SL g190 ( .A(n_141), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_167), .Y(n_191) );
XNOR2xp5_ASAP7_75t_L g192 ( .A(n_128), .B(n_90), .Y(n_192) );
OR2x2_ASAP7_75t_L g193 ( .A(n_140), .B(n_90), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_164), .Y(n_194) );
OR2x6_ASAP7_75t_L g195 ( .A(n_137), .B(n_96), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_133), .B(n_111), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g197 ( .A1(n_168), .A2(n_95), .B1(n_115), .B2(n_107), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_165), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_135), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_154), .B(n_117), .Y(n_200) );
AND2x6_ASAP7_75t_L g201 ( .A(n_170), .B(n_116), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_135), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_171), .B(n_94), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_147), .B(n_94), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_138), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_153), .B(n_98), .Y(n_206) );
BUFx2_ASAP7_75t_L g207 ( .A(n_143), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_153), .B(n_98), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_138), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_148), .B(n_115), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_142), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_150), .Y(n_212) );
BUFx4f_ASAP7_75t_L g213 ( .A(n_170), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_150), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_157), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_157), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_166), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_172), .Y(n_218) );
INVx2_ASAP7_75t_SL g219 ( .A(n_153), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_151), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_160), .Y(n_221) );
AND2x6_ASAP7_75t_L g222 ( .A(n_127), .B(n_80), .Y(n_222) );
AO22x2_ASAP7_75t_L g223 ( .A1(n_146), .A2(n_107), .B1(n_83), .B2(n_108), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_140), .Y(n_224) );
AND2x6_ASAP7_75t_L g225 ( .A(n_127), .B(n_114), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_143), .B(n_114), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_131), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_127), .Y(n_228) );
OAI22xp5_ASAP7_75t_SL g229 ( .A1(n_142), .A2(n_91), .B1(n_110), .B2(n_104), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_127), .Y(n_230) );
AND2x4_ASAP7_75t_L g231 ( .A(n_130), .B(n_91), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_130), .B(n_110), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_173), .Y(n_233) );
BUFx2_ASAP7_75t_L g234 ( .A(n_207), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_197), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_173), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_176), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_180), .Y(n_238) );
BUFx2_ASAP7_75t_L g239 ( .A(n_190), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_211), .Y(n_240) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_219), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_220), .B(n_161), .Y(n_242) );
INVx5_ASAP7_75t_L g243 ( .A(n_222), .Y(n_243) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_208), .A2(n_82), .B(n_104), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_217), .B(n_161), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_190), .B(n_134), .Y(n_246) );
INVx3_ASAP7_75t_L g247 ( .A(n_205), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_203), .B(n_134), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_180), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_203), .B(n_132), .Y(n_250) );
AND3x2_ASAP7_75t_SL g251 ( .A(n_192), .B(n_132), .C(n_147), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_221), .B(n_156), .Y(n_252) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_222), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_199), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_202), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_197), .Y(n_256) );
OR2x2_ASAP7_75t_SL g257 ( .A(n_193), .B(n_155), .Y(n_257) );
INVx3_ASAP7_75t_L g258 ( .A(n_209), .Y(n_258) );
INVx2_ASAP7_75t_SL g259 ( .A(n_213), .Y(n_259) );
AND2x6_ASAP7_75t_L g260 ( .A(n_196), .B(n_82), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_222), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_212), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_200), .B(n_156), .Y(n_263) );
OR2x2_ASAP7_75t_L g264 ( .A(n_184), .B(n_155), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_214), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_232), .B(n_112), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_177), .A2(n_89), .B1(n_93), .B2(n_112), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_215), .Y(n_268) );
OR2x6_ASAP7_75t_L g269 ( .A(n_195), .B(n_93), .Y(n_269) );
OR2x6_ASAP7_75t_L g270 ( .A(n_195), .B(n_89), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_200), .B(n_139), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_216), .Y(n_272) );
BUFx2_ASAP7_75t_L g273 ( .A(n_177), .Y(n_273) );
BUFx10_ASAP7_75t_L g274 ( .A(n_187), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_222), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_177), .A2(n_84), .B1(n_158), .B2(n_152), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_208), .B(n_159), .Y(n_277) );
INVxp67_ASAP7_75t_L g278 ( .A(n_210), .Y(n_278) );
NOR2xp33_ASAP7_75t_R g279 ( .A(n_224), .B(n_5), .Y(n_279) );
NOR3xp33_ASAP7_75t_SL g280 ( .A(n_229), .B(n_6), .C(n_7), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_213), .B(n_159), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_177), .B(n_159), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_195), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_177), .B(n_159), .Y(n_284) );
NOR2xp33_ASAP7_75t_R g285 ( .A(n_227), .B(n_8), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_210), .Y(n_286) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_222), .Y(n_287) );
INVxp67_ASAP7_75t_L g288 ( .A(n_231), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_194), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_188), .Y(n_290) );
AND2x6_ASAP7_75t_L g291 ( .A(n_196), .B(n_159), .Y(n_291) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_225), .Y(n_292) );
NOR3xp33_ASAP7_75t_SL g293 ( .A(n_204), .B(n_9), .C(n_10), .Y(n_293) );
BUFx2_ASAP7_75t_L g294 ( .A(n_201), .Y(n_294) );
BUFx2_ASAP7_75t_L g295 ( .A(n_201), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_232), .B(n_9), .Y(n_296) );
NOR2xp33_ASAP7_75t_SL g297 ( .A(n_231), .B(n_158), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_181), .Y(n_298) );
AO22x1_ASAP7_75t_L g299 ( .A1(n_201), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_258), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_239), .B(n_226), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_277), .A2(n_206), .B(n_183), .Y(n_302) );
NAND2x1p5_ASAP7_75t_L g303 ( .A(n_238), .B(n_226), .Y(n_303) );
INVx2_ASAP7_75t_SL g304 ( .A(n_269), .Y(n_304) );
AOI21x1_ASAP7_75t_L g305 ( .A1(n_282), .A2(n_183), .B(n_175), .Y(n_305) );
A2O1A1Ixp33_ASAP7_75t_SL g306 ( .A1(n_266), .A2(n_204), .B(n_182), .C(n_218), .Y(n_306) );
AND2x4_ASAP7_75t_L g307 ( .A(n_249), .B(n_201), .Y(n_307) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_253), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_268), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_245), .B(n_186), .Y(n_310) );
BUFx12f_ASAP7_75t_L g311 ( .A(n_234), .Y(n_311) );
CKINVDCx11_ASAP7_75t_R g312 ( .A(n_235), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_269), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_269), .Y(n_314) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_253), .Y(n_315) );
A2O1A1Ixp33_ASAP7_75t_L g316 ( .A1(n_293), .A2(n_175), .B(n_189), .C(n_185), .Y(n_316) );
INVx2_ASAP7_75t_SL g317 ( .A(n_269), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_256), .B(n_174), .Y(n_318) );
INVx3_ASAP7_75t_L g319 ( .A(n_298), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_242), .B(n_201), .Y(n_320) );
AOI221x1_ASAP7_75t_L g321 ( .A1(n_284), .A2(n_223), .B1(n_198), .B2(n_191), .C(n_127), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_260), .B(n_179), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_253), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_260), .B(n_174), .Y(n_324) );
BUFx2_ASAP7_75t_L g325 ( .A(n_270), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_260), .A2(n_223), .B1(n_178), .B2(n_225), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_253), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_298), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_240), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_260), .A2(n_223), .B1(n_225), .B2(n_158), .Y(n_330) );
BUFx2_ASAP7_75t_L g331 ( .A(n_270), .Y(n_331) );
BUFx3_ASAP7_75t_L g332 ( .A(n_291), .Y(n_332) );
CKINVDCx11_ASAP7_75t_R g333 ( .A(n_235), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g334 ( .A1(n_260), .A2(n_225), .B1(n_158), .B2(n_152), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_261), .Y(n_335) );
INVx8_ASAP7_75t_L g336 ( .A(n_270), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_289), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_283), .B(n_158), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_298), .Y(n_339) );
INVx2_ASAP7_75t_SL g340 ( .A(n_270), .Y(n_340) );
OR2x6_ASAP7_75t_L g341 ( .A(n_273), .B(n_152), .Y(n_341) );
AND2x4_ASAP7_75t_L g342 ( .A(n_259), .B(n_11), .Y(n_342) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_261), .Y(n_343) );
AND2x6_ASAP7_75t_L g344 ( .A(n_241), .B(n_152), .Y(n_344) );
BUFx2_ASAP7_75t_L g345 ( .A(n_286), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g346 ( .A(n_240), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g347 ( .A(n_294), .B(n_152), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_260), .B(n_225), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_296), .B(n_12), .Y(n_349) );
NAND2xp5_ASAP7_75t_SL g350 ( .A(n_295), .B(n_230), .Y(n_350) );
INVx6_ASAP7_75t_SL g351 ( .A(n_274), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_258), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_258), .Y(n_353) );
OR2x6_ASAP7_75t_L g354 ( .A(n_259), .B(n_13), .Y(n_354) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_261), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_318), .A2(n_256), .B1(n_296), .B2(n_254), .Y(n_356) );
A2O1A1Ixp33_ASAP7_75t_L g357 ( .A1(n_316), .A2(n_262), .B(n_265), .C(n_272), .Y(n_357) );
CKINVDCx11_ASAP7_75t_R g358 ( .A(n_311), .Y(n_358) );
AND2x4_ASAP7_75t_SL g359 ( .A(n_313), .B(n_274), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_337), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_310), .A2(n_265), .B1(n_262), .B2(n_255), .Y(n_361) );
OAI211xp5_ASAP7_75t_SL g362 ( .A1(n_312), .A2(n_280), .B(n_278), .C(n_252), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_310), .A2(n_255), .B1(n_254), .B2(n_272), .Y(n_363) );
INVxp67_ASAP7_75t_L g364 ( .A(n_345), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_336), .A2(n_267), .B1(n_286), .B2(n_288), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_301), .B(n_264), .Y(n_366) );
OAI222xp33_ASAP7_75t_L g367 ( .A1(n_354), .A2(n_251), .B1(n_246), .B2(n_248), .C1(n_250), .C2(n_263), .Y(n_367) );
INVx8_ASAP7_75t_L g368 ( .A(n_336), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_336), .A2(n_257), .B1(n_247), .B2(n_271), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_309), .B(n_291), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_303), .B(n_251), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_303), .B(n_279), .Y(n_372) );
NAND3xp33_ASAP7_75t_SL g373 ( .A(n_346), .B(n_279), .C(n_285), .Y(n_373) );
INVx3_ASAP7_75t_L g374 ( .A(n_336), .Y(n_374) );
NAND2x1_ASAP7_75t_L g375 ( .A(n_344), .B(n_291), .Y(n_375) );
OAI22xp33_ASAP7_75t_L g376 ( .A1(n_354), .A2(n_297), .B1(n_241), .B2(n_247), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_304), .B(n_291), .Y(n_377) );
INVx4_ASAP7_75t_L g378 ( .A(n_314), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_349), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_311), .Y(n_380) );
INVx6_ASAP7_75t_L g381 ( .A(n_307), .Y(n_381) );
OAI21xp5_ASAP7_75t_L g382 ( .A1(n_302), .A2(n_237), .B(n_290), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_342), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_342), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_317), .B(n_291), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_320), .A2(n_291), .B1(n_241), .B2(n_244), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_340), .B(n_244), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_324), .A2(n_247), .B1(n_241), .B2(n_237), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_342), .A2(n_244), .B1(n_233), .B2(n_285), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_320), .B(n_274), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_325), .A2(n_236), .B1(n_299), .B2(n_233), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_360), .Y(n_392) );
AOI22xp33_ASAP7_75t_SL g393 ( .A1(n_369), .A2(n_346), .B1(n_354), .B2(n_331), .Y(n_393) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_375), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_370), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_362), .A2(n_333), .B1(n_312), .B2(n_329), .Y(n_396) );
BUFx3_ASAP7_75t_L g397 ( .A(n_368), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_383), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_356), .A2(n_333), .B1(n_329), .B2(n_307), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_356), .B(n_307), .Y(n_400) );
AOI22xp33_ASAP7_75t_SL g401 ( .A1(n_368), .A2(n_332), .B1(n_328), .B2(n_319), .Y(n_401) );
AND2x4_ASAP7_75t_L g402 ( .A(n_374), .B(n_319), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_373), .A2(n_330), .B1(n_326), .B2(n_319), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_371), .B(n_306), .Y(n_404) );
OA21x2_ASAP7_75t_L g405 ( .A1(n_357), .A2(n_321), .B(n_316), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_366), .A2(n_306), .B1(n_339), .B2(n_281), .C(n_328), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_384), .Y(n_407) );
OAI22xp33_ASAP7_75t_L g408 ( .A1(n_368), .A2(n_351), .B1(n_328), .B2(n_352), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_379), .Y(n_409) );
OAI21xp5_ASAP7_75t_L g410 ( .A1(n_357), .A2(n_305), .B(n_353), .Y(n_410) );
OAI22xp33_ASAP7_75t_L g411 ( .A1(n_365), .A2(n_351), .B1(n_353), .B2(n_352), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_382), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_372), .A2(n_351), .B1(n_300), .B2(n_281), .Y(n_413) );
CKINVDCx8_ASAP7_75t_R g414 ( .A(n_380), .Y(n_414) );
OAI21x1_ASAP7_75t_L g415 ( .A1(n_388), .A2(n_300), .B(n_350), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_361), .A2(n_363), .B1(n_390), .B2(n_391), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_361), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_367), .A2(n_322), .B1(n_338), .B2(n_290), .C(n_347), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_363), .B(n_332), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_387), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_392), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_392), .B(n_389), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_392), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_393), .A2(n_390), .B1(n_389), .B2(n_378), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_397), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_417), .B(n_374), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_409), .A2(n_364), .B1(n_376), .B2(n_378), .C(n_359), .Y(n_427) );
INVx2_ASAP7_75t_SL g428 ( .A(n_397), .Y(n_428) );
INVx1_ASAP7_75t_SL g429 ( .A(n_420), .Y(n_429) );
INVxp67_ASAP7_75t_L g430 ( .A(n_404), .Y(n_430) );
OAI33xp33_ASAP7_75t_L g431 ( .A1(n_404), .A2(n_338), .A3(n_385), .B1(n_377), .B2(n_347), .B3(n_350), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_420), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_400), .A2(n_381), .B1(n_358), .B2(n_359), .Y(n_433) );
AO21x2_ASAP7_75t_L g434 ( .A1(n_410), .A2(n_386), .B(n_334), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_409), .B(n_420), .Y(n_435) );
NAND3xp33_ASAP7_75t_L g436 ( .A(n_406), .B(n_276), .C(n_341), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_398), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_398), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_412), .Y(n_439) );
OAI221xp5_ASAP7_75t_L g440 ( .A1(n_399), .A2(n_381), .B1(n_348), .B2(n_341), .C(n_358), .Y(n_440) );
INVxp67_ASAP7_75t_SL g441 ( .A(n_411), .Y(n_441) );
OAI22xp33_ASAP7_75t_L g442 ( .A1(n_416), .A2(n_381), .B1(n_341), .B2(n_343), .Y(n_442) );
AOI222xp33_ASAP7_75t_L g443 ( .A1(n_396), .A2(n_344), .B1(n_15), .B2(n_16), .C1(n_17), .C2(n_18), .Y(n_443) );
AOI211xp5_ASAP7_75t_L g444 ( .A1(n_408), .A2(n_261), .B(n_275), .C(n_287), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_407), .Y(n_445) );
AOI21x1_ASAP7_75t_L g446 ( .A1(n_405), .A2(n_341), .B(n_228), .Y(n_446) );
OAI221xp5_ASAP7_75t_L g447 ( .A1(n_416), .A2(n_355), .B1(n_343), .B2(n_335), .C(n_327), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_410), .A2(n_355), .B(n_308), .Y(n_448) );
NAND4xp25_ASAP7_75t_L g449 ( .A(n_406), .B(n_14), .C(n_15), .D(n_16), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_417), .B(n_14), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_400), .B(n_20), .Y(n_451) );
INVx3_ASAP7_75t_L g452 ( .A(n_394), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_407), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_395), .B(n_22), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_395), .Y(n_455) );
NOR3xp33_ASAP7_75t_L g456 ( .A(n_449), .B(n_418), .C(n_401), .Y(n_456) );
INVx1_ASAP7_75t_SL g457 ( .A(n_429), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_432), .B(n_412), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_432), .B(n_394), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_440), .B(n_414), .Y(n_460) );
NAND4xp25_ASAP7_75t_L g461 ( .A(n_443), .B(n_418), .C(n_403), .D(n_413), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_432), .Y(n_462) );
NAND4xp25_ASAP7_75t_L g463 ( .A(n_443), .B(n_397), .C(n_419), .D(n_401), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_452), .B(n_439), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_435), .B(n_419), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_429), .B(n_405), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_421), .B(n_405), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_425), .Y(n_468) );
INVx4_ASAP7_75t_L g469 ( .A(n_452), .Y(n_469) );
AOI21xp33_ASAP7_75t_L g470 ( .A1(n_441), .A2(n_405), .B(n_394), .Y(n_470) );
NAND3xp33_ASAP7_75t_L g471 ( .A(n_430), .B(n_394), .C(n_402), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_423), .B(n_415), .Y(n_472) );
OAI31xp33_ASAP7_75t_L g473 ( .A1(n_449), .A2(n_402), .A3(n_24), .B(n_23), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_435), .Y(n_474) );
INVx3_ASAP7_75t_L g475 ( .A(n_452), .Y(n_475) );
INVx3_ASAP7_75t_L g476 ( .A(n_452), .Y(n_476) );
INVx1_ASAP7_75t_SL g477 ( .A(n_428), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_451), .A2(n_402), .B1(n_344), .B2(n_415), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_428), .B(n_394), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_423), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_439), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_439), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_422), .B(n_438), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_422), .B(n_394), .Y(n_484) );
INVx2_ASAP7_75t_SL g485 ( .A(n_450), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_437), .Y(n_486) );
INVx4_ASAP7_75t_L g487 ( .A(n_450), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_437), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_438), .B(n_402), .Y(n_489) );
OAI221xp5_ASAP7_75t_L g490 ( .A1(n_424), .A2(n_433), .B1(n_427), .B2(n_444), .C(n_426), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_445), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_451), .B(n_23), .Y(n_492) );
INVx2_ASAP7_75t_SL g493 ( .A(n_426), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_455), .B(n_344), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_455), .B(n_344), .Y(n_495) );
AND2x2_ASAP7_75t_SL g496 ( .A(n_454), .B(n_323), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_445), .Y(n_497) );
AOI33xp33_ASAP7_75t_L g498 ( .A1(n_453), .A2(n_24), .A3(n_414), .B1(n_30), .B2(n_31), .B3(n_35), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_453), .B(n_26), .Y(n_499) );
NOR2x1_ASAP7_75t_SL g500 ( .A(n_454), .B(n_355), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_434), .B(n_36), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_446), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_434), .B(n_40), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_483), .B(n_434), .Y(n_504) );
INVx2_ASAP7_75t_SL g505 ( .A(n_468), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_488), .Y(n_506) );
OR2x6_ASAP7_75t_L g507 ( .A(n_487), .B(n_448), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_486), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_474), .B(n_442), .Y(n_509) );
OR2x4_ASAP7_75t_L g510 ( .A(n_460), .B(n_431), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g511 ( .A1(n_463), .A2(n_436), .B1(n_444), .B2(n_434), .Y(n_511) );
INVx1_ASAP7_75t_SL g512 ( .A(n_477), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_483), .B(n_446), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_488), .B(n_436), .Y(n_514) );
NOR3xp33_ASAP7_75t_L g515 ( .A(n_498), .B(n_447), .C(n_48), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_489), .B(n_47), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_489), .B(n_51), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_486), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_486), .Y(n_519) );
OAI31xp33_ASAP7_75t_L g520 ( .A1(n_473), .A2(n_54), .A3(n_55), .B(n_56), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_484), .B(n_58), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_465), .B(n_59), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_480), .B(n_60), .Y(n_523) );
AOI22x1_ASAP7_75t_L g524 ( .A1(n_492), .A2(n_355), .B1(n_343), .B2(n_335), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_491), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_491), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_491), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_463), .B(n_63), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_492), .B(n_64), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_497), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_497), .Y(n_531) );
NOR2xp33_ASAP7_75t_R g532 ( .A(n_496), .B(n_69), .Y(n_532) );
OR2x6_ASAP7_75t_L g533 ( .A(n_487), .B(n_308), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_479), .A2(n_308), .B(n_335), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_484), .B(n_230), .Y(n_535) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_457), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_467), .B(n_464), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_471), .A2(n_315), .B(n_335), .Y(n_538) );
OR2x6_ASAP7_75t_L g539 ( .A(n_487), .B(n_343), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_462), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_461), .A2(n_327), .B1(n_323), .B2(n_315), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_487), .B(n_327), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_485), .B(n_315), .Y(n_543) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_499), .Y(n_544) );
NAND2xp33_ASAP7_75t_R g545 ( .A(n_501), .B(n_323), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_490), .B(n_230), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_490), .B(n_275), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_457), .B(n_275), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_458), .B(n_292), .Y(n_549) );
NAND2xp33_ASAP7_75t_SL g550 ( .A(n_501), .B(n_292), .Y(n_550) );
INVxp67_ASAP7_75t_SL g551 ( .A(n_536), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_528), .A2(n_456), .B1(n_461), .B2(n_493), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_506), .Y(n_553) );
INVx2_ASAP7_75t_SL g554 ( .A(n_505), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_540), .Y(n_555) );
OAI22xp33_ASAP7_75t_L g556 ( .A1(n_544), .A2(n_471), .B1(n_478), .B2(n_473), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_537), .B(n_464), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_544), .A2(n_456), .B1(n_478), .B2(n_493), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_537), .B(n_505), .Y(n_559) );
CKINVDCx16_ASAP7_75t_R g560 ( .A(n_532), .Y(n_560) );
NAND4xp25_ASAP7_75t_L g561 ( .A(n_528), .B(n_470), .C(n_503), .D(n_499), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_504), .B(n_493), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_512), .B(n_469), .Y(n_563) );
AOI222xp33_ASAP7_75t_L g564 ( .A1(n_504), .A2(n_509), .B1(n_546), .B2(n_547), .C1(n_514), .C2(n_513), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_521), .B(n_464), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_519), .Y(n_566) );
INVx1_ASAP7_75t_SL g567 ( .A(n_532), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_525), .Y(n_568) );
AOI221xp5_ASAP7_75t_L g569 ( .A1(n_547), .A2(n_482), .B1(n_481), .B2(n_472), .C(n_458), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_526), .B(n_482), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_521), .B(n_464), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_527), .Y(n_572) );
OR2x6_ASAP7_75t_L g573 ( .A(n_533), .B(n_469), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_540), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_530), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_508), .B(n_462), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_531), .B(n_462), .Y(n_577) );
AOI322xp5_ASAP7_75t_L g578 ( .A1(n_511), .A2(n_502), .A3(n_495), .B1(n_494), .B2(n_459), .C1(n_475), .C2(n_476), .Y(n_578) );
OAI22xp5_ASAP7_75t_SL g579 ( .A1(n_510), .A2(n_469), .B1(n_495), .B2(n_494), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_518), .B(n_466), .Y(n_580) );
NOR3xp33_ASAP7_75t_L g581 ( .A(n_515), .B(n_476), .C(n_475), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_518), .Y(n_582) );
NAND2xp33_ASAP7_75t_L g583 ( .A(n_529), .B(n_476), .Y(n_583) );
A2O1A1Ixp33_ASAP7_75t_L g584 ( .A1(n_520), .A2(n_475), .B(n_459), .C(n_466), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_545), .A2(n_459), .B1(n_502), .B2(n_500), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_535), .B(n_543), .Y(n_586) );
NOR2x1p5_ASAP7_75t_L g587 ( .A(n_522), .B(n_459), .Y(n_587) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_550), .A2(n_500), .B(n_287), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_523), .Y(n_589) );
INVx1_ASAP7_75t_SL g590 ( .A(n_542), .Y(n_590) );
NOR3xp33_ASAP7_75t_L g591 ( .A(n_516), .B(n_243), .C(n_517), .Y(n_591) );
NOR2x1_ASAP7_75t_L g592 ( .A(n_533), .B(n_243), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_553), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_564), .B(n_535), .Y(n_594) );
AOI21xp33_ASAP7_75t_SL g595 ( .A1(n_560), .A2(n_539), .B(n_533), .Y(n_595) );
CKINVDCx20_ASAP7_75t_R g596 ( .A(n_590), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_557), .B(n_507), .Y(n_597) );
NOR3xp33_ASAP7_75t_SL g598 ( .A(n_556), .B(n_549), .C(n_538), .Y(n_598) );
INVx1_ASAP7_75t_SL g599 ( .A(n_554), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_559), .B(n_539), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_555), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_562), .B(n_507), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_566), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_562), .B(n_507), .Y(n_604) );
INVxp67_ASAP7_75t_L g605 ( .A(n_551), .Y(n_605) );
OAI211xp5_ASAP7_75t_SL g606 ( .A1(n_552), .A2(n_541), .B(n_534), .C(n_507), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_574), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_565), .B(n_539), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_568), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_582), .Y(n_610) );
NOR3xp33_ASAP7_75t_L g611 ( .A(n_558), .B(n_548), .C(n_524), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_572), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_575), .Y(n_613) );
INVx1_ASAP7_75t_SL g614 ( .A(n_563), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_580), .B(n_586), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_563), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_571), .B(n_586), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_569), .B(n_589), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_576), .B(n_577), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_569), .B(n_558), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_577), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_578), .B(n_570), .Y(n_622) );
AOI221x1_ASAP7_75t_L g623 ( .A1(n_595), .A2(n_581), .B1(n_579), .B2(n_591), .C(n_561), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_615), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_615), .Y(n_625) );
AO22x1_ASAP7_75t_L g626 ( .A1(n_599), .A2(n_567), .B1(n_573), .B2(n_583), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_622), .B(n_584), .Y(n_627) );
XNOR2xp5_ASAP7_75t_L g628 ( .A(n_596), .B(n_587), .Y(n_628) );
OAI22x1_ASAP7_75t_SL g629 ( .A1(n_596), .A2(n_573), .B1(n_585), .B2(n_588), .Y(n_629) );
NOR2x1_ASAP7_75t_L g630 ( .A(n_606), .B(n_588), .Y(n_630) );
INVx2_ASAP7_75t_SL g631 ( .A(n_614), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_601), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_621), .Y(n_633) );
XNOR2xp5_ASAP7_75t_L g634 ( .A(n_594), .B(n_592), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_611), .A2(n_618), .B1(n_604), .B2(n_602), .Y(n_635) );
INVxp67_ASAP7_75t_L g636 ( .A(n_605), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_617), .B(n_602), .Y(n_637) );
XNOR2xp5_ASAP7_75t_L g638 ( .A(n_617), .B(n_597), .Y(n_638) );
NOR2x1_ASAP7_75t_L g639 ( .A(n_629), .B(n_616), .Y(n_639) );
AND2x4_ASAP7_75t_L g640 ( .A(n_636), .B(n_604), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_635), .A2(n_597), .B1(n_598), .B2(n_600), .Y(n_641) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_633), .Y(n_642) );
AOI322xp5_ASAP7_75t_L g643 ( .A1(n_627), .A2(n_593), .A3(n_608), .B1(n_612), .B2(n_603), .C1(n_609), .C2(n_613), .Y(n_643) );
CKINVDCx20_ASAP7_75t_R g644 ( .A(n_628), .Y(n_644) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_632), .Y(n_645) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_631), .Y(n_646) );
AO22x2_ASAP7_75t_L g647 ( .A1(n_623), .A2(n_619), .B1(n_610), .B2(n_607), .Y(n_647) );
NAND4xp25_ASAP7_75t_L g648 ( .A(n_630), .B(n_624), .C(n_625), .D(n_637), .Y(n_648) );
NAND4xp25_ASAP7_75t_L g649 ( .A(n_634), .B(n_623), .C(n_635), .D(n_630), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_638), .B(n_634), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g651 ( .A1(n_626), .A2(n_635), .B1(n_627), .B2(n_594), .C(n_629), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_638), .A2(n_635), .B1(n_628), .B2(n_596), .Y(n_652) );
OAI222xp33_ASAP7_75t_L g653 ( .A1(n_635), .A2(n_628), .B1(n_627), .B2(n_620), .C1(n_634), .C2(n_638), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_639), .B(n_647), .Y(n_654) );
CKINVDCx5p33_ASAP7_75t_R g655 ( .A(n_644), .Y(n_655) );
NAND2x1p5_ASAP7_75t_L g656 ( .A(n_645), .B(n_640), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_642), .Y(n_657) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_646), .Y(n_658) );
NOR3xp33_ASAP7_75t_L g659 ( .A(n_654), .B(n_649), .C(n_653), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_654), .A2(n_651), .B1(n_652), .B2(n_641), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_658), .B(n_643), .Y(n_661) );
OR2x2_ASAP7_75t_L g662 ( .A(n_661), .B(n_648), .Y(n_662) );
OR3x1_ASAP7_75t_L g663 ( .A(n_659), .B(n_657), .C(n_655), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_663), .Y(n_664) );
OAI21xp5_ASAP7_75t_L g665 ( .A1(n_662), .A2(n_660), .B(n_656), .Y(n_665) );
XNOR2xp5_ASAP7_75t_L g666 ( .A(n_664), .B(n_650), .Y(n_666) );
AOI21xp5_ASAP7_75t_L g667 ( .A1(n_666), .A2(n_665), .B(n_647), .Y(n_667) );
endmodule