module real_aes_7419_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_746;
wire n_153;
wire n_532;
wire n_284;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_283;
wire n_252;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g112 ( .A(n_0), .Y(n_112) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_1), .A2(n_148), .B(n_151), .C(n_226), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_2), .A2(n_176), .B(n_177), .Y(n_175) );
INVx1_ASAP7_75t_L g507 ( .A(n_3), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_4), .B(n_187), .Y(n_186) );
AOI21xp33_ASAP7_75t_L g484 ( .A1(n_5), .A2(n_176), .B(n_485), .Y(n_484) );
AND2x6_ASAP7_75t_L g148 ( .A(n_6), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g251 ( .A(n_7), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_8), .B(n_42), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_8), .B(n_42), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_9), .A2(n_275), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_10), .B(n_160), .Y(n_228) );
INVx1_ASAP7_75t_L g489 ( .A(n_11), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_12), .B(n_181), .Y(n_540) );
INVx1_ASAP7_75t_L g140 ( .A(n_13), .Y(n_140) );
INVx1_ASAP7_75t_L g552 ( .A(n_14), .Y(n_552) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_15), .A2(n_195), .B(n_236), .C(n_238), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_16), .B(n_187), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_17), .B(n_478), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_18), .B(n_176), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_19), .B(n_283), .Y(n_282) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_20), .A2(n_181), .B(n_212), .C(n_215), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_21), .B(n_187), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_22), .B(n_160), .Y(n_159) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_23), .A2(n_214), .B(n_238), .C(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_24), .B(n_160), .Y(n_196) );
CKINVDCx16_ASAP7_75t_R g142 ( .A(n_25), .Y(n_142) );
INVx1_ASAP7_75t_L g193 ( .A(n_26), .Y(n_193) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_27), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_28), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_29), .B(n_160), .Y(n_508) );
INVx1_ASAP7_75t_L g280 ( .A(n_30), .Y(n_280) );
INVx1_ASAP7_75t_L g497 ( .A(n_31), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g123 ( .A1(n_32), .A2(n_124), .B1(n_125), .B2(n_450), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_32), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_33), .A2(n_104), .B1(n_117), .B2(n_763), .Y(n_103) );
INVx2_ASAP7_75t_L g146 ( .A(n_34), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_35), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_36), .B(n_458), .Y(n_457) );
A2O1A1Ixp33_ASAP7_75t_L g180 ( .A1(n_37), .A2(n_181), .B(n_182), .C(n_184), .Y(n_180) );
INVxp67_ASAP7_75t_L g281 ( .A(n_38), .Y(n_281) );
CKINVDCx14_ASAP7_75t_R g178 ( .A(n_39), .Y(n_178) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_40), .A2(n_151), .B(n_192), .C(n_199), .Y(n_191) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_41), .A2(n_148), .B(n_151), .C(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g496 ( .A(n_43), .Y(n_496) );
OAI22xp5_ASAP7_75t_SL g447 ( .A1(n_44), .A2(n_52), .B1(n_448), .B2(n_449), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_44), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_45), .A2(n_65), .B1(n_753), .B2(n_754), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_45), .Y(n_754) );
OAI22xp5_ASAP7_75t_SL g750 ( .A1(n_46), .A2(n_751), .B1(n_752), .B2(n_755), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_46), .Y(n_755) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_47), .A2(n_162), .B(n_249), .C(n_250), .Y(n_248) );
AOI222xp33_ASAP7_75t_L g460 ( .A1(n_48), .A2(n_461), .B1(n_749), .B2(n_750), .C1(n_756), .C2(n_759), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_49), .B(n_160), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_50), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g277 ( .A(n_51), .Y(n_277) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_52), .Y(n_448) );
INVx1_ASAP7_75t_L g210 ( .A(n_53), .Y(n_210) );
CKINVDCx16_ASAP7_75t_R g498 ( .A(n_54), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_55), .B(n_176), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_56), .A2(n_151), .B1(n_215), .B2(n_495), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_57), .Y(n_523) );
CKINVDCx16_ASAP7_75t_R g504 ( .A(n_58), .Y(n_504) );
CKINVDCx14_ASAP7_75t_R g247 ( .A(n_59), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_60), .A2(n_184), .B(n_249), .C(n_488), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_61), .Y(n_532) );
INVx1_ASAP7_75t_L g486 ( .A(n_62), .Y(n_486) );
INVx1_ASAP7_75t_L g149 ( .A(n_63), .Y(n_149) );
INVx1_ASAP7_75t_L g139 ( .A(n_64), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_65), .Y(n_753) );
INVx1_ASAP7_75t_SL g183 ( .A(n_66), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_67), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_68), .B(n_187), .Y(n_217) );
INVx1_ASAP7_75t_L g155 ( .A(n_69), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_SL g477 ( .A1(n_70), .A2(n_184), .B(n_478), .C(n_479), .Y(n_477) );
INVxp67_ASAP7_75t_L g480 ( .A(n_71), .Y(n_480) );
INVx1_ASAP7_75t_L g116 ( .A(n_72), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_73), .A2(n_176), .B(n_246), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_74), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_75), .A2(n_176), .B(n_233), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_76), .Y(n_500) );
INVx1_ASAP7_75t_L g526 ( .A(n_77), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_78), .A2(n_275), .B(n_276), .Y(n_274) );
CKINVDCx16_ASAP7_75t_R g190 ( .A(n_79), .Y(n_190) );
INVx1_ASAP7_75t_L g234 ( .A(n_80), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_81), .A2(n_148), .B(n_151), .C(n_528), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_82), .A2(n_176), .B(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g237 ( .A(n_83), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_84), .B(n_194), .Y(n_520) );
INVx2_ASAP7_75t_L g137 ( .A(n_85), .Y(n_137) );
INVx1_ASAP7_75t_L g227 ( .A(n_86), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_87), .B(n_478), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_88), .A2(n_148), .B(n_151), .C(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g113 ( .A(n_89), .Y(n_113) );
OR2x2_ASAP7_75t_L g453 ( .A(n_89), .B(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g747 ( .A(n_89), .B(n_455), .Y(n_747) );
A2O1A1Ixp33_ASAP7_75t_L g150 ( .A1(n_90), .A2(n_151), .B(n_154), .C(n_164), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_91), .B(n_169), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_92), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_93), .A2(n_148), .B(n_151), .C(n_538), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_94), .Y(n_544) );
INVx1_ASAP7_75t_L g476 ( .A(n_95), .Y(n_476) );
CKINVDCx16_ASAP7_75t_R g549 ( .A(n_96), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_97), .B(n_194), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_98), .B(n_135), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_99), .B(n_135), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_100), .B(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g213 ( .A(n_101), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_102), .A2(n_176), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g763 ( .A(n_106), .Y(n_763) );
CKINVDCx9p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
CKINVDCx14_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_112), .B(n_113), .C(n_114), .Y(n_111) );
AND2x2_ASAP7_75t_L g455 ( .A(n_112), .B(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g464 ( .A(n_113), .B(n_455), .Y(n_464) );
NOR2x2_ASAP7_75t_L g758 ( .A(n_113), .B(n_454), .Y(n_758) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
AO21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_122), .B(n_459), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx3_ASAP7_75t_L g762 ( .A(n_119), .Y(n_762) );
INVx2_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI21xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_451), .B(n_457), .Y(n_122) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
XNOR2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_447), .Y(n_125) );
INVx3_ASAP7_75t_L g748 ( .A(n_126), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_126), .A2(n_463), .B1(n_746), .B2(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_SL g126 ( .A(n_127), .B(n_402), .Y(n_126) );
NOR4xp25_ASAP7_75t_L g127 ( .A(n_128), .B(n_339), .C(n_373), .D(n_389), .Y(n_127) );
NAND4xp25_ASAP7_75t_SL g128 ( .A(n_129), .B(n_265), .C(n_303), .D(n_319), .Y(n_128) );
AOI222xp33_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_202), .B1(n_240), .B2(n_253), .C1(n_258), .C2(n_264), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AOI31xp33_ASAP7_75t_L g435 ( .A1(n_131), .A2(n_436), .A3(n_437), .B(n_439), .Y(n_435) );
OR2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_170), .Y(n_131) );
AND2x2_ASAP7_75t_L g410 ( .A(n_132), .B(n_172), .Y(n_410) );
BUFx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_SL g257 ( .A(n_133), .Y(n_257) );
AND2x2_ASAP7_75t_L g264 ( .A(n_133), .B(n_188), .Y(n_264) );
AND2x2_ASAP7_75t_L g324 ( .A(n_133), .B(n_173), .Y(n_324) );
AO21x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_141), .B(n_166), .Y(n_133) );
INVx3_ASAP7_75t_L g187 ( .A(n_134), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_134), .B(n_201), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_134), .B(n_230), .Y(n_229) );
NOR2xp33_ASAP7_75t_SL g522 ( .A(n_134), .B(n_523), .Y(n_522) );
INVx4_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_135), .Y(n_174) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_135), .A2(n_474), .B(n_481), .Y(n_473) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g273 ( .A(n_136), .Y(n_273) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
AND2x2_ASAP7_75t_SL g169 ( .A(n_137), .B(n_138), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
OAI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_150), .Y(n_141) );
O2A1O1Ixp33_ASAP7_75t_L g189 ( .A1(n_143), .A2(n_169), .B(n_190), .C(n_191), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g223 ( .A1(n_143), .A2(n_224), .B(n_225), .Y(n_223) );
OAI22xp33_ASAP7_75t_L g493 ( .A1(n_143), .A2(n_165), .B1(n_494), .B2(n_498), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g503 ( .A1(n_143), .A2(n_504), .B(n_505), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_143), .A2(n_526), .B(n_527), .Y(n_525) );
NAND2x1p5_ASAP7_75t_L g143 ( .A(n_144), .B(n_148), .Y(n_143) );
AND2x4_ASAP7_75t_L g176 ( .A(n_144), .B(n_148), .Y(n_176) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
INVx1_ASAP7_75t_L g198 ( .A(n_145), .Y(n_198) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g152 ( .A(n_146), .Y(n_152) );
INVx1_ASAP7_75t_L g216 ( .A(n_146), .Y(n_216) );
INVx1_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_147), .Y(n_158) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_147), .Y(n_160) );
INVx3_ASAP7_75t_L g195 ( .A(n_147), .Y(n_195) );
INVx1_ASAP7_75t_L g478 ( .A(n_147), .Y(n_478) );
INVx4_ASAP7_75t_SL g165 ( .A(n_148), .Y(n_165) );
BUFx3_ASAP7_75t_L g199 ( .A(n_148), .Y(n_199) );
INVx5_ASAP7_75t_L g179 ( .A(n_151), .Y(n_179) );
AND2x6_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
BUFx3_ASAP7_75t_L g163 ( .A(n_152), .Y(n_163) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_152), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_159), .C(n_161), .Y(n_154) );
O2A1O1Ixp5_ASAP7_75t_L g226 ( .A1(n_156), .A2(n_161), .B(n_227), .C(n_228), .Y(n_226) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
OAI22xp5_ASAP7_75t_SL g495 ( .A1(n_157), .A2(n_158), .B1(n_496), .B2(n_497), .Y(n_495) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx4_ASAP7_75t_L g214 ( .A(n_158), .Y(n_214) );
INVx4_ASAP7_75t_L g181 ( .A(n_160), .Y(n_181) );
INVx2_ASAP7_75t_L g249 ( .A(n_160), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_161), .A2(n_520), .B(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_161), .A2(n_529), .B(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g238 ( .A(n_163), .Y(n_238) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_L g177 ( .A1(n_165), .A2(n_178), .B(n_179), .C(n_180), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_SL g209 ( .A1(n_165), .A2(n_179), .B(n_210), .C(n_211), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_SL g233 ( .A1(n_165), .A2(n_179), .B(n_234), .C(n_235), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_SL g246 ( .A1(n_165), .A2(n_179), .B(n_247), .C(n_248), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_SL g276 ( .A1(n_165), .A2(n_179), .B(n_277), .C(n_278), .Y(n_276) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_165), .A2(n_179), .B(n_476), .C(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g485 ( .A1(n_165), .A2(n_179), .B(n_486), .C(n_487), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_L g548 ( .A1(n_165), .A2(n_179), .B(n_549), .C(n_550), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
INVx1_ASAP7_75t_L g283 ( .A(n_168), .Y(n_283) );
AO21x2_ASAP7_75t_L g535 ( .A1(n_168), .A2(n_536), .B(n_543), .Y(n_535) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g222 ( .A(n_169), .Y(n_222) );
OA21x2_ASAP7_75t_L g244 ( .A1(n_169), .A2(n_245), .B(n_252), .Y(n_244) );
OA21x2_ASAP7_75t_L g546 ( .A1(n_169), .A2(n_547), .B(n_553), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_170), .B(n_354), .Y(n_353) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_171), .B(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_171), .B(n_268), .Y(n_314) );
AND2x2_ASAP7_75t_L g407 ( .A(n_171), .B(n_347), .Y(n_407) );
OAI321xp33_ASAP7_75t_L g441 ( .A1(n_171), .A2(n_257), .A3(n_414), .B1(n_442), .B2(n_444), .C(n_445), .Y(n_441) );
NAND4xp25_ASAP7_75t_L g445 ( .A(n_171), .B(n_243), .C(n_354), .D(n_446), .Y(n_445) );
AND2x4_ASAP7_75t_L g171 ( .A(n_172), .B(n_188), .Y(n_171) );
AND2x2_ASAP7_75t_L g309 ( .A(n_172), .B(n_255), .Y(n_309) );
AND2x2_ASAP7_75t_L g328 ( .A(n_172), .B(n_257), .Y(n_328) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g256 ( .A(n_173), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g284 ( .A(n_173), .B(n_188), .Y(n_284) );
AND2x2_ASAP7_75t_L g370 ( .A(n_173), .B(n_255), .Y(n_370) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_186), .Y(n_173) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_174), .A2(n_208), .B(n_217), .Y(n_207) );
OA21x2_ASAP7_75t_L g231 ( .A1(n_174), .A2(n_232), .B(n_239), .Y(n_231) );
BUFx2_ASAP7_75t_L g275 ( .A(n_176), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_181), .B(n_183), .Y(n_182) );
INVx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_185), .Y(n_541) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_187), .A2(n_484), .B(n_490), .Y(n_483) );
INVx3_ASAP7_75t_SL g255 ( .A(n_188), .Y(n_255) );
AND2x2_ASAP7_75t_L g302 ( .A(n_188), .B(n_289), .Y(n_302) );
OR2x2_ASAP7_75t_L g335 ( .A(n_188), .B(n_257), .Y(n_335) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_188), .Y(n_342) );
AND2x2_ASAP7_75t_L g371 ( .A(n_188), .B(n_256), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_188), .B(n_344), .Y(n_386) );
AND2x2_ASAP7_75t_L g418 ( .A(n_188), .B(n_410), .Y(n_418) );
AND2x2_ASAP7_75t_L g427 ( .A(n_188), .B(n_269), .Y(n_427) );
OR2x6_ASAP7_75t_L g188 ( .A(n_189), .B(n_200), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_196), .C(n_197), .Y(n_192) );
OAI22xp33_ASAP7_75t_L g279 ( .A1(n_194), .A2(n_214), .B1(n_280), .B2(n_281), .Y(n_279) );
O2A1O1Ixp33_ASAP7_75t_L g506 ( .A1(n_194), .A2(n_507), .B(n_508), .C(n_509), .Y(n_506) );
INVx5_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_195), .B(n_251), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_195), .B(n_480), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_195), .B(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_198), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_204), .B(n_218), .Y(n_203) );
INVx1_ASAP7_75t_SL g395 ( .A(n_204), .Y(n_395) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g260 ( .A(n_205), .B(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g242 ( .A(n_206), .B(n_220), .Y(n_242) );
AND2x2_ASAP7_75t_L g331 ( .A(n_206), .B(n_244), .Y(n_331) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g301 ( .A(n_207), .B(n_231), .Y(n_301) );
OR2x2_ASAP7_75t_L g312 ( .A(n_207), .B(n_244), .Y(n_312) );
AND2x2_ASAP7_75t_L g338 ( .A(n_207), .B(n_244), .Y(n_338) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_207), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_214), .B(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_214), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g509 ( .A(n_215), .Y(n_509) );
INVx3_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_218), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_218), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_SL g218 ( .A(n_219), .Y(n_218) );
OR2x2_ASAP7_75t_L g311 ( .A(n_219), .B(n_312), .Y(n_311) );
AOI322xp5_ASAP7_75t_L g397 ( .A1(n_219), .A2(n_301), .A3(n_307), .B1(n_338), .B2(n_388), .C1(n_398), .C2(n_400), .Y(n_397) );
OR2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_231), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_220), .B(n_243), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_220), .B(n_244), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_220), .B(n_261), .Y(n_318) );
AND2x2_ASAP7_75t_L g372 ( .A(n_220), .B(n_338), .Y(n_372) );
INVx1_ASAP7_75t_L g376 ( .A(n_220), .Y(n_376) );
AND2x2_ASAP7_75t_L g388 ( .A(n_220), .B(n_231), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_220), .B(n_260), .Y(n_420) );
INVx4_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g285 ( .A(n_221), .B(n_231), .Y(n_285) );
BUFx3_ASAP7_75t_L g299 ( .A(n_221), .Y(n_299) );
AND3x2_ASAP7_75t_L g381 ( .A(n_221), .B(n_361), .C(n_382), .Y(n_381) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_229), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_222), .B(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_222), .B(n_532), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_222), .B(n_544), .Y(n_543) );
NAND3xp33_ASAP7_75t_L g241 ( .A(n_231), .B(n_242), .C(n_243), .Y(n_241) );
INVx1_ASAP7_75t_SL g261 ( .A(n_231), .Y(n_261) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_231), .Y(n_366) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g360 ( .A(n_242), .B(n_361), .Y(n_360) );
INVxp67_ASAP7_75t_L g367 ( .A(n_242), .Y(n_367) );
AND2x2_ASAP7_75t_L g405 ( .A(n_243), .B(n_383), .Y(n_405) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
BUFx3_ASAP7_75t_L g286 ( .A(n_244), .Y(n_286) );
AND2x2_ASAP7_75t_L g361 ( .A(n_244), .B(n_261), .Y(n_361) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
OR2x2_ASAP7_75t_L g305 ( .A(n_255), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g424 ( .A(n_255), .B(n_324), .Y(n_424) );
AND2x2_ASAP7_75t_L g438 ( .A(n_255), .B(n_257), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_256), .B(n_269), .Y(n_379) );
AND2x2_ASAP7_75t_L g426 ( .A(n_256), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g289 ( .A(n_257), .B(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g306 ( .A(n_257), .B(n_269), .Y(n_306) );
INVx1_ASAP7_75t_L g316 ( .A(n_257), .Y(n_316) );
AND2x2_ASAP7_75t_L g347 ( .A(n_257), .B(n_269), .Y(n_347) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OAI221xp5_ASAP7_75t_L g389 ( .A1(n_259), .A2(n_390), .B1(n_394), .B2(n_396), .C(n_397), .Y(n_389) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_260), .B(n_262), .Y(n_259) );
AND2x2_ASAP7_75t_L g293 ( .A(n_260), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_263), .B(n_300), .Y(n_443) );
AOI322xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_285), .A3(n_286), .B1(n_287), .B2(n_293), .C1(n_295), .C2(n_302), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_284), .Y(n_267) );
NAND2x1p5_ASAP7_75t_L g323 ( .A(n_268), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_268), .B(n_334), .Y(n_333) );
O2A1O1Ixp33_ASAP7_75t_L g357 ( .A1(n_268), .A2(n_284), .B(n_358), .C(n_359), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_268), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_268), .B(n_328), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_268), .B(n_410), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_268), .B(n_438), .Y(n_437) );
BUFx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_269), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_269), .B(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g399 ( .A(n_269), .B(n_286), .Y(n_399) );
OA21x2_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_274), .B(n_282), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AO21x2_ASAP7_75t_L g290 ( .A1(n_271), .A2(n_291), .B(n_292), .Y(n_290) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_271), .A2(n_525), .B(n_531), .Y(n_524) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AOI21xp5_ASAP7_75t_SL g516 ( .A1(n_272), .A2(n_517), .B(n_518), .Y(n_516) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_273), .A2(n_493), .B(n_499), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_273), .B(n_500), .Y(n_499) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_273), .A2(n_503), .B(n_510), .Y(n_502) );
INVx1_ASAP7_75t_L g291 ( .A(n_274), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_282), .Y(n_292) );
INVx1_ASAP7_75t_L g374 ( .A(n_284), .Y(n_374) );
OAI31xp33_ASAP7_75t_L g384 ( .A1(n_284), .A2(n_309), .A3(n_385), .B(n_387), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_284), .B(n_290), .Y(n_436) );
INVx1_ASAP7_75t_SL g297 ( .A(n_285), .Y(n_297) );
AND2x2_ASAP7_75t_L g330 ( .A(n_285), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g411 ( .A(n_285), .B(n_412), .Y(n_411) );
OR2x2_ASAP7_75t_L g296 ( .A(n_286), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g321 ( .A(n_286), .Y(n_321) );
AND2x2_ASAP7_75t_L g348 ( .A(n_286), .B(n_301), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_286), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g440 ( .A(n_286), .B(n_388), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_288), .B(n_358), .Y(n_431) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g327 ( .A(n_290), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_SL g345 ( .A(n_290), .Y(n_345) );
NAND2xp33_ASAP7_75t_SL g295 ( .A(n_296), .B(n_298), .Y(n_295) );
OAI211xp5_ASAP7_75t_SL g339 ( .A1(n_297), .A2(n_340), .B(n_346), .C(n_362), .Y(n_339) );
OR2x2_ASAP7_75t_L g414 ( .A(n_297), .B(n_395), .Y(n_414) );
OR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
CKINVDCx16_ASAP7_75t_R g351 ( .A(n_299), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_299), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g320 ( .A(n_301), .B(n_321), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_307), .B(n_310), .C(n_313), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_SL g354 ( .A(n_306), .Y(n_354) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_309), .B(n_347), .Y(n_352) );
INVx1_ASAP7_75t_L g358 ( .A(n_309), .Y(n_358) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g317 ( .A(n_312), .B(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g350 ( .A(n_312), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g412 ( .A(n_312), .Y(n_412) );
AOI21xp33_ASAP7_75t_SL g313 ( .A1(n_314), .A2(n_315), .B(n_317), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_315), .A2(n_326), .B(n_329), .Y(n_325) );
AOI211xp5_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_322), .B(n_325), .C(n_332), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_320), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_323), .B(n_414), .Y(n_413) );
INVx2_ASAP7_75t_SL g336 ( .A(n_324), .Y(n_336) );
OAI21xp5_ASAP7_75t_L g391 ( .A1(n_326), .A2(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_331), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g356 ( .A(n_331), .Y(n_356) );
AOI21xp33_ASAP7_75t_SL g332 ( .A1(n_333), .A2(n_336), .B(n_337), .Y(n_332) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g387 ( .A(n_338), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_344), .B(n_370), .Y(n_396) );
AND2x2_ASAP7_75t_L g409 ( .A(n_344), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g423 ( .A(n_344), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g433 ( .A(n_344), .B(n_371), .Y(n_433) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI211xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_348), .B(n_349), .C(n_357), .Y(n_346) );
INVx1_ASAP7_75t_L g393 ( .A(n_347), .Y(n_393) );
OAI22xp33_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_352), .B1(n_353), .B2(n_355), .Y(n_349) );
OR2x2_ASAP7_75t_L g355 ( .A(n_351), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_351), .B(n_412), .Y(n_434) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g428 ( .A(n_361), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_368), .B1(n_371), .B2(n_372), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
INVx1_ASAP7_75t_L g446 ( .A(n_366), .Y(n_446) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g392 ( .A(n_370), .Y(n_392) );
OAI211xp5_ASAP7_75t_SL g373 ( .A1(n_374), .A2(n_375), .B(n_377), .C(n_384), .Y(n_373) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx2_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
INVxp67_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVxp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_392), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NOR5xp2_ASAP7_75t_L g402 ( .A(n_403), .B(n_421), .C(n_429), .D(n_435), .E(n_441), .Y(n_402) );
OAI211xp5_ASAP7_75t_SL g403 ( .A1(n_404), .A2(n_406), .B(n_408), .C(n_415), .Y(n_403) );
INVxp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_411), .B(n_413), .Y(n_408) );
OAI21xp33_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_418), .B(n_419), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_418), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AOI21xp33_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_425), .B(n_428), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_SL g444 ( .A(n_424), .Y(n_444) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_432), .B(n_434), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g458 ( .A(n_453), .Y(n_458) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AOI21xp33_ASAP7_75t_L g459 ( .A1(n_457), .A2(n_460), .B(n_762), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_465), .B1(n_746), .B2(n_748), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g761 ( .A(n_465), .Y(n_761) );
INVx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND4x1_ASAP7_75t_L g466 ( .A(n_467), .B(n_664), .C(n_711), .D(n_731), .Y(n_466) );
NOR3xp33_ASAP7_75t_SL g467 ( .A(n_468), .B(n_594), .C(n_619), .Y(n_467) );
OAI211xp5_ASAP7_75t_SL g468 ( .A1(n_469), .A2(n_512), .B(n_554), .C(n_584), .Y(n_468) );
INVxp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_491), .Y(n_470) );
INVx3_ASAP7_75t_SL g636 ( .A(n_471), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_471), .B(n_567), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_471), .B(n_501), .Y(n_717) );
AND2x2_ASAP7_75t_L g740 ( .A(n_471), .B(n_606), .Y(n_740) );
AND2x4_ASAP7_75t_L g471 ( .A(n_472), .B(n_482), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g558 ( .A(n_473), .B(n_483), .Y(n_558) );
INVx3_ASAP7_75t_L g571 ( .A(n_473), .Y(n_571) );
AND2x2_ASAP7_75t_L g576 ( .A(n_473), .B(n_482), .Y(n_576) );
OR2x2_ASAP7_75t_L g627 ( .A(n_473), .B(n_568), .Y(n_627) );
BUFx2_ASAP7_75t_L g647 ( .A(n_473), .Y(n_647) );
AND2x2_ASAP7_75t_L g657 ( .A(n_473), .B(n_568), .Y(n_657) );
AND2x2_ASAP7_75t_L g663 ( .A(n_473), .B(n_492), .Y(n_663) );
INVx1_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_483), .B(n_568), .Y(n_582) );
INVx2_ASAP7_75t_L g592 ( .A(n_483), .Y(n_592) );
AND2x2_ASAP7_75t_L g605 ( .A(n_483), .B(n_571), .Y(n_605) );
OR2x2_ASAP7_75t_L g616 ( .A(n_483), .B(n_568), .Y(n_616) );
AND2x2_ASAP7_75t_SL g662 ( .A(n_483), .B(n_663), .Y(n_662) );
BUFx2_ASAP7_75t_L g674 ( .A(n_483), .Y(n_674) );
AND2x2_ASAP7_75t_L g720 ( .A(n_483), .B(n_492), .Y(n_720) );
INVx3_ASAP7_75t_SL g593 ( .A(n_491), .Y(n_593) );
OR2x2_ASAP7_75t_L g646 ( .A(n_491), .B(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_501), .Y(n_491) );
INVx3_ASAP7_75t_L g568 ( .A(n_492), .Y(n_568) );
AND2x2_ASAP7_75t_L g635 ( .A(n_492), .B(n_502), .Y(n_635) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_492), .Y(n_703) );
AOI33xp33_ASAP7_75t_L g707 ( .A1(n_492), .A2(n_636), .A3(n_643), .B1(n_652), .B2(n_708), .B3(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g556 ( .A(n_501), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_501), .B(n_571), .Y(n_570) );
NOR3xp33_ASAP7_75t_L g630 ( .A(n_501), .B(n_631), .C(n_633), .Y(n_630) );
AND2x2_ASAP7_75t_L g656 ( .A(n_501), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_501), .B(n_663), .Y(n_666) );
AND2x2_ASAP7_75t_L g719 ( .A(n_501), .B(n_720), .Y(n_719) );
INVx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx3_ASAP7_75t_L g575 ( .A(n_502), .Y(n_575) );
OR2x2_ASAP7_75t_L g669 ( .A(n_502), .B(n_568), .Y(n_669) );
OR2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_533), .Y(n_512) );
AOI32xp33_ASAP7_75t_L g620 ( .A1(n_513), .A2(n_621), .A3(n_623), .B1(n_625), .B2(n_628), .Y(n_620) );
NOR2xp67_ASAP7_75t_L g693 ( .A(n_513), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g723 ( .A(n_513), .Y(n_723) );
INVx4_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g655 ( .A(n_514), .B(n_639), .Y(n_655) );
AND2x2_ASAP7_75t_L g675 ( .A(n_514), .B(n_601), .Y(n_675) );
AND2x2_ASAP7_75t_L g743 ( .A(n_514), .B(n_661), .Y(n_743) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_524), .Y(n_514) );
INVx3_ASAP7_75t_L g564 ( .A(n_515), .Y(n_564) );
AND2x2_ASAP7_75t_L g578 ( .A(n_515), .B(n_562), .Y(n_578) );
OR2x2_ASAP7_75t_L g583 ( .A(n_515), .B(n_561), .Y(n_583) );
INVx1_ASAP7_75t_L g590 ( .A(n_515), .Y(n_590) );
AND2x2_ASAP7_75t_L g598 ( .A(n_515), .B(n_572), .Y(n_598) );
AND2x2_ASAP7_75t_L g600 ( .A(n_515), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_515), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g653 ( .A(n_515), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_515), .B(n_738), .Y(n_737) );
OR2x6_ASAP7_75t_L g515 ( .A(n_516), .B(n_522), .Y(n_515) );
INVx2_ASAP7_75t_L g562 ( .A(n_524), .Y(n_562) );
AND2x2_ASAP7_75t_L g608 ( .A(n_524), .B(n_534), .Y(n_608) );
AND2x2_ASAP7_75t_L g618 ( .A(n_524), .B(n_546), .Y(n_618) );
INVx2_ASAP7_75t_L g738 ( .A(n_533), .Y(n_738) );
OR2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_545), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_534), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g579 ( .A(n_534), .Y(n_579) );
AND2x2_ASAP7_75t_L g623 ( .A(n_534), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g639 ( .A(n_534), .B(n_602), .Y(n_639) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g587 ( .A(n_535), .Y(n_587) );
AND2x2_ASAP7_75t_L g601 ( .A(n_535), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g652 ( .A(n_535), .B(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_535), .B(n_562), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_542), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_540), .B(n_541), .Y(n_538) );
AND2x2_ASAP7_75t_L g563 ( .A(n_545), .B(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g624 ( .A(n_545), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_545), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g661 ( .A(n_545), .Y(n_661) );
INVx1_ASAP7_75t_L g694 ( .A(n_545), .Y(n_694) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g572 ( .A(n_546), .B(n_562), .Y(n_572) );
INVx1_ASAP7_75t_L g602 ( .A(n_546), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_559), .B1(n_565), .B2(n_572), .C(n_573), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_556), .B(n_576), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_556), .B(n_639), .Y(n_716) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_558), .B(n_606), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_558), .B(n_567), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_558), .B(n_581), .Y(n_710) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g632 ( .A(n_562), .Y(n_632) );
AND2x2_ASAP7_75t_L g607 ( .A(n_563), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g685 ( .A(n_563), .Y(n_685) );
AND2x2_ASAP7_75t_L g617 ( .A(n_564), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_564), .B(n_587), .Y(n_633) );
AND2x2_ASAP7_75t_L g697 ( .A(n_564), .B(n_623), .Y(n_697) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
BUFx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g606 ( .A(n_568), .B(n_575), .Y(n_606) );
AND2x2_ASAP7_75t_L g702 ( .A(n_569), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_571), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_572), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_572), .B(n_579), .Y(n_667) );
AND2x2_ASAP7_75t_L g687 ( .A(n_572), .B(n_587), .Y(n_687) );
AND2x2_ASAP7_75t_L g708 ( .A(n_572), .B(n_652), .Y(n_708) );
OAI32xp33_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_577), .A3(n_579), .B1(n_580), .B2(n_583), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx1_ASAP7_75t_SL g581 ( .A(n_575), .Y(n_581) );
NAND2x1_ASAP7_75t_L g622 ( .A(n_575), .B(n_605), .Y(n_622) );
OR2x2_ASAP7_75t_L g626 ( .A(n_575), .B(n_627), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_575), .B(n_674), .Y(n_727) );
INVx1_ASAP7_75t_L g595 ( .A(n_576), .Y(n_595) );
OAI221xp5_ASAP7_75t_SL g713 ( .A1(n_577), .A2(n_668), .B1(n_714), .B2(n_717), .C(n_718), .Y(n_713) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g585 ( .A(n_578), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g628 ( .A(n_578), .B(n_601), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_578), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g706 ( .A(n_578), .B(n_639), .Y(n_706) );
INVxp67_ASAP7_75t_L g642 ( .A(n_579), .Y(n_642) );
OR2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
AND2x2_ASAP7_75t_L g712 ( .A(n_581), .B(n_699), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_581), .B(n_662), .Y(n_735) );
INVx1_ASAP7_75t_L g610 ( .A(n_583), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_583), .B(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g728 ( .A(n_583), .B(n_729), .Y(n_728) );
OAI21xp5_ASAP7_75t_SL g584 ( .A1(n_585), .A2(n_588), .B(n_591), .Y(n_584) );
AND2x2_ASAP7_75t_L g597 ( .A(n_586), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g681 ( .A(n_590), .B(n_601), .Y(n_681) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
AND2x2_ASAP7_75t_L g699 ( .A(n_592), .B(n_657), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_592), .B(n_656), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_593), .B(n_605), .Y(n_679) );
OAI211xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B(n_599), .C(n_609), .Y(n_594) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_595), .A2(n_630), .B1(n_634), .B2(n_637), .C(n_640), .Y(n_629) );
AOI31xp33_ASAP7_75t_L g724 ( .A1(n_595), .A2(n_725), .A3(n_726), .B(n_728), .Y(n_724) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_603), .B1(n_605), .B2(n_607), .Y(n_599) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx1_ASAP7_75t_L g725 ( .A(n_605), .Y(n_725) );
INVx1_ASAP7_75t_L g688 ( .A(n_606), .Y(n_688) );
O2A1O1Ixp33_ASAP7_75t_L g731 ( .A1(n_608), .A2(n_732), .B(n_734), .C(n_736), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B1(n_613), .B2(n_617), .Y(n_609) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_614), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OAI221xp5_ASAP7_75t_SL g704 ( .A1(n_616), .A2(n_650), .B1(n_669), .B2(n_705), .C(n_707), .Y(n_704) );
INVx1_ASAP7_75t_L g700 ( .A(n_617), .Y(n_700) );
INVx1_ASAP7_75t_L g654 ( .A(n_618), .Y(n_654) );
NAND3xp33_ASAP7_75t_SL g619 ( .A(n_620), .B(n_629), .C(n_644), .Y(n_619) );
OAI21xp33_ASAP7_75t_L g670 ( .A1(n_621), .A2(n_671), .B(n_675), .Y(n_670) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_623), .B(n_723), .Y(n_722) );
INVxp67_ASAP7_75t_L g730 ( .A(n_624), .Y(n_730) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g668 ( .A(n_631), .B(n_651), .Y(n_668) );
INVx1_ASAP7_75t_L g643 ( .A(n_632), .Y(n_643) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g641 ( .A(n_635), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_635), .B(n_673), .Y(n_672) );
NOR4xp25_ASAP7_75t_L g640 ( .A(n_636), .B(n_641), .C(n_642), .D(n_643), .Y(n_640) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AOI222xp33_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_649), .B1(n_655), .B2(n_656), .C1(n_658), .C2(n_662), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_646), .B(n_648), .Y(n_645) );
INVx1_ASAP7_75t_L g742 ( .A(n_646), .Y(n_742) );
INVx1_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_654), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_658), .B(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OAI21xp5_ASAP7_75t_SL g718 ( .A1(n_663), .A2(n_719), .B(n_721), .Y(n_718) );
NOR4xp25_ASAP7_75t_L g664 ( .A(n_665), .B(n_676), .C(n_689), .D(n_704), .Y(n_664) );
OAI221xp5_ASAP7_75t_SL g665 ( .A1(n_666), .A2(n_667), .B1(n_668), .B2(n_669), .C(n_670), .Y(n_665) );
INVx1_ASAP7_75t_L g745 ( .A(n_666), .Y(n_745) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_673), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
OAI222xp33_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_680), .B1(n_682), .B2(n_683), .C1(n_686), .C2(n_688), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AOI211xp5_ASAP7_75t_L g711 ( .A1(n_681), .A2(n_712), .B(n_713), .C(n_724), .Y(n_711) );
OR2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
INVx1_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
OAI222xp33_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_695), .B1(n_696), .B2(n_698), .C1(n_700), .C2(n_701), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVxp67_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_706), .A2(n_709), .B1(n_742), .B2(n_743), .Y(n_741) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
OAI211xp5_ASAP7_75t_SL g736 ( .A1(n_737), .A2(n_739), .B(n_741), .C(n_744), .Y(n_736) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx3_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
endmodule