module fake_jpeg_124_n_353 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_353);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_353;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_11),
.B(n_7),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_43),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_14),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_52),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_16),
.B(n_20),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_47),
.B(n_51),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_48),
.Y(n_116)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_16),
.B(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_15),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_54),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_57),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_30),
.B(n_15),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_27),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_74),
.Y(n_87)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_20),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_64),
.B(n_73),
.Y(n_114)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_0),
.Y(n_68)
);

AND2x4_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_31),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

NAND2xp33_ASAP7_75t_SL g109 ( 
.A(n_70),
.B(n_71),
.Y(n_109)
);

CKINVDCx6p67_ASAP7_75t_R g71 ( 
.A(n_35),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_34),
.B(n_18),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_38),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_18),
.B(n_10),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_76),
.B(n_77),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_36),
.B(n_13),
.Y(n_77)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_24),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_88),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_24),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_68),
.A2(n_62),
.B1(n_72),
.B2(n_44),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_90),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_68),
.A2(n_41),
.B1(n_19),
.B2(n_26),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_94),
.A2(n_107),
.B1(n_123),
.B2(n_60),
.Y(n_129)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_32),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_97),
.B(n_104),
.Y(n_140)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_45),
.A2(n_18),
.B1(n_21),
.B2(n_17),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_113),
.B1(n_121),
.B2(n_66),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_32),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_71),
.A2(n_38),
.B1(n_23),
.B2(n_39),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_105),
.A2(n_110),
.B1(n_115),
.B2(n_117),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_48),
.A2(n_41),
.B1(n_19),
.B2(n_26),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_71),
.A2(n_38),
.B1(n_23),
.B2(n_39),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_111),
.Y(n_151)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_67),
.A2(n_17),
.B1(n_21),
.B2(n_26),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_71),
.A2(n_38),
.B1(n_23),
.B2(n_31),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_61),
.A2(n_63),
.B1(n_38),
.B2(n_28),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_61),
.A2(n_40),
.B1(n_28),
.B2(n_26),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_70),
.A2(n_41),
.B1(n_19),
.B2(n_40),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_59),
.A2(n_35),
.B1(n_13),
.B2(n_2),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_129),
.A2(n_165),
.B1(n_143),
.B2(n_151),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_131),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_63),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_139),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_133),
.A2(n_146),
.B1(n_154),
.B2(n_160),
.Y(n_177)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

INVx13_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_55),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_136),
.B(n_153),
.Y(n_202)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_91),
.Y(n_138)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_138),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_80),
.B(n_0),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_84),
.B(n_1),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_150),
.Y(n_172)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_142),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_88),
.A2(n_55),
.B1(n_2),
.B2(n_3),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_147),
.B(n_109),
.Y(n_174)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g190 ( 
.A(n_149),
.Y(n_190)
);

NOR2x1_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_1),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_120),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_86),
.A2(n_90),
.B1(n_104),
.B2(n_97),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_3),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_156),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_120),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_159),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_123),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_161),
.A2(n_79),
.B(n_81),
.Y(n_197)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_82),
.Y(n_163)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_78),
.Y(n_164)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_164),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_94),
.A2(n_100),
.B1(n_112),
.B2(n_107),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_85),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_83),
.Y(n_198)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_119),
.Y(n_167)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_83),
.Y(n_168)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_92),
.C(n_103),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_169),
.B(n_187),
.C(n_206),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_134),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_188),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_174),
.B(n_175),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_140),
.B(n_111),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_176),
.A2(n_130),
.B1(n_202),
.B2(n_174),
.Y(n_214)
);

AND2x6_ASAP7_75t_L g185 ( 
.A(n_136),
.B(n_111),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_185),
.B(n_203),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_137),
.B(n_98),
.C(n_99),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_109),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_146),
.B(n_93),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_189),
.B(n_119),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_131),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_193),
.Y(n_231)
);

INVxp33_ASAP7_75t_L g193 ( 
.A(n_127),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_147),
.B(n_100),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_142),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_163),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_198),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_129),
.A2(n_106),
.B1(n_116),
.B2(n_124),
.Y(n_201)
);

A2O1A1Ixp33_ASAP7_75t_SL g223 ( 
.A1(n_201),
.A2(n_128),
.B(n_158),
.C(n_124),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_137),
.B(n_108),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_162),
.B(n_93),
.C(n_108),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_177),
.A2(n_130),
.B1(n_161),
.B2(n_165),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_208),
.A2(n_219),
.B1(n_223),
.B2(n_227),
.Y(n_258)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_210),
.Y(n_242)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_211),
.Y(n_260)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_196),
.Y(n_212)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_213),
.Y(n_245)
);

OA22x2_ASAP7_75t_L g253 ( 
.A1(n_214),
.A2(n_216),
.B1(n_173),
.B2(n_159),
.Y(n_253)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_190),
.A2(n_160),
.B1(n_149),
.B2(n_135),
.Y(n_216)
);

AOI21x1_ASAP7_75t_L g247 ( 
.A1(n_218),
.A2(n_181),
.B(n_195),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_177),
.A2(n_171),
.B1(n_176),
.B2(n_189),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_169),
.B(n_128),
.C(n_127),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_232),
.C(n_178),
.Y(n_240)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_194),
.A2(n_166),
.B1(n_156),
.B2(n_153),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_222),
.A2(n_237),
.B(n_180),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_225),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_175),
.B(n_164),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_126),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_233),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_201),
.A2(n_116),
.B1(n_106),
.B2(n_145),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_187),
.B(n_144),
.C(n_168),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_170),
.B(n_126),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_192),
.B(n_144),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_234),
.B(n_235),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_206),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_238),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_185),
.A2(n_148),
.B(n_138),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_197),
.B(n_157),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_172),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_264),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_240),
.B(n_251),
.C(n_252),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_224),
.A2(n_186),
.B1(n_179),
.B2(n_181),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_243),
.A2(n_231),
.B1(n_210),
.B2(n_227),
.Y(n_282)
);

AND2x2_ASAP7_75t_SL g246 ( 
.A(n_218),
.B(n_236),
.Y(n_246)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_246),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_247),
.A2(n_231),
.B(n_222),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_214),
.A2(n_181),
.B1(n_179),
.B2(n_173),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_249),
.A2(n_254),
.B1(n_261),
.B2(n_218),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_178),
.C(n_204),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_204),
.C(n_182),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_229),
.A2(n_182),
.B1(n_183),
.B2(n_200),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_200),
.C(n_205),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_259),
.C(n_212),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_205),
.C(n_180),
.Y(n_259)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_207),
.Y(n_263)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_263),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_234),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_261),
.A2(n_237),
.B(n_238),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_266),
.A2(n_279),
.B(n_286),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_275),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_265),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_284),
.C(n_257),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_219),
.Y(n_270)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_270),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_265),
.B(n_209),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_276),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_255),
.B(n_209),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_280),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_225),
.Y(n_274)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_252),
.B(n_251),
.Y(n_276)
);

NOR3xp33_ASAP7_75t_SL g277 ( 
.A(n_241),
.B(n_230),
.C(n_233),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_278),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_228),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_247),
.A2(n_230),
.B(n_226),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_256),
.B(n_235),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_282),
.A2(n_258),
.B1(n_254),
.B2(n_243),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_249),
.A2(n_213),
.B(n_208),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_287),
.A2(n_301),
.B1(n_268),
.B2(n_286),
.Y(n_307)
);

AOI322xp5_ASAP7_75t_L g292 ( 
.A1(n_270),
.A2(n_262),
.A3(n_246),
.B1(n_253),
.B2(n_258),
.C1(n_263),
.C2(n_242),
.Y(n_292)
);

OAI322xp33_ASAP7_75t_L g311 ( 
.A1(n_292),
.A2(n_300),
.A3(n_302),
.B1(n_281),
.B2(n_274),
.C1(n_285),
.C2(n_277),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_267),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_280),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_283),
.C(n_284),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_276),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_298),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_246),
.Y(n_298)
);

AOI322xp5_ASAP7_75t_L g300 ( 
.A1(n_267),
.A2(n_253),
.A3(n_242),
.B1(n_241),
.B2(n_245),
.C1(n_244),
.C2(n_250),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_271),
.A2(n_259),
.B1(n_253),
.B2(n_250),
.Y(n_301)
);

AOI322xp5_ASAP7_75t_L g302 ( 
.A1(n_278),
.A2(n_245),
.A3(n_244),
.B1(n_248),
.B2(n_260),
.C1(n_221),
.C2(n_223),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_266),
.A2(n_223),
.B1(n_248),
.B2(n_260),
.Y(n_303)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_303),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_312),
.C(n_314),
.Y(n_320)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_306),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_290),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_293),
.B(n_294),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_309),
.B(n_313),
.Y(n_321)
);

OAI21x1_ASAP7_75t_L g310 ( 
.A1(n_294),
.A2(n_299),
.B(n_281),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_316),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_311),
.A2(n_317),
.B1(n_289),
.B2(n_295),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_272),
.C(n_279),
.Y(n_312)
);

OA21x2_ASAP7_75t_SL g313 ( 
.A1(n_299),
.A2(n_273),
.B(n_285),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_275),
.C(n_282),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_215),
.C(n_152),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_304),
.C(n_312),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_291),
.B(n_183),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_301),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_318),
.A2(n_223),
.B1(n_183),
.B2(n_167),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_307),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_308),
.A2(n_288),
.B(n_290),
.Y(n_323)
);

AOI21xp33_ASAP7_75t_SL g337 ( 
.A1(n_323),
.A2(n_223),
.B(n_81),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_291),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_327),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_326),
.B(n_328),
.C(n_316),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_290),
.C(n_288),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_304),
.B(n_289),
.C(n_295),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_330),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_319),
.A2(n_317),
.B1(n_287),
.B2(n_308),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_326),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_331),
.B(n_335),
.Y(n_338)
);

OAI21xp33_ASAP7_75t_L g333 ( 
.A1(n_327),
.A2(n_314),
.B(n_303),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_333),
.A2(n_9),
.B(n_5),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_334),
.B(n_320),
.C(n_328),
.Y(n_342)
);

AND2x6_ASAP7_75t_L g336 ( 
.A(n_321),
.B(n_211),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_336),
.B(n_324),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_337),
.B(n_322),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_340),
.B(n_333),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_341),
.A2(n_343),
.B(n_336),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_342),
.B(n_334),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_344),
.B(n_345),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_339),
.B(n_332),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_346),
.A2(n_347),
.B(n_341),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_349),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_348),
.C(n_338),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_8),
.C(n_9),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_9),
.Y(n_353)
);


endmodule