module fake_jpeg_13366_n_206 (n_13, n_21, n_57, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_55, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_56, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_206);

input n_13;
input n_21;
input n_57;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_55;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_56;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_31),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_22),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_14),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_25),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_5),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_26),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

BUFx4f_ASAP7_75t_SL g75 ( 
.A(n_33),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_10),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_13),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_18),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_8),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_12),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_88),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_94),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_0),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_66),
.C(n_78),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_70),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_96),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_71),
.B1(n_86),
.B2(n_59),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_104),
.B1(n_69),
.B2(n_67),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_93),
.A2(n_78),
.B1(n_59),
.B2(n_80),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_100),
.A2(n_74),
.B1(n_65),
.B2(n_81),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_92),
.A2(n_86),
.B1(n_80),
.B2(n_66),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_101),
.A2(n_105),
.B1(n_110),
.B2(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_103),
.B(n_65),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_93),
.A2(n_85),
.B1(n_79),
.B2(n_83),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_58),
.B1(n_63),
.B2(n_77),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_111),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_88),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_84),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_132),
.B1(n_37),
.B2(n_45),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_117),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_115),
.A2(n_119),
.B1(n_128),
.B2(n_130),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_107),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_1),
.C(n_6),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_111),
.A2(n_76),
.B1(n_81),
.B2(n_72),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_109),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_123),
.Y(n_143)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_64),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_126),
.Y(n_153)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_94),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_129),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_98),
.A2(n_75),
.B1(n_96),
.B2(n_3),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_94),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_28),
.B1(n_55),
.B2(n_54),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_108),
.B(n_94),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_42),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_52),
.B1(n_51),
.B2(n_50),
.Y(n_132)
);

OA22x2_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_49),
.B1(n_48),
.B2(n_46),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_133),
.A2(n_126),
.B1(n_114),
.B2(n_116),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_0),
.Y(n_134)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_119),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_147),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_145),
.B1(n_146),
.B2(n_155),
.Y(n_158)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_133),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_141),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_142),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_127),
.A2(n_106),
.B1(n_3),
.B2(n_4),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_115),
.A2(n_106),
.B1(n_4),
.B2(n_5),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_128),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_7),
.Y(n_159)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_151),
.B(n_156),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_1),
.B1(n_6),
.B2(n_7),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_159),
.B(n_161),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_151),
.A2(n_141),
.B1(n_150),
.B2(n_154),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_8),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_169),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_40),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_170),
.C(n_13),
.Y(n_180)
);

A2O1A1O1Ixp25_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_39),
.B(n_38),
.C(n_36),
.D(n_34),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_166),
.A2(n_163),
.B(n_157),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_152),
.B(n_9),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_171),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_11),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_32),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_156),
.B(n_12),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_30),
.B1(n_29),
.B2(n_24),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_14),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_144),
.A2(n_139),
.B(n_148),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_140),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_179),
.B(n_180),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_137),
.Y(n_182)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_183),
.A2(n_172),
.B1(n_158),
.B2(n_167),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_137),
.Y(n_184)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_15),
.Y(n_185)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

OAI21xp33_ASAP7_75t_SL g186 ( 
.A1(n_162),
.A2(n_16),
.B(n_17),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_186),
.A2(n_162),
.B1(n_166),
.B2(n_158),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_188),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_181),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_190),
.A2(n_181),
.B1(n_186),
.B2(n_178),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_194),
.A2(n_196),
.B1(n_189),
.B2(n_188),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_198),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_180),
.C(n_193),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_195),
.B(n_187),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_193),
.B1(n_191),
.B2(n_177),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_175),
.B(n_173),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_202),
.A2(n_18),
.B(n_20),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_20),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_204),
.B(n_21),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_21),
.Y(n_206)
);


endmodule