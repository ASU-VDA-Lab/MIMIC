module fake_netlist_6_2378_n_108 (n_16, n_1, n_9, n_8, n_18, n_10, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_7, n_2, n_5, n_19, n_108);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_7;
input n_2;
input n_5;
input n_19;

output n_108;

wire n_52;
wire n_91;
wire n_46;
wire n_21;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_20;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_94;
wire n_97;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_40;
wire n_25;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVxp33_ASAP7_75t_SL g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVxp67_ASAP7_75t_SL g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVxp67_ASAP7_75t_SL g35 ( 
.A(n_12),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_2),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_20),
.B(n_4),
.Y(n_40)
);

AND2x4_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_13),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_7),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_23),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_28),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_20),
.B1(n_26),
.B2(n_35),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_30),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_46),
.B(n_39),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_50),
.Y(n_63)
);

AND2x4_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_53),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_53),
.B(n_55),
.Y(n_65)
);

CKINVDCx6p67_ASAP7_75t_R g66 ( 
.A(n_61),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_53),
.B1(n_50),
.B2(n_52),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_59),
.Y(n_70)
);

BUFx4f_ASAP7_75t_SL g71 ( 
.A(n_66),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_59),
.B(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_64),
.B(n_67),
.C(n_32),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_67),
.Y(n_76)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_74),
.A2(n_64),
.B(n_45),
.C(n_33),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_76),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_77),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_78),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_78),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_74),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_82),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_71),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_87),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_88),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_38),
.C(n_80),
.Y(n_96)
);

AOI221xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_33),
.B1(n_34),
.B2(n_48),
.C(n_47),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_93),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_85),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

OAI211xp5_ASAP7_75t_SL g101 ( 
.A1(n_97),
.A2(n_34),
.B(n_47),
.C(n_44),
.Y(n_101)
);

OAI211xp5_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_95),
.B(n_44),
.C(n_37),
.Y(n_102)
);

NOR2xp67_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_86),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_103),
.B1(n_99),
.B2(n_101),
.Y(n_104)
);

AOI211xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_86),
.B(n_56),
.C(n_73),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_71),
.B(n_19),
.C(n_17),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_72),
.B(n_105),
.Y(n_107)
);

AOI221xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_72),
.B1(n_106),
.B2(n_105),
.C(n_38),
.Y(n_108)
);


endmodule