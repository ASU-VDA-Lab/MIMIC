module real_aes_7105_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_404;
wire n_288;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI222xp33_ASAP7_75t_L g452 ( .A1(n_0), .A2(n_453), .B1(n_733), .B2(n_734), .C1(n_743), .C2(n_746), .Y(n_452) );
INVx1_ASAP7_75t_L g118 ( .A(n_1), .Y(n_118) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_2), .A2(n_140), .B(n_144), .C(n_239), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_3), .A2(n_176), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g465 ( .A(n_4), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_5), .B(n_216), .Y(n_273) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_6), .A2(n_735), .B1(n_736), .B2(n_742), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_6), .Y(n_742) );
AOI21xp33_ASAP7_75t_L g492 ( .A1(n_7), .A2(n_176), .B(n_493), .Y(n_492) );
AND2x6_ASAP7_75t_L g140 ( .A(n_8), .B(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g199 ( .A(n_9), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_10), .B(n_42), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_10), .B(n_42), .Y(n_752) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_11), .A2(n_175), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_12), .B(n_152), .Y(n_243) );
INVx1_ASAP7_75t_L g497 ( .A(n_13), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_14), .B(n_210), .Y(n_520) );
INVx1_ASAP7_75t_L g160 ( .A(n_15), .Y(n_160) );
INVx1_ASAP7_75t_L g541 ( .A(n_16), .Y(n_541) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_17), .A2(n_150), .B(n_224), .C(n_226), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_18), .B(n_216), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_19), .B(n_476), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_20), .B(n_176), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_21), .B(n_189), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_22), .A2(n_210), .B(n_211), .C(n_213), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_23), .B(n_216), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_24), .B(n_152), .Y(n_260) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_25), .A2(n_184), .B(n_226), .C(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_26), .B(n_152), .Y(n_151) );
CKINVDCx16_ASAP7_75t_R g256 ( .A(n_27), .Y(n_256) );
INVx1_ASAP7_75t_L g148 ( .A(n_28), .Y(n_148) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_29), .A2(n_737), .B1(n_738), .B2(n_739), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_29), .Y(n_737) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_30), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_31), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_32), .B(n_152), .Y(n_466) );
INVx1_ASAP7_75t_L g182 ( .A(n_33), .Y(n_182) );
INVx1_ASAP7_75t_L g487 ( .A(n_34), .Y(n_487) );
INVx2_ASAP7_75t_L g138 ( .A(n_35), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_36), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_37), .A2(n_210), .B(n_269), .C(n_271), .Y(n_268) );
INVxp67_ASAP7_75t_L g183 ( .A(n_38), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g143 ( .A1(n_39), .A2(n_144), .B(n_147), .C(n_155), .Y(n_143) );
CKINVDCx14_ASAP7_75t_R g267 ( .A(n_40), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_41), .A2(n_140), .B(n_144), .C(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g486 ( .A(n_43), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_44), .A2(n_197), .B(n_198), .C(n_200), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_45), .B(n_152), .Y(n_531) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_46), .A2(n_50), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_46), .Y(n_127) );
AOI22xp5_ASAP7_75t_SL g104 ( .A1(n_47), .A2(n_105), .B1(n_750), .B2(n_751), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_48), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_49), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_50), .Y(n_126) );
INVx1_ASAP7_75t_L g208 ( .A(n_51), .Y(n_208) );
CKINVDCx16_ASAP7_75t_R g488 ( .A(n_52), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_53), .B(n_176), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_54), .A2(n_144), .B1(n_213), .B2(n_485), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_55), .Y(n_514) );
CKINVDCx16_ASAP7_75t_R g462 ( .A(n_56), .Y(n_462) );
CKINVDCx14_ASAP7_75t_R g195 ( .A(n_57), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_58), .A2(n_197), .B(n_271), .C(n_496), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_59), .Y(n_534) );
INVx1_ASAP7_75t_L g494 ( .A(n_60), .Y(n_494) );
INVx1_ASAP7_75t_L g141 ( .A(n_61), .Y(n_141) );
INVx1_ASAP7_75t_L g159 ( .A(n_62), .Y(n_159) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_63), .A2(n_92), .B1(n_740), .B2(n_741), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_63), .Y(n_740) );
INVx1_ASAP7_75t_SL g270 ( .A(n_64), .Y(n_270) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_65), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_66), .B(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g259 ( .A(n_67), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_SL g475 ( .A1(n_68), .A2(n_271), .B(n_476), .C(n_477), .Y(n_475) );
INVxp67_ASAP7_75t_L g478 ( .A(n_69), .Y(n_478) );
INVx1_ASAP7_75t_L g756 ( .A(n_70), .Y(n_756) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_71), .A2(n_176), .B(n_194), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_72), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_73), .A2(n_176), .B(n_221), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_74), .Y(n_490) );
INVx1_ASAP7_75t_L g528 ( .A(n_75), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_76), .A2(n_175), .B(n_177), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g142 ( .A(n_77), .Y(n_142) );
INVx1_ASAP7_75t_L g222 ( .A(n_78), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_79), .A2(n_140), .B(n_144), .C(n_530), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_80), .A2(n_176), .B(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g225 ( .A(n_81), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_82), .B(n_149), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_83), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g157 ( .A(n_84), .Y(n_157) );
INVx1_ASAP7_75t_L g240 ( .A(n_85), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_86), .B(n_476), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g463 ( .A1(n_87), .A2(n_140), .B(n_144), .C(n_464), .Y(n_463) );
OR2x2_ASAP7_75t_L g115 ( .A(n_88), .B(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g729 ( .A(n_88), .Y(n_729) );
OR2x2_ASAP7_75t_L g732 ( .A(n_88), .B(n_117), .Y(n_732) );
NAND3xp33_ASAP7_75t_SL g753 ( .A(n_88), .B(n_118), .C(n_754), .Y(n_753) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_89), .A2(n_144), .B(n_258), .C(n_261), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_90), .B(n_156), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_91), .Y(n_469) );
CKINVDCx14_ASAP7_75t_R g741 ( .A(n_92), .Y(n_741) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_93), .A2(n_103), .B1(n_122), .B2(n_123), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_93), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_94), .A2(n_140), .B(n_144), .C(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g474 ( .A(n_95), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g538 ( .A(n_96), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_97), .B(n_149), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_98), .B(n_164), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_99), .B(n_164), .Y(n_542) );
INVx2_ASAP7_75t_L g212 ( .A(n_100), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_101), .A2(n_176), .B(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_102), .B(n_756), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_103), .Y(n_123) );
OA21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_111), .B(n_451), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
BUFx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g749 ( .A(n_110), .Y(n_749) );
OAI21xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_120), .B(n_448), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_115), .Y(n_450) );
NOR2x2_ASAP7_75t_L g745 ( .A(n_116), .B(n_729), .Y(n_745) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OR2x2_ASAP7_75t_L g728 ( .A(n_117), .B(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
AOI22xp33_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_124), .B1(n_446), .B2(n_447), .Y(n_120) );
INVx1_ASAP7_75t_L g446 ( .A(n_121), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_122), .B(n_235), .Y(n_523) );
INVx1_ASAP7_75t_L g447 ( .A(n_124), .Y(n_447) );
XNOR2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_128), .Y(n_124) );
OAI22xp5_ASAP7_75t_SL g453 ( .A1(n_128), .A2(n_454), .B1(n_726), .B2(n_730), .Y(n_453) );
INVx1_ASAP7_75t_SL g748 ( .A(n_128), .Y(n_748) );
OR5x1_ASAP7_75t_L g128 ( .A(n_129), .B(n_340), .C(n_404), .D(n_420), .E(n_435), .Y(n_128) );
NAND4xp25_ASAP7_75t_L g129 ( .A(n_130), .B(n_274), .C(n_301), .D(n_324), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_217), .B(n_228), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_166), .Y(n_131) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx3_ASAP7_75t_SL g251 ( .A(n_133), .Y(n_251) );
AND2x4_ASAP7_75t_L g287 ( .A(n_133), .B(n_276), .Y(n_287) );
OR2x2_ASAP7_75t_L g297 ( .A(n_133), .B(n_253), .Y(n_297) );
OR2x2_ASAP7_75t_L g343 ( .A(n_133), .B(n_169), .Y(n_343) );
AND2x2_ASAP7_75t_L g357 ( .A(n_133), .B(n_252), .Y(n_357) );
AND2x2_ASAP7_75t_L g400 ( .A(n_133), .B(n_290), .Y(n_400) );
AND2x2_ASAP7_75t_L g407 ( .A(n_133), .B(n_264), .Y(n_407) );
AND2x2_ASAP7_75t_L g426 ( .A(n_133), .B(n_316), .Y(n_426) );
AND2x2_ASAP7_75t_L g444 ( .A(n_133), .B(n_286), .Y(n_444) );
OR2x6_ASAP7_75t_L g133 ( .A(n_134), .B(n_161), .Y(n_133) );
O2A1O1Ixp33_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_142), .B(n_143), .C(n_156), .Y(n_134) );
OAI21xp5_ASAP7_75t_L g236 ( .A1(n_135), .A2(n_237), .B(n_238), .Y(n_236) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_135), .A2(n_256), .B(n_257), .Y(n_255) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_135), .A2(n_462), .B(n_463), .Y(n_461) );
OAI22xp33_ASAP7_75t_L g483 ( .A1(n_135), .A2(n_186), .B1(n_484), .B2(n_488), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g527 ( .A1(n_135), .A2(n_528), .B(n_529), .Y(n_527) );
NAND2x1p5_ASAP7_75t_L g135 ( .A(n_136), .B(n_140), .Y(n_135) );
AND2x4_ASAP7_75t_L g176 ( .A(n_136), .B(n_140), .Y(n_176) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx1_ASAP7_75t_L g154 ( .A(n_137), .Y(n_154) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g145 ( .A(n_138), .Y(n_145) );
INVx1_ASAP7_75t_L g214 ( .A(n_138), .Y(n_214) );
INVx1_ASAP7_75t_L g146 ( .A(n_139), .Y(n_146) );
INVx3_ASAP7_75t_L g150 ( .A(n_139), .Y(n_150) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_139), .Y(n_152) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_139), .Y(n_185) );
INVx1_ASAP7_75t_L g476 ( .A(n_139), .Y(n_476) );
BUFx3_ASAP7_75t_L g155 ( .A(n_140), .Y(n_155) );
INVx4_ASAP7_75t_SL g186 ( .A(n_140), .Y(n_186) );
INVx5_ASAP7_75t_L g179 ( .A(n_144), .Y(n_179) );
AND2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
BUFx3_ASAP7_75t_L g201 ( .A(n_145), .Y(n_201) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_145), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B(n_151), .C(n_153), .Y(n_147) );
OAI22xp33_ASAP7_75t_L g181 ( .A1(n_149), .A2(n_182), .B1(n_183), .B2(n_184), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_L g464 ( .A1(n_149), .A2(n_465), .B(n_466), .C(n_467), .Y(n_464) );
INVx5_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_150), .B(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_150), .B(n_478), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_150), .B(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g197 ( .A(n_152), .Y(n_197) );
INVx4_ASAP7_75t_L g210 ( .A(n_152), .Y(n_210) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_154), .B(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g190 ( .A(n_156), .Y(n_190) );
OA21x2_ASAP7_75t_L g192 ( .A1(n_156), .A2(n_193), .B(n_202), .Y(n_192) );
INVx1_ASAP7_75t_L g235 ( .A(n_156), .Y(n_235) );
OA21x2_ASAP7_75t_L g535 ( .A1(n_156), .A2(n_536), .B(n_542), .Y(n_535) );
AND2x2_ASAP7_75t_SL g156 ( .A(n_157), .B(n_158), .Y(n_156) );
AND2x2_ASAP7_75t_L g165 ( .A(n_157), .B(n_158), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
INVx3_ASAP7_75t_L g216 ( .A(n_163), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_163), .B(n_246), .Y(n_245) );
AO21x2_ASAP7_75t_L g254 ( .A1(n_163), .A2(n_255), .B(n_262), .Y(n_254) );
NOR2xp33_ASAP7_75t_SL g513 ( .A(n_163), .B(n_514), .Y(n_513) );
INVx4_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_164), .Y(n_205) );
OA21x2_ASAP7_75t_L g471 ( .A1(n_164), .A2(n_472), .B(n_479), .Y(n_471) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g172 ( .A(n_165), .Y(n_172) );
INVx1_ASAP7_75t_L g409 ( .A(n_166), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_167), .B(n_191), .Y(n_166) );
AND2x2_ASAP7_75t_L g319 ( .A(n_167), .B(n_252), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_167), .B(n_339), .Y(n_338) );
AOI32xp33_ASAP7_75t_L g352 ( .A1(n_167), .A2(n_353), .A3(n_356), .B1(n_358), .B2(n_362), .Y(n_352) );
AND2x2_ASAP7_75t_L g422 ( .A(n_167), .B(n_316), .Y(n_422) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_SL g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g286 ( .A(n_169), .B(n_253), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_169), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g328 ( .A(n_169), .B(n_275), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_169), .B(n_407), .Y(n_406) );
AO21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_173), .B(n_187), .Y(n_169) );
INVx1_ASAP7_75t_L g291 ( .A(n_170), .Y(n_291) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_170), .A2(n_527), .B(n_533), .Y(n_526) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AOI21xp5_ASAP7_75t_SL g507 ( .A1(n_171), .A2(n_508), .B(n_509), .Y(n_507) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AO21x2_ASAP7_75t_L g460 ( .A1(n_172), .A2(n_461), .B(n_468), .Y(n_460) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_172), .A2(n_483), .B(n_489), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_172), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
OA21x2_ASAP7_75t_L g290 ( .A1(n_174), .A2(n_188), .B(n_291), .Y(n_290) );
BUFx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_SL g177 ( .A1(n_178), .A2(n_179), .B(n_180), .C(n_186), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_SL g194 ( .A1(n_179), .A2(n_186), .B(n_195), .C(n_196), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_SL g207 ( .A1(n_179), .A2(n_186), .B(n_208), .C(n_209), .Y(n_207) );
O2A1O1Ixp33_ASAP7_75t_SL g221 ( .A1(n_179), .A2(n_186), .B(n_222), .C(n_223), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g266 ( .A1(n_179), .A2(n_186), .B(n_267), .C(n_268), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_179), .A2(n_186), .B(n_474), .C(n_475), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_179), .A2(n_186), .B(n_494), .C(n_495), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_L g537 ( .A1(n_179), .A2(n_186), .B(n_538), .C(n_539), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_184), .B(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_184), .B(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_184), .B(n_541), .Y(n_540) );
INVx4_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g242 ( .A(n_185), .Y(n_242) );
OAI22xp5_ASAP7_75t_SL g485 ( .A1(n_185), .A2(n_242), .B1(n_486), .B2(n_487), .Y(n_485) );
INVx1_ASAP7_75t_L g261 ( .A(n_186), .Y(n_261) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_190), .B(n_263), .Y(n_262) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_190), .A2(n_516), .B(n_523), .Y(n_515) );
AND2x2_ASAP7_75t_L g293 ( .A(n_191), .B(n_232), .Y(n_293) );
AND2x2_ASAP7_75t_L g369 ( .A(n_191), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_SL g441 ( .A(n_191), .Y(n_441) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_203), .Y(n_191) );
OR2x2_ASAP7_75t_L g231 ( .A(n_192), .B(n_204), .Y(n_231) );
AND2x2_ASAP7_75t_L g248 ( .A(n_192), .B(n_249), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_192), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g300 ( .A(n_192), .Y(n_300) );
AND2x2_ASAP7_75t_L g327 ( .A(n_192), .B(n_204), .Y(n_327) );
BUFx3_ASAP7_75t_L g330 ( .A(n_192), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_192), .B(n_305), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_192), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g244 ( .A(n_200), .Y(n_244) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g226 ( .A(n_201), .Y(n_226) );
INVx2_ASAP7_75t_L g281 ( .A(n_203), .Y(n_281) );
AND2x2_ASAP7_75t_L g299 ( .A(n_203), .B(n_279), .Y(n_299) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g310 ( .A(n_204), .B(n_219), .Y(n_310) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_204), .Y(n_323) );
OA21x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_215), .Y(n_204) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_205), .A2(n_220), .B(n_227), .Y(n_219) );
OA21x2_ASAP7_75t_L g264 ( .A1(n_205), .A2(n_265), .B(n_273), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_210), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g467 ( .A(n_213), .Y(n_467) );
INVx3_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_216), .A2(n_492), .B(n_498), .Y(n_491) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_218), .B(n_330), .Y(n_380) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_SL g249 ( .A(n_219), .Y(n_249) );
NAND3xp33_ASAP7_75t_L g298 ( .A(n_219), .B(n_299), .C(n_300), .Y(n_298) );
OR2x2_ASAP7_75t_L g306 ( .A(n_219), .B(n_279), .Y(n_306) );
AND2x2_ASAP7_75t_L g326 ( .A(n_219), .B(n_279), .Y(n_326) );
AND2x2_ASAP7_75t_L g370 ( .A(n_219), .B(n_234), .Y(n_370) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_247), .B(n_250), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_230), .B(n_232), .Y(n_229) );
AND2x2_ASAP7_75t_L g445 ( .A(n_230), .B(n_370), .Y(n_445) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_231), .A2(n_343), .B1(n_385), .B2(n_387), .Y(n_384) );
OR2x2_ASAP7_75t_L g391 ( .A(n_231), .B(n_306), .Y(n_391) );
OR2x2_ASAP7_75t_L g415 ( .A(n_231), .B(n_416), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_231), .B(n_335), .Y(n_428) );
AND2x2_ASAP7_75t_L g321 ( .A(n_232), .B(n_322), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_232), .A2(n_394), .B(n_409), .Y(n_408) );
AOI32xp33_ASAP7_75t_L g429 ( .A1(n_232), .A2(n_319), .A3(n_430), .B1(n_432), .B2(n_433), .Y(n_429) );
OR2x2_ASAP7_75t_L g440 ( .A(n_232), .B(n_441), .Y(n_440) );
CKINVDCx16_ASAP7_75t_R g232 ( .A(n_233), .Y(n_232) );
OR2x2_ASAP7_75t_L g308 ( .A(n_233), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_233), .B(n_322), .Y(n_387) );
BUFx3_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx4_ASAP7_75t_L g279 ( .A(n_234), .Y(n_279) );
AND2x2_ASAP7_75t_L g345 ( .A(n_234), .B(n_310), .Y(n_345) );
AND3x2_ASAP7_75t_L g354 ( .A(n_234), .B(n_248), .C(n_355), .Y(n_354) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_245), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_235), .B(n_469), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_235), .B(n_534), .Y(n_533) );
O2A1O1Ixp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_243), .C(n_244), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g258 ( .A1(n_241), .A2(n_244), .B(n_259), .C(n_260), .Y(n_258) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_244), .A2(n_511), .B(n_512), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_244), .A2(n_531), .B(n_532), .Y(n_530) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g280 ( .A(n_249), .B(n_281), .Y(n_280) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_249), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_249), .B(n_279), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
AND2x2_ASAP7_75t_L g275 ( .A(n_251), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g315 ( .A(n_251), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g333 ( .A(n_251), .B(n_264), .Y(n_333) );
AND2x2_ASAP7_75t_L g351 ( .A(n_251), .B(n_253), .Y(n_351) );
OR2x2_ASAP7_75t_L g365 ( .A(n_251), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g411 ( .A(n_251), .B(n_339), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_252), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_264), .Y(n_252) );
AND2x2_ASAP7_75t_L g312 ( .A(n_253), .B(n_290), .Y(n_312) );
OR2x2_ASAP7_75t_L g366 ( .A(n_253), .B(n_290), .Y(n_366) );
AND2x2_ASAP7_75t_L g419 ( .A(n_253), .B(n_276), .Y(n_419) );
INVx2_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
BUFx2_ASAP7_75t_L g317 ( .A(n_254), .Y(n_317) );
AND2x2_ASAP7_75t_L g339 ( .A(n_254), .B(n_264), .Y(n_339) );
INVx2_ASAP7_75t_L g276 ( .A(n_264), .Y(n_276) );
INVx1_ASAP7_75t_L g296 ( .A(n_264), .Y(n_296) );
INVx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_272), .Y(n_521) );
AOI211xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_277), .B(n_282), .C(n_294), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_275), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g438 ( .A(n_275), .Y(n_438) );
AND2x2_ASAP7_75t_L g316 ( .A(n_276), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_279), .B(n_280), .Y(n_288) );
INVx1_ASAP7_75t_L g373 ( .A(n_279), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_279), .B(n_300), .Y(n_397) );
AND2x2_ASAP7_75t_L g413 ( .A(n_279), .B(n_327), .Y(n_413) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_280), .B(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g304 ( .A(n_281), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_288), .B1(n_289), .B2(n_292), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_285), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_286), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g311 ( .A(n_287), .B(n_312), .Y(n_311) );
AOI221xp5_ASAP7_75t_SL g376 ( .A1(n_287), .A2(n_329), .B1(n_377), .B2(n_382), .C(n_384), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_287), .B(n_350), .Y(n_383) );
INVx1_ASAP7_75t_L g443 ( .A(n_289), .Y(n_443) );
BUFx3_ASAP7_75t_L g350 ( .A(n_290), .Y(n_350) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI21xp33_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_297), .B(n_298), .Y(n_294) );
INVx1_ASAP7_75t_L g359 ( .A(n_296), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_296), .B(n_350), .Y(n_403) );
INVx1_ASAP7_75t_L g360 ( .A(n_297), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g361 ( .A(n_297), .B(n_350), .Y(n_361) );
INVxp67_ASAP7_75t_L g381 ( .A(n_299), .Y(n_381) );
AND2x2_ASAP7_75t_L g322 ( .A(n_300), .B(n_323), .Y(n_322) );
O2A1O1Ixp33_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_307), .B(n_311), .C(n_313), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_SL g336 ( .A(n_304), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_305), .B(n_336), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_305), .B(n_327), .Y(n_378) );
INVx2_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_308), .A2(n_314), .B1(n_318), .B2(n_320), .Y(n_313) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g329 ( .A(n_310), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g374 ( .A(n_310), .B(n_375), .Y(n_374) );
OAI21xp33_ASAP7_75t_L g377 ( .A1(n_312), .A2(n_378), .B(n_379), .Y(n_377) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
AOI221xp5_ASAP7_75t_L g324 ( .A1(n_316), .A2(n_325), .B1(n_328), .B2(n_329), .C(n_331), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_316), .B(n_350), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_316), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g432 ( .A(n_322), .Y(n_432) );
INVxp67_ASAP7_75t_L g355 ( .A(n_323), .Y(n_355) );
INVx1_ASAP7_75t_L g362 ( .A(n_325), .Y(n_362) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
AND2x2_ASAP7_75t_L g401 ( .A(n_326), .B(n_330), .Y(n_401) );
INVx1_ASAP7_75t_L g375 ( .A(n_330), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_330), .B(n_345), .Y(n_405) );
OAI32xp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_334), .A3(n_336), .B1(n_337), .B2(n_338), .Y(n_331) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx2_ASAP7_75t_SL g344 ( .A(n_339), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_339), .B(n_371), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_339), .B(n_400), .Y(n_431) );
NAND2x1p5_ASAP7_75t_L g439 ( .A(n_339), .B(n_350), .Y(n_439) );
NAND5xp2_ASAP7_75t_L g340 ( .A(n_341), .B(n_363), .C(n_376), .D(n_388), .E(n_389), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_345), .B1(n_346), .B2(n_348), .C(n_352), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp33_ASAP7_75t_SL g367 ( .A(n_347), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_350), .B(n_419), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_351), .A2(n_364), .B1(n_367), .B2(n_371), .Y(n_363) );
INVx2_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
OAI211xp5_ASAP7_75t_SL g358 ( .A1(n_354), .A2(n_359), .B(n_360), .C(n_361), .Y(n_358) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_SL g386 ( .A(n_366), .Y(n_386) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_375), .B(n_424), .Y(n_434) );
OR2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AOI222xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_392), .B1(n_394), .B2(n_398), .C1(n_401), .C2(n_402), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OAI221xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B1(n_408), .B2(n_410), .C(n_412), .Y(n_404) );
INVx1_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
OAI21xp33_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_414), .B(n_417), .Y(n_412) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g424 ( .A(n_416), .Y(n_424) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI221xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_423), .B1(n_425), .B2(n_427), .C(n_429), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
A2O1A1Ixp33_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_439), .B(n_440), .C(n_442), .Y(n_435) );
INVxp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI21xp33_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B(n_445), .Y(n_442) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_448), .B(n_452), .C(n_749), .Y(n_451) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g747 ( .A(n_454), .Y(n_747) );
OR4x1_ASAP7_75t_L g454 ( .A(n_455), .B(n_615), .C(n_675), .D(n_702), .Y(n_454) );
NAND4xp25_ASAP7_75t_SL g455 ( .A(n_456), .B(n_563), .C(n_594), .D(n_611), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_499), .B(n_501), .C(n_543), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_480), .Y(n_457) );
INVx1_ASAP7_75t_L g605 ( .A(n_458), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_458), .A2(n_646), .B1(n_694), .B2(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_470), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_459), .B(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g556 ( .A(n_459), .B(n_482), .Y(n_556) );
AND2x2_ASAP7_75t_L g598 ( .A(n_459), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_459), .B(n_500), .Y(n_610) );
INVx1_ASAP7_75t_L g650 ( .A(n_459), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_459), .B(n_704), .Y(n_703) );
INVx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g578 ( .A(n_460), .B(n_482), .Y(n_578) );
INVx3_ASAP7_75t_L g582 ( .A(n_460), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_460), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g669 ( .A(n_470), .B(n_491), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_470), .B(n_582), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_470), .B(n_697), .Y(n_696) );
INVx3_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g500 ( .A(n_471), .B(n_482), .Y(n_500) );
INVx1_ASAP7_75t_L g551 ( .A(n_471), .Y(n_551) );
BUFx2_ASAP7_75t_L g555 ( .A(n_471), .Y(n_555) );
AND2x2_ASAP7_75t_L g599 ( .A(n_471), .B(n_481), .Y(n_599) );
OR2x2_ASAP7_75t_L g638 ( .A(n_471), .B(n_481), .Y(n_638) );
AND2x2_ASAP7_75t_L g663 ( .A(n_471), .B(n_491), .Y(n_663) );
AND2x2_ASAP7_75t_L g722 ( .A(n_471), .B(n_552), .Y(n_722) );
INVx1_ASAP7_75t_L g697 ( .A(n_480), .Y(n_697) );
OR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_491), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_481), .B(n_491), .Y(n_583) );
AND2x2_ASAP7_75t_L g593 ( .A(n_481), .B(n_582), .Y(n_593) );
BUFx2_ASAP7_75t_L g604 ( .A(n_481), .Y(n_604) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g626 ( .A(n_482), .B(n_491), .Y(n_626) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_482), .Y(n_681) );
AND2x2_ASAP7_75t_SL g499 ( .A(n_491), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_SL g552 ( .A(n_491), .Y(n_552) );
BUFx2_ASAP7_75t_L g577 ( .A(n_491), .Y(n_577) );
INVx2_ASAP7_75t_L g596 ( .A(n_491), .Y(n_596) );
AND2x2_ASAP7_75t_L g658 ( .A(n_491), .B(n_582), .Y(n_658) );
AOI321xp33_ASAP7_75t_L g677 ( .A1(n_499), .A2(n_678), .A3(n_679), .B1(n_680), .B2(n_682), .C(n_683), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_500), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_500), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g671 ( .A(n_500), .B(n_650), .Y(n_671) );
AND2x2_ASAP7_75t_L g704 ( .A(n_500), .B(n_596), .Y(n_704) );
INVx1_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_524), .Y(n_502) );
OR2x2_ASAP7_75t_L g606 ( .A(n_503), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_515), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx3_ASAP7_75t_L g558 ( .A(n_506), .Y(n_558) );
AND2x2_ASAP7_75t_L g568 ( .A(n_506), .B(n_526), .Y(n_568) );
AND2x2_ASAP7_75t_L g573 ( .A(n_506), .B(n_548), .Y(n_573) );
INVx1_ASAP7_75t_L g590 ( .A(n_506), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_506), .B(n_571), .Y(n_609) );
AND2x2_ASAP7_75t_L g614 ( .A(n_506), .B(n_547), .Y(n_614) );
OR2x2_ASAP7_75t_L g646 ( .A(n_506), .B(n_635), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_506), .B(n_559), .Y(n_685) );
AND2x2_ASAP7_75t_L g719 ( .A(n_506), .B(n_545), .Y(n_719) );
OR2x6_ASAP7_75t_L g506 ( .A(n_507), .B(n_513), .Y(n_506) );
INVx1_ASAP7_75t_L g546 ( .A(n_515), .Y(n_546) );
INVx2_ASAP7_75t_L g561 ( .A(n_515), .Y(n_561) );
AND2x2_ASAP7_75t_L g601 ( .A(n_515), .B(n_572), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_515), .B(n_548), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_522), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B(n_521), .Y(n_518) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g707 ( .A(n_525), .B(n_558), .Y(n_707) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_535), .Y(n_525) );
INVx2_ASAP7_75t_L g548 ( .A(n_526), .Y(n_548) );
AND2x2_ASAP7_75t_L g701 ( .A(n_526), .B(n_561), .Y(n_701) );
AND2x2_ASAP7_75t_L g547 ( .A(n_535), .B(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g562 ( .A(n_535), .Y(n_562) );
INVx1_ASAP7_75t_L g572 ( .A(n_535), .Y(n_572) );
OAI22xp33_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_549), .B1(n_553), .B2(n_557), .Y(n_543) );
OAI22xp33_ASAP7_75t_L g698 ( .A1(n_544), .A2(n_662), .B1(n_699), .B2(n_700), .Y(n_698) );
INVx1_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
INVx1_ASAP7_75t_L g613 ( .A(n_546), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_547), .B(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g608 ( .A(n_548), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_548), .B(n_561), .Y(n_635) );
INVx1_ASAP7_75t_L g651 ( .A(n_548), .Y(n_651) );
AND2x2_ASAP7_75t_L g592 ( .A(n_550), .B(n_593), .Y(n_592) );
INVx3_ASAP7_75t_SL g631 ( .A(n_550), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_550), .B(n_556), .Y(n_708) );
AND2x4_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
INVx1_ASAP7_75t_L g717 ( .A(n_553), .Y(n_717) );
OR2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_554), .B(n_650), .Y(n_692) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx3_ASAP7_75t_SL g597 ( .A(n_556), .Y(n_597) );
NAND2x1_ASAP7_75t_SL g557 ( .A(n_558), .B(n_559), .Y(n_557) );
AND2x2_ASAP7_75t_L g618 ( .A(n_558), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g625 ( .A(n_558), .B(n_562), .Y(n_625) );
AND2x2_ASAP7_75t_L g630 ( .A(n_558), .B(n_571), .Y(n_630) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_558), .Y(n_679) );
OAI311xp33_ASAP7_75t_L g702 ( .A1(n_559), .A2(n_703), .A3(n_705), .B1(n_706), .C1(n_716), .Y(n_702) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OR2x2_ASAP7_75t_L g715 ( .A(n_560), .B(n_588), .Y(n_715) );
OR2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
AND2x2_ASAP7_75t_L g571 ( .A(n_561), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g619 ( .A(n_561), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g674 ( .A(n_561), .Y(n_674) );
INVx1_ASAP7_75t_L g567 ( .A(n_562), .Y(n_567) );
INVx1_ASAP7_75t_L g587 ( .A(n_562), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_562), .B(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g620 ( .A(n_562), .Y(n_620) );
AOI221xp5_ASAP7_75t_SL g563 ( .A1(n_564), .A2(n_566), .B1(n_574), .B2(n_579), .C(n_584), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_569), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx4_ASAP7_75t_L g588 ( .A(n_568), .Y(n_588) );
AND2x2_ASAP7_75t_L g682 ( .A(n_568), .B(n_601), .Y(n_682) );
AND2x2_ASAP7_75t_L g689 ( .A(n_568), .B(n_571), .Y(n_689) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_571), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g600 ( .A(n_573), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_578), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_576), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g725 ( .A(n_578), .B(n_669), .Y(n_725) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g710 ( .A(n_582), .B(n_638), .Y(n_710) );
OAI211xp5_ASAP7_75t_L g675 ( .A1(n_583), .A2(n_676), .B(n_677), .C(n_690), .Y(n_675) );
AOI21xp33_ASAP7_75t_SL g584 ( .A1(n_585), .A2(n_589), .B(n_591), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NOR2xp67_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g654 ( .A(n_588), .Y(n_654) );
OAI221xp5_ASAP7_75t_L g683 ( .A1(n_589), .A2(n_684), .B1(n_685), .B2(n_686), .C(n_687), .Y(n_683) );
AND2x2_ASAP7_75t_L g660 ( .A(n_590), .B(n_601), .Y(n_660) );
AND2x2_ASAP7_75t_L g713 ( .A(n_590), .B(n_608), .Y(n_713) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_593), .B(n_631), .Y(n_655) );
O2A1O1Ixp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_598), .B(n_600), .C(n_602), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
AND2x2_ASAP7_75t_L g641 ( .A(n_596), .B(n_599), .Y(n_641) );
OR2x2_ASAP7_75t_L g684 ( .A(n_596), .B(n_638), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_597), .B(n_663), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_597), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_SL g628 ( .A(n_598), .Y(n_628) );
INVx1_ASAP7_75t_L g694 ( .A(n_601), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_606), .B1(n_609), .B2(n_610), .Y(n_602) );
INVx1_ASAP7_75t_L g617 ( .A(n_603), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_604), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g680 ( .A(n_605), .B(n_681), .Y(n_680) );
INVxp67_ASAP7_75t_L g666 ( .A(n_607), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_608), .B(n_694), .Y(n_693) );
OAI22xp33_ASAP7_75t_L g667 ( .A1(n_609), .A2(n_668), .B1(n_670), .B2(n_672), .Y(n_667) );
INVx1_ASAP7_75t_L g676 ( .A(n_612), .Y(n_676) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
AND2x2_ASAP7_75t_L g718 ( .A(n_613), .B(n_713), .Y(n_718) );
AOI222xp33_ASAP7_75t_L g647 ( .A1(n_614), .A2(n_648), .B1(n_651), .B2(n_652), .C1(n_655), .C2(n_656), .Y(n_647) );
NAND4xp25_ASAP7_75t_SL g615 ( .A(n_616), .B(n_636), .C(n_647), .D(n_659), .Y(n_615) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B1(n_621), .B2(n_626), .C(n_627), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_619), .B(n_654), .Y(n_653) );
INVxp67_ASAP7_75t_L g645 ( .A(n_620), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_621), .A2(n_691), .B1(n_693), .B2(n_695), .C(n_698), .Y(n_690) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g633 ( .A(n_625), .B(n_634), .Y(n_633) );
OAI21xp33_ASAP7_75t_L g687 ( .A1(n_626), .A2(n_688), .B(n_689), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .B1(n_631), .B2(n_632), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI21xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_639), .B(n_642), .Y(n_636) );
INVxp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g678 ( .A(n_649), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_650), .B(n_669), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_650), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_654), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_SL g686 ( .A(n_658), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_661), .B1(n_664), .B2(n_666), .C(n_667), .Y(n_659) );
INVxp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AOI222xp33_ASAP7_75t_L g706 ( .A1(n_669), .A2(n_707), .B1(n_708), .B2(n_709), .C1(n_711), .C2(n_714), .Y(n_706) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_673), .B(n_713), .Y(n_712) );
INVxp67_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g705 ( .A(n_679), .Y(n_705) );
INVxp67_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVxp33_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AOI221xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B1(n_719), .B2(n_720), .C(n_723), .Y(n_716) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVxp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
OAI22xp5_ASAP7_75t_SL g746 ( .A1(n_726), .A2(n_732), .B1(n_747), .B2(n_748), .Y(n_746) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
CKINVDCx16_ASAP7_75t_R g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
INVx3_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
OR2x2_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
endmodule