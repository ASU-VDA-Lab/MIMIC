module real_aes_7657_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_755;
wire n_153;
wire n_316;
wire n_532;
wire n_284;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_0), .B(n_109), .C(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g447 ( .A(n_0), .Y(n_447) );
INVx1_ASAP7_75t_L g537 ( .A(n_1), .Y(n_537) );
INVx1_ASAP7_75t_L g199 ( .A(n_2), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_3), .A2(n_40), .B1(n_161), .B2(n_479), .Y(n_496) );
AOI21xp33_ASAP7_75t_L g140 ( .A1(n_4), .A2(n_141), .B(n_148), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_5), .B(n_134), .Y(n_528) );
AND2x6_ASAP7_75t_L g146 ( .A(n_6), .B(n_147), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_7), .A2(n_240), .B(n_241), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_8), .B(n_107), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_8), .B(n_42), .Y(n_448) );
INVx1_ASAP7_75t_L g158 ( .A(n_9), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_10), .B(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g139 ( .A(n_11), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_12), .B(n_171), .Y(n_474) );
INVx1_ASAP7_75t_L g246 ( .A(n_13), .Y(n_246) );
INVx1_ASAP7_75t_L g532 ( .A(n_14), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_15), .B(n_135), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_16), .A2(n_748), .B1(n_749), .B2(n_752), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_16), .Y(n_752) );
AO32x2_ASAP7_75t_L g494 ( .A1(n_17), .A2(n_134), .A3(n_168), .B1(n_495), .B2(n_499), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_18), .B(n_161), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_19), .B(n_187), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_20), .B(n_135), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_21), .A2(n_53), .B1(n_161), .B2(n_479), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_22), .B(n_141), .Y(n_211) );
AOI22xp33_ASAP7_75t_SL g507 ( .A1(n_23), .A2(n_79), .B1(n_161), .B2(n_171), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_24), .B(n_161), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_25), .B(n_132), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_26), .A2(n_244), .B(n_245), .C(n_247), .Y(n_243) );
OAI22xp5_ASAP7_75t_SL g749 ( .A1(n_27), .A2(n_77), .B1(n_750), .B2(n_751), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_27), .Y(n_751) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_28), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_29), .B(n_164), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_30), .B(n_156), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_31), .A2(n_104), .B1(n_113), .B2(n_761), .Y(n_103) );
INVx1_ASAP7_75t_L g177 ( .A(n_32), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_33), .B(n_164), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_34), .B(n_443), .Y(n_452) );
INVx2_ASAP7_75t_L g144 ( .A(n_35), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_36), .B(n_161), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_37), .B(n_164), .Y(n_480) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_38), .A2(n_65), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_38), .Y(n_123) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_39), .A2(n_146), .B(n_151), .C(n_213), .Y(n_212) );
AOI222xp33_ASAP7_75t_L g454 ( .A1(n_41), .A2(n_455), .B1(n_746), .B2(n_747), .C1(n_753), .C2(n_757), .Y(n_454) );
INVx1_ASAP7_75t_L g107 ( .A(n_42), .Y(n_107) );
INVx1_ASAP7_75t_L g175 ( .A(n_43), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_44), .B(n_156), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_45), .B(n_161), .Y(n_522) );
OAI321xp33_ASAP7_75t_L g119 ( .A1(n_46), .A2(n_120), .A3(n_443), .B1(n_449), .B2(n_450), .C(n_452), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g449 ( .A(n_46), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_47), .A2(n_89), .B1(n_218), .B2(n_479), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_48), .B(n_161), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_49), .B(n_161), .Y(n_533) );
CKINVDCx16_ASAP7_75t_R g178 ( .A(n_50), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_51), .B(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_52), .B(n_141), .Y(n_234) );
AOI22xp33_ASAP7_75t_SL g517 ( .A1(n_54), .A2(n_63), .B1(n_161), .B2(n_171), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_55), .A2(n_151), .B1(n_171), .B2(n_173), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_56), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_57), .B(n_161), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g196 ( .A(n_58), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_59), .B(n_161), .Y(n_550) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_60), .A2(n_155), .B(n_157), .C(n_160), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g264 ( .A(n_61), .Y(n_264) );
INVx1_ASAP7_75t_L g149 ( .A(n_62), .Y(n_149) );
INVx1_ASAP7_75t_L g147 ( .A(n_64), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_65), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_66), .B(n_161), .Y(n_538) );
INVx1_ASAP7_75t_L g138 ( .A(n_67), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_68), .Y(n_118) );
AO32x2_ASAP7_75t_L g504 ( .A1(n_69), .A2(n_134), .A3(n_226), .B1(n_499), .B2(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g549 ( .A(n_70), .Y(n_549) );
INVx1_ASAP7_75t_L g487 ( .A(n_71), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_SL g186 ( .A1(n_72), .A2(n_160), .B(n_187), .C(n_188), .Y(n_186) );
INVxp67_ASAP7_75t_L g189 ( .A(n_73), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_74), .B(n_171), .Y(n_488) );
INVx1_ASAP7_75t_L g112 ( .A(n_75), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_76), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_77), .Y(n_750) );
INVx1_ASAP7_75t_L g257 ( .A(n_78), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_80), .A2(n_146), .B(n_151), .C(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_81), .B(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_82), .B(n_171), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_83), .B(n_200), .Y(n_214) );
INVx2_ASAP7_75t_L g136 ( .A(n_84), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_85), .B(n_187), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_86), .B(n_171), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_87), .A2(n_146), .B(n_151), .C(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g109 ( .A(n_88), .Y(n_109) );
OR2x2_ASAP7_75t_L g444 ( .A(n_88), .B(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g460 ( .A(n_88), .B(n_446), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_90), .A2(n_102), .B1(n_171), .B2(n_172), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_91), .B(n_164), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_92), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_93), .A2(n_146), .B(n_151), .C(n_229), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_94), .Y(n_236) );
INVx1_ASAP7_75t_L g185 ( .A(n_95), .Y(n_185) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_96), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_97), .B(n_200), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_98), .B(n_171), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_99), .B(n_134), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_100), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_101), .A2(n_141), .B(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g761 ( .A(n_104), .Y(n_761) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
OR2x2_ASAP7_75t_L g462 ( .A(n_109), .B(n_446), .Y(n_462) );
NOR2x2_ASAP7_75t_L g759 ( .A(n_109), .B(n_445), .Y(n_759) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AO21x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_119), .B(n_453), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_SL g760 ( .A(n_117), .Y(n_760) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_120), .B(n_451), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_122), .B1(n_125), .B2(n_442), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_125), .A2(n_464), .B1(n_755), .B2(n_756), .Y(n_754) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx2_ASAP7_75t_L g442 ( .A(n_126), .Y(n_442) );
AND3x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_364), .C(n_409), .Y(n_126) );
NOR4xp25_ASAP7_75t_L g127 ( .A(n_128), .B(n_287), .C(n_328), .D(n_345), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_191), .B(n_207), .C(n_249), .Y(n_128) );
OR2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_165), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_130), .B(n_192), .Y(n_191) );
NOR4xp25_ASAP7_75t_L g311 ( .A(n_130), .B(n_305), .C(n_312), .D(n_318), .Y(n_311) );
AND2x2_ASAP7_75t_L g384 ( .A(n_130), .B(n_273), .Y(n_384) );
AND2x2_ASAP7_75t_L g403 ( .A(n_130), .B(n_349), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_130), .B(n_398), .Y(n_412) );
AND2x2_ASAP7_75t_L g425 ( .A(n_130), .B(n_206), .Y(n_425) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_SL g270 ( .A(n_131), .Y(n_270) );
AND2x2_ASAP7_75t_L g277 ( .A(n_131), .B(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g327 ( .A(n_131), .B(n_166), .Y(n_327) );
AND2x2_ASAP7_75t_SL g338 ( .A(n_131), .B(n_273), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_131), .B(n_166), .Y(n_342) );
AND2x2_ASAP7_75t_L g351 ( .A(n_131), .B(n_276), .Y(n_351) );
BUFx2_ASAP7_75t_L g374 ( .A(n_131), .Y(n_374) );
AND2x2_ASAP7_75t_L g378 ( .A(n_131), .B(n_182), .Y(n_378) );
OA21x2_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_140), .B(n_163), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NOR2xp33_ASAP7_75t_SL g220 ( .A(n_133), .B(n_221), .Y(n_220) );
NAND3xp33_ASAP7_75t_L g514 ( .A(n_133), .B(n_499), .C(n_515), .Y(n_514) );
AO21x1_ASAP7_75t_L g552 ( .A1(n_133), .A2(n_515), .B(n_553), .Y(n_552) );
INVx4_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OA21x2_ASAP7_75t_L g182 ( .A1(n_134), .A2(n_183), .B(n_190), .Y(n_182) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_134), .A2(n_520), .B(n_528), .Y(n_519) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g168 ( .A(n_135), .Y(n_168) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x2_ASAP7_75t_SL g164 ( .A(n_136), .B(n_137), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
BUFx2_ASAP7_75t_L g240 ( .A(n_141), .Y(n_240) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_146), .Y(n_141) );
NAND2x1p5_ASAP7_75t_L g179 ( .A(n_142), .B(n_146), .Y(n_179) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
INVx1_ASAP7_75t_L g527 ( .A(n_143), .Y(n_527) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
INVx1_ASAP7_75t_L g172 ( .A(n_144), .Y(n_172) );
INVx1_ASAP7_75t_L g153 ( .A(n_145), .Y(n_153) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_145), .Y(n_156) );
INVx3_ASAP7_75t_L g159 ( .A(n_145), .Y(n_159) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_145), .Y(n_174) );
INVx1_ASAP7_75t_L g187 ( .A(n_145), .Y(n_187) );
INVx4_ASAP7_75t_SL g162 ( .A(n_146), .Y(n_162) );
OAI21xp5_ASAP7_75t_L g471 ( .A1(n_146), .A2(n_472), .B(n_476), .Y(n_471) );
OAI21xp5_ASAP7_75t_L g485 ( .A1(n_146), .A2(n_486), .B(n_489), .Y(n_485) );
BUFx3_ASAP7_75t_L g499 ( .A(n_146), .Y(n_499) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_146), .A2(n_521), .B(n_524), .Y(n_520) );
OAI21xp5_ASAP7_75t_L g530 ( .A1(n_146), .A2(n_531), .B(n_535), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_154), .C(n_162), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_150), .A2(n_162), .B(n_185), .C(n_186), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g241 ( .A1(n_150), .A2(n_162), .B(n_242), .C(n_243), .Y(n_241) );
INVx5_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x6_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_152), .Y(n_161) );
BUFx3_ASAP7_75t_L g218 ( .A(n_152), .Y(n_218) );
INVx1_ASAP7_75t_L g479 ( .A(n_152), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_155), .A2(n_477), .B(n_478), .Y(n_476) );
O2A1O1Ixp5_ASAP7_75t_L g548 ( .A1(n_155), .A2(n_536), .B(n_549), .C(n_550), .Y(n_548) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx4_ASAP7_75t_L g232 ( .A(n_156), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_156), .A2(n_496), .B1(n_497), .B2(n_498), .Y(n_495) );
OAI22xp5_ASAP7_75t_SL g505 ( .A1(n_156), .A2(n_159), .B1(n_506), .B2(n_507), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_156), .A2(n_497), .B1(n_516), .B2(n_517), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_159), .B(n_189), .Y(n_188) );
INVx5_ASAP7_75t_L g200 ( .A(n_159), .Y(n_200) );
O2A1O1Ixp5_ASAP7_75t_SL g486 ( .A1(n_160), .A2(n_200), .B(n_487), .C(n_488), .Y(n_486) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_161), .Y(n_233) );
OAI22xp33_ASAP7_75t_L g169 ( .A1(n_162), .A2(n_170), .B1(n_178), .B2(n_179), .Y(n_169) );
INVx1_ASAP7_75t_L g205 ( .A(n_164), .Y(n_205) );
INVx2_ASAP7_75t_L g226 ( .A(n_164), .Y(n_226) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_164), .A2(n_239), .B(n_248), .Y(n_238) );
OA21x2_ASAP7_75t_L g470 ( .A1(n_164), .A2(n_471), .B(n_480), .Y(n_470) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_164), .A2(n_485), .B(n_492), .Y(n_484) );
OR2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_182), .Y(n_165) );
AND2x2_ASAP7_75t_L g206 ( .A(n_166), .B(n_182), .Y(n_206) );
BUFx2_ASAP7_75t_L g280 ( .A(n_166), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_166), .A2(n_313), .B1(n_315), .B2(n_316), .Y(n_312) );
OR2x2_ASAP7_75t_L g334 ( .A(n_166), .B(n_194), .Y(n_334) );
AND2x2_ASAP7_75t_L g398 ( .A(n_166), .B(n_276), .Y(n_398) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g266 ( .A(n_167), .B(n_194), .Y(n_266) );
AND2x2_ASAP7_75t_L g273 ( .A(n_167), .B(n_182), .Y(n_273) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_167), .Y(n_315) );
OR2x2_ASAP7_75t_L g350 ( .A(n_167), .B(n_193), .Y(n_350) );
AO21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_180), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_168), .B(n_181), .Y(n_180) );
AO21x2_ASAP7_75t_L g194 ( .A1(n_168), .A2(n_195), .B(n_203), .Y(n_194) );
INVx2_ASAP7_75t_L g219 ( .A(n_168), .Y(n_219) );
INVx2_ASAP7_75t_L g202 ( .A(n_171), .Y(n_202) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OAI22xp5_ASAP7_75t_SL g173 ( .A1(n_174), .A2(n_175), .B1(n_176), .B2(n_177), .Y(n_173) );
INVx2_ASAP7_75t_L g176 ( .A(n_174), .Y(n_176) );
INVx4_ASAP7_75t_L g244 ( .A(n_174), .Y(n_244) );
OAI21xp5_ASAP7_75t_L g195 ( .A1(n_179), .A2(n_196), .B(n_197), .Y(n_195) );
OAI21xp5_ASAP7_75t_L g256 ( .A1(n_179), .A2(n_257), .B(n_258), .Y(n_256) );
INVx1_ASAP7_75t_L g269 ( .A(n_182), .Y(n_269) );
INVx3_ASAP7_75t_L g278 ( .A(n_182), .Y(n_278) );
BUFx2_ASAP7_75t_L g302 ( .A(n_182), .Y(n_302) );
AND2x2_ASAP7_75t_L g335 ( .A(n_182), .B(n_270), .Y(n_335) );
INVx1_ASAP7_75t_L g475 ( .A(n_187), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_191), .A2(n_421), .B1(n_422), .B2(n_423), .Y(n_420) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_206), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_193), .B(n_278), .Y(n_282) );
INVx1_ASAP7_75t_L g310 ( .A(n_193), .Y(n_310) );
INVx3_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx3_ASAP7_75t_L g276 ( .A(n_194), .Y(n_276) );
O2A1O1Ixp33_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_201), .C(n_202), .Y(n_198) );
INVx2_ASAP7_75t_L g497 ( .A(n_200), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_200), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_200), .A2(n_546), .B(n_547), .Y(n_545) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_202), .A2(n_532), .B(n_533), .C(n_534), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_205), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_205), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g288 ( .A(n_206), .Y(n_288) );
NAND2x1_ASAP7_75t_SL g207 ( .A(n_208), .B(n_222), .Y(n_207) );
AND2x2_ASAP7_75t_L g286 ( .A(n_208), .B(n_237), .Y(n_286) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_208), .Y(n_360) );
AND2x2_ASAP7_75t_L g387 ( .A(n_208), .B(n_307), .Y(n_387) );
AND2x2_ASAP7_75t_L g395 ( .A(n_208), .B(n_357), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_208), .B(n_252), .Y(n_422) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g253 ( .A(n_209), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g271 ( .A(n_209), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g292 ( .A(n_209), .Y(n_292) );
INVx1_ASAP7_75t_L g298 ( .A(n_209), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_209), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g331 ( .A(n_209), .B(n_255), .Y(n_331) );
OR2x2_ASAP7_75t_L g369 ( .A(n_209), .B(n_324), .Y(n_369) );
AOI32xp33_ASAP7_75t_L g381 ( .A1(n_209), .A2(n_382), .A3(n_385), .B1(n_386), .B2(n_387), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_209), .B(n_357), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_209), .B(n_317), .Y(n_432) );
OR2x6_ASAP7_75t_L g209 ( .A(n_210), .B(n_220), .Y(n_209) );
AOI21xp5_ASAP7_75t_SL g210 ( .A1(n_211), .A2(n_212), .B(n_219), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_216), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_216), .A2(n_260), .B(n_261), .Y(n_259) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g247 ( .A(n_218), .Y(n_247) );
INVx1_ASAP7_75t_L g262 ( .A(n_219), .Y(n_262) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_219), .A2(n_530), .B(n_539), .Y(n_529) );
OA21x2_ASAP7_75t_L g543 ( .A1(n_219), .A2(n_544), .B(n_551), .Y(n_543) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
OR2x2_ASAP7_75t_L g343 ( .A(n_223), .B(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_237), .Y(n_223) );
INVx1_ASAP7_75t_L g305 ( .A(n_224), .Y(n_305) );
AND2x2_ASAP7_75t_L g307 ( .A(n_224), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_224), .B(n_254), .Y(n_324) );
AND2x2_ASAP7_75t_L g357 ( .A(n_224), .B(n_333), .Y(n_357) );
AND2x2_ASAP7_75t_L g394 ( .A(n_224), .B(n_255), .Y(n_394) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g252 ( .A(n_225), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_225), .B(n_254), .Y(n_284) );
AND2x2_ASAP7_75t_L g291 ( .A(n_225), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g332 ( .A(n_225), .B(n_333), .Y(n_332) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_235), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_228), .B(n_234), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_233), .Y(n_229) );
INVx2_ASAP7_75t_L g308 ( .A(n_237), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_237), .B(n_254), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_237), .B(n_299), .Y(n_380) );
INVx1_ASAP7_75t_L g402 ( .A(n_237), .Y(n_402) );
INVx1_ASAP7_75t_L g419 ( .A(n_237), .Y(n_419) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g272 ( .A(n_238), .B(n_254), .Y(n_272) );
AND2x2_ASAP7_75t_L g294 ( .A(n_238), .B(n_255), .Y(n_294) );
INVx1_ASAP7_75t_L g333 ( .A(n_238), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_244), .B(n_246), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_244), .A2(n_490), .B(n_491), .Y(n_489) );
INVx1_ASAP7_75t_L g534 ( .A(n_244), .Y(n_534) );
AOI221x1_ASAP7_75t_SL g249 ( .A1(n_250), .A2(n_265), .B1(n_271), .B2(n_273), .C(n_274), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_250), .A2(n_338), .B1(n_405), .B2(n_406), .Y(n_404) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_253), .Y(n_250) );
AND2x2_ASAP7_75t_L g296 ( .A(n_251), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g391 ( .A(n_251), .B(n_271), .Y(n_391) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g347 ( .A(n_252), .B(n_272), .Y(n_347) );
INVx1_ASAP7_75t_L g359 ( .A(n_253), .Y(n_359) );
AND2x2_ASAP7_75t_L g370 ( .A(n_253), .B(n_357), .Y(n_370) );
AND2x2_ASAP7_75t_L g437 ( .A(n_253), .B(n_332), .Y(n_437) );
INVx2_ASAP7_75t_L g299 ( .A(n_254), .Y(n_299) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_262), .B(n_263), .Y(n_255) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_266), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g389 ( .A(n_266), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_267), .B(n_350), .Y(n_353) );
INVx3_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_268), .A2(n_389), .B(n_434), .Y(n_433) );
AND2x4_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
NOR2xp33_ASAP7_75t_SL g411 ( .A(n_271), .B(n_297), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_272), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g363 ( .A(n_272), .B(n_291), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_272), .B(n_298), .Y(n_440) );
AND2x2_ASAP7_75t_L g309 ( .A(n_273), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g376 ( .A(n_273), .Y(n_376) );
AOI21xp33_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_279), .B(n_283), .Y(n_274) );
NAND2x1_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_276), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g325 ( .A(n_276), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g337 ( .A(n_276), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_276), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g361 ( .A(n_277), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_277), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_277), .B(n_280), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
AOI211xp5_ASAP7_75t_L g348 ( .A1(n_280), .A2(n_319), .B(n_349), .C(n_351), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_280), .A2(n_367), .B1(n_370), .B2(n_371), .C(n_375), .Y(n_366) );
AND2x2_ASAP7_75t_L g362 ( .A(n_281), .B(n_315), .Y(n_362) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g322 ( .A(n_286), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g393 ( .A(n_286), .B(n_394), .Y(n_393) );
OAI211xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_289), .B(n_295), .C(n_320), .Y(n_287) );
NAND3xp33_ASAP7_75t_SL g406 ( .A(n_288), .B(n_407), .C(n_408), .Y(n_406) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_293), .Y(n_289) );
OR2x2_ASAP7_75t_L g379 ( .A(n_290), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_300), .B1(n_303), .B2(n_309), .C(n_311), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_297), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_297), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g319 ( .A(n_302), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_302), .A2(n_359), .B1(n_360), .B2(n_361), .Y(n_358) );
OR2x2_ASAP7_75t_L g439 ( .A(n_302), .B(n_350), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_304), .B(n_306), .Y(n_303) );
INVxp67_ASAP7_75t_L g413 ( .A(n_305), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_307), .B(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g314 ( .A(n_308), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_310), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_310), .B(n_357), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_310), .B(n_377), .Y(n_416) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_314), .Y(n_340) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g430 ( .A(n_319), .B(n_350), .Y(n_430) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_325), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_SL g408 ( .A(n_325), .Y(n_408) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OAI322xp33_ASAP7_75t_SL g328 ( .A1(n_329), .A2(n_334), .A3(n_335), .B1(n_336), .B2(n_339), .C1(n_341), .C2(n_343), .Y(n_328) );
OAI322xp33_ASAP7_75t_L g410 ( .A1(n_329), .A2(n_411), .A3(n_412), .B1(n_413), .B2(n_414), .C1(n_415), .C2(n_417), .Y(n_410) );
CKINVDCx16_ASAP7_75t_R g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx4_ASAP7_75t_L g344 ( .A(n_331), .Y(n_344) );
AND2x2_ASAP7_75t_L g405 ( .A(n_331), .B(n_357), .Y(n_405) );
AND2x2_ASAP7_75t_L g418 ( .A(n_331), .B(n_419), .Y(n_418) );
CKINVDCx16_ASAP7_75t_R g429 ( .A(n_334), .Y(n_429) );
INVx1_ASAP7_75t_L g407 ( .A(n_335), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
OR2x2_ASAP7_75t_L g341 ( .A(n_337), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g424 ( .A(n_337), .B(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_337), .B(n_378), .Y(n_435) );
OR2x2_ASAP7_75t_L g368 ( .A(n_340), .B(n_369), .Y(n_368) );
INVxp33_ASAP7_75t_L g385 ( .A(n_340), .Y(n_385) );
OAI221xp5_ASAP7_75t_SL g345 ( .A1(n_344), .A2(n_346), .B1(n_348), .B2(n_352), .C(n_354), .Y(n_345) );
NOR2xp67_ASAP7_75t_L g401 ( .A(n_344), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g428 ( .A(n_344), .Y(n_428) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
INVx3_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
AOI322xp5_ASAP7_75t_L g392 ( .A1(n_351), .A2(n_376), .A3(n_393), .B1(n_395), .B2(n_396), .C1(n_399), .C2(n_403), .Y(n_392) );
INVxp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_358), .B1(n_362), .B2(n_363), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_365), .B(n_388), .Y(n_364) );
NAND2xp5_ASAP7_75t_SL g365 ( .A(n_366), .B(n_381), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_369), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
NAND2xp33_ASAP7_75t_SL g386 ( .A(n_372), .B(n_383), .Y(n_386) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
OAI322xp33_ASAP7_75t_L g426 ( .A1(n_374), .A2(n_427), .A3(n_429), .B1(n_430), .B2(n_431), .C1(n_433), .C2(n_436), .Y(n_426) );
AOI21xp33_ASAP7_75t_SL g375 ( .A1(n_376), .A2(n_377), .B(n_379), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_384), .B(n_432), .Y(n_441) );
OAI211xp5_ASAP7_75t_SL g388 ( .A1(n_389), .A2(n_390), .B(n_392), .C(n_404), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NOR4xp25_ASAP7_75t_L g409 ( .A(n_410), .B(n_420), .C(n_426), .D(n_438), .Y(n_409) );
INVxp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
CKINVDCx14_ASAP7_75t_R g436 ( .A(n_437), .Y(n_436) );
OAI21xp5_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_440), .B(n_441), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_442), .A2(n_457), .B1(n_461), .B2(n_463), .Y(n_456) );
INVx1_ASAP7_75t_L g451 ( .A(n_443), .Y(n_451) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
AOI21xp33_ASAP7_75t_L g453 ( .A1(n_452), .A2(n_454), .B(n_760), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g755 ( .A(n_460), .Y(n_755) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx6_ASAP7_75t_L g756 ( .A(n_462), .Y(n_756) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_668), .Y(n_464) );
NAND5xp2_ASAP7_75t_L g465 ( .A(n_466), .B(n_587), .C(n_602), .D(n_628), .E(n_650), .Y(n_465) );
NOR2xp33_ASAP7_75t_SL g466 ( .A(n_467), .B(n_567), .Y(n_466) );
OAI221xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_508), .B1(n_540), .B2(n_556), .C(n_557), .Y(n_467) );
NOR2xp33_ASAP7_75t_SL g468 ( .A(n_469), .B(n_500), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_469), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_SL g744 ( .A(n_469), .Y(n_744) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_481), .Y(n_469) );
INVx1_ASAP7_75t_L g584 ( .A(n_470), .Y(n_584) );
AND2x2_ASAP7_75t_L g586 ( .A(n_470), .B(n_494), .Y(n_586) );
AND2x2_ASAP7_75t_L g596 ( .A(n_470), .B(n_493), .Y(n_596) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_470), .Y(n_614) );
INVx1_ASAP7_75t_L g624 ( .A(n_470), .Y(n_624) );
OR2x2_ASAP7_75t_L g662 ( .A(n_470), .B(n_561), .Y(n_662) );
INVx2_ASAP7_75t_L g712 ( .A(n_470), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_470), .B(n_560), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B(n_475), .Y(n_472) );
NOR2xp67_ASAP7_75t_L g481 ( .A(n_482), .B(n_493), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_483), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_483), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_SL g644 ( .A(n_483), .B(n_584), .Y(n_644) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_484), .Y(n_502) );
INVx2_ASAP7_75t_L g561 ( .A(n_484), .Y(n_561) );
OR2x2_ASAP7_75t_L g623 ( .A(n_484), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g562 ( .A(n_493), .B(n_504), .Y(n_562) );
AND2x2_ASAP7_75t_L g579 ( .A(n_493), .B(n_559), .Y(n_579) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g503 ( .A(n_494), .B(n_504), .Y(n_503) );
BUFx2_ASAP7_75t_L g582 ( .A(n_494), .Y(n_582) );
AND2x2_ASAP7_75t_L g711 ( .A(n_494), .B(n_712), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_497), .A2(n_525), .B(n_526), .Y(n_524) );
O2A1O1Ixp33_ASAP7_75t_L g535 ( .A1(n_497), .A2(n_536), .B(n_537), .C(n_538), .Y(n_535) );
OAI21xp5_ASAP7_75t_L g544 ( .A1(n_499), .A2(n_545), .B(n_548), .Y(n_544) );
INVx1_ASAP7_75t_L g556 ( .A(n_500), .Y(n_556) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_503), .Y(n_500) );
AND2x2_ASAP7_75t_L g674 ( .A(n_501), .B(n_562), .Y(n_674) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g675 ( .A(n_502), .B(n_586), .Y(n_675) );
O2A1O1Ixp33_ASAP7_75t_L g642 ( .A1(n_503), .A2(n_643), .B(n_645), .C(n_647), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_503), .B(n_643), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g715 ( .A1(n_503), .A2(n_573), .B1(n_716), .B2(n_717), .C(n_719), .Y(n_715) );
INVx1_ASAP7_75t_L g559 ( .A(n_504), .Y(n_559) );
INVx1_ASAP7_75t_L g595 ( .A(n_504), .Y(n_595) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_504), .Y(n_604) );
INVx1_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_518), .Y(n_509) );
AND2x2_ASAP7_75t_L g621 ( .A(n_510), .B(n_566), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_510), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_511), .B(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g713 ( .A(n_511), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g745 ( .A(n_511), .Y(n_745) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx3_ASAP7_75t_L g575 ( .A(n_512), .Y(n_575) );
AND2x2_ASAP7_75t_L g601 ( .A(n_512), .B(n_555), .Y(n_601) );
NOR2x1_ASAP7_75t_L g610 ( .A(n_512), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g617 ( .A(n_512), .B(n_618), .Y(n_617) );
AND2x4_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
INVx1_ASAP7_75t_L g553 ( .A(n_513), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_518), .B(n_657), .Y(n_692) );
INVx1_ASAP7_75t_SL g696 ( .A(n_518), .Y(n_696) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_529), .Y(n_518) );
INVx3_ASAP7_75t_L g555 ( .A(n_519), .Y(n_555) );
AND2x2_ASAP7_75t_L g566 ( .A(n_519), .B(n_543), .Y(n_566) );
AND2x2_ASAP7_75t_L g588 ( .A(n_519), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g633 ( .A(n_519), .B(n_627), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_519), .B(n_565), .Y(n_714) );
INVx2_ASAP7_75t_L g536 ( .A(n_527), .Y(n_536) );
AND2x2_ASAP7_75t_L g554 ( .A(n_529), .B(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g565 ( .A(n_529), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_529), .B(n_543), .Y(n_590) );
AND2x2_ASAP7_75t_L g626 ( .A(n_529), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_554), .Y(n_541) );
INVx1_ASAP7_75t_L g606 ( .A(n_542), .Y(n_606) );
AND2x2_ASAP7_75t_L g648 ( .A(n_542), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_542), .B(n_569), .Y(n_654) );
AOI21xp5_ASAP7_75t_SL g728 ( .A1(n_542), .A2(n_560), .B(n_583), .Y(n_728) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_552), .Y(n_542) );
OR2x2_ASAP7_75t_L g571 ( .A(n_543), .B(n_552), .Y(n_571) );
AND2x2_ASAP7_75t_L g618 ( .A(n_543), .B(n_555), .Y(n_618) );
INVx2_ASAP7_75t_L g627 ( .A(n_543), .Y(n_627) );
INVx1_ASAP7_75t_L g733 ( .A(n_543), .Y(n_733) );
AND2x2_ASAP7_75t_L g657 ( .A(n_552), .B(n_627), .Y(n_657) );
INVx1_ASAP7_75t_L g682 ( .A(n_552), .Y(n_682) );
AND2x2_ASAP7_75t_L g591 ( .A(n_554), .B(n_575), .Y(n_591) );
AND2x2_ASAP7_75t_L g603 ( .A(n_554), .B(n_604), .Y(n_603) );
INVx2_ASAP7_75t_SL g721 ( .A(n_554), .Y(n_721) );
INVx2_ASAP7_75t_L g611 ( .A(n_555), .Y(n_611) );
AND2x2_ASAP7_75t_L g649 ( .A(n_555), .B(n_565), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_555), .B(n_733), .Y(n_732) );
OAI21xp33_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_562), .B(n_563), .Y(n_557) );
AND2x2_ASAP7_75t_L g664 ( .A(n_558), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g718 ( .A(n_558), .Y(n_718) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
INVx1_ASAP7_75t_L g638 ( .A(n_559), .Y(n_638) );
BUFx2_ASAP7_75t_L g737 ( .A(n_559), .Y(n_737) );
BUFx2_ASAP7_75t_L g608 ( .A(n_560), .Y(n_608) );
AND2x2_ASAP7_75t_L g710 ( .A(n_560), .B(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g693 ( .A(n_561), .Y(n_693) );
AND2x4_ASAP7_75t_L g620 ( .A(n_562), .B(n_583), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_562), .B(n_644), .Y(n_656) );
AOI32xp33_ASAP7_75t_L g580 ( .A1(n_563), .A2(n_581), .A3(n_583), .B1(n_585), .B2(n_586), .Y(n_580) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .Y(n_563) );
INVx3_ASAP7_75t_L g569 ( .A(n_564), .Y(n_569) );
OR2x2_ASAP7_75t_L g705 ( .A(n_564), .B(n_661), .Y(n_705) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g574 ( .A(n_565), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g681 ( .A(n_565), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g573 ( .A(n_566), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g585 ( .A(n_566), .B(n_575), .Y(n_585) );
INVx1_ASAP7_75t_L g706 ( .A(n_566), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_566), .B(n_681), .Y(n_739) );
A2O1A1Ixp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_572), .B(n_576), .C(n_580), .Y(n_567) );
OAI322xp33_ASAP7_75t_L g676 ( .A1(n_568), .A2(n_613), .A3(n_677), .B1(n_679), .B2(n_683), .C1(n_684), .C2(n_688), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVxp67_ASAP7_75t_L g641 ( .A(n_569), .Y(n_641) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g695 ( .A(n_571), .B(n_696), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_571), .B(n_611), .Y(n_742) );
INVxp67_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g634 ( .A(n_574), .Y(n_634) );
OR2x2_ASAP7_75t_L g720 ( .A(n_575), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_578), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g629 ( .A(n_579), .B(n_608), .Y(n_629) );
AND2x2_ASAP7_75t_L g700 ( .A(n_579), .B(n_613), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_579), .B(n_687), .Y(n_722) );
AOI221xp5_ASAP7_75t_L g587 ( .A1(n_581), .A2(n_588), .B1(n_591), .B2(n_592), .C(n_597), .Y(n_587) );
OR2x2_ASAP7_75t_L g598 ( .A(n_581), .B(n_594), .Y(n_598) );
AND2x2_ASAP7_75t_L g686 ( .A(n_581), .B(n_687), .Y(n_686) );
AOI32xp33_ASAP7_75t_L g725 ( .A1(n_581), .A2(n_611), .A3(n_726), .B1(n_727), .B2(n_730), .Y(n_725) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND3xp33_ASAP7_75t_L g659 ( .A(n_582), .B(n_618), .C(n_641), .Y(n_659) );
AND2x2_ASAP7_75t_L g685 ( .A(n_582), .B(n_678), .Y(n_685) );
INVxp67_ASAP7_75t_L g665 ( .A(n_583), .Y(n_665) );
BUFx3_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_586), .B(n_638), .Y(n_694) );
INVx2_ASAP7_75t_L g704 ( .A(n_586), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_586), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g673 ( .A(n_589), .Y(n_673) );
OR2x2_ASAP7_75t_L g599 ( .A(n_590), .B(n_600), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_592), .B(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_596), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_595), .Y(n_678) );
AND2x2_ASAP7_75t_L g637 ( .A(n_596), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g683 ( .A(n_596), .Y(n_683) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_596), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
AOI21xp33_ASAP7_75t_SL g622 ( .A1(n_598), .A2(n_623), .B(n_625), .Y(n_622) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g716 ( .A(n_601), .B(n_626), .Y(n_716) );
AOI211xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_605), .B(n_615), .C(n_622), .Y(n_602) );
AND2x2_ASAP7_75t_L g646 ( .A(n_604), .B(n_614), .Y(n_646) );
INVx2_ASAP7_75t_L g661 ( .A(n_604), .Y(n_661) );
OR2x2_ASAP7_75t_L g699 ( .A(n_604), .B(n_662), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_604), .B(n_742), .Y(n_741) );
AOI211xp5_ASAP7_75t_SL g605 ( .A1(n_606), .A2(n_607), .B(n_609), .C(n_612), .Y(n_605) );
INVxp67_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_608), .B(n_646), .Y(n_645) );
OAI211xp5_ASAP7_75t_L g727 ( .A1(n_609), .A2(n_704), .B(n_728), .C(n_729), .Y(n_727) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2x1p5_ASAP7_75t_L g625 ( .A(n_610), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g667 ( .A(n_611), .B(n_657), .Y(n_667) );
INVx1_ASAP7_75t_L g672 ( .A(n_611), .Y(n_672) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g615 ( .A(n_616), .B(n_619), .Y(n_615) );
INVxp33_ASAP7_75t_L g723 ( .A(n_617), .Y(n_723) );
AND2x2_ASAP7_75t_L g702 ( .A(n_618), .B(n_681), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_623), .A2(n_685), .B(n_686), .Y(n_684) );
OAI322xp33_ASAP7_75t_L g703 ( .A1(n_625), .A2(n_704), .A3(n_705), .B1(n_706), .B2(n_707), .C1(n_709), .C2(n_713), .Y(n_703) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B1(n_635), .B2(n_639), .C(n_642), .Y(n_628) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g680 ( .A(n_633), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g724 ( .A(n_637), .Y(n_724) );
INVxp67_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_640), .B(n_660), .Y(n_726) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g689 ( .A(n_649), .B(n_657), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_653), .B1(n_655), .B2(n_657), .C(n_658), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_653), .A2(n_670), .B1(n_674), .B2(n_675), .C(n_676), .Y(n_669) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVxp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_657), .B(n_672), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B1(n_663), .B2(n_666), .Y(n_658) );
OR2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
INVx2_ASAP7_75t_SL g687 ( .A(n_662), .Y(n_687) );
INVxp67_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND5xp2_ASAP7_75t_L g668 ( .A(n_669), .B(n_690), .C(n_715), .D(n_725), .E(n_735), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_671), .B(n_673), .Y(n_670) );
NOR4xp25_ASAP7_75t_L g743 ( .A(n_672), .B(n_678), .C(n_744), .D(n_745), .Y(n_743) );
AOI221xp5_ASAP7_75t_L g735 ( .A1(n_675), .A2(n_736), .B1(n_738), .B2(n_740), .C(n_743), .Y(n_735) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g734 ( .A(n_681), .Y(n_734) );
OAI322xp33_ASAP7_75t_L g691 ( .A1(n_685), .A2(n_692), .A3(n_693), .B1(n_694), .B2(n_695), .C1(n_697), .C2(n_701), .Y(n_691) );
INVx1_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_703), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_700), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g736 ( .A(n_711), .B(n_737), .Y(n_736) );
OAI22xp33_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_722), .B1(n_723), .B2(n_724), .Y(n_719) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
OR2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_734), .Y(n_731) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVxp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
endmodule