module fake_jpeg_8372_n_229 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_SL g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_36),
.B(n_48),
.Y(n_72)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_31),
.Y(n_57)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

CKINVDCx6p67_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_50),
.Y(n_75)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_40),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_52),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_48),
.B(n_21),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_67),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_23),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_54),
.A2(n_21),
.B(n_32),
.Y(n_101)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_59),
.Y(n_74)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_65),
.Y(n_95)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_30),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_31),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_90),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_30),
.B(n_24),
.C(n_25),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_78),
.B(n_79),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_30),
.B(n_24),
.C(n_25),
.Y(n_79)
);

O2A1O1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_36),
.B(n_23),
.C(n_29),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_81),
.Y(n_125)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_93),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_39),
.B(n_45),
.C(n_43),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_85),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_64),
.A2(n_45),
.B1(n_37),
.B2(n_43),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_34),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_37),
.B1(n_42),
.B2(n_46),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_86),
.A2(n_87),
.B1(n_61),
.B2(n_63),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_49),
.A2(n_42),
.B1(n_39),
.B2(n_29),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_34),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_91),
.C(n_35),
.Y(n_116)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_97),
.Y(n_118)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_103),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_56),
.Y(n_97)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_0),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_101),
.B(n_28),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_51),
.A2(n_18),
.B(n_32),
.Y(n_102)
);

NOR3xp33_ASAP7_75t_SL g110 ( 
.A(n_102),
.B(n_18),
.C(n_39),
.Y(n_110)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_107),
.B(n_112),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_119),
.B1(n_92),
.B2(n_90),
.Y(n_134)
);

NAND2xp33_ASAP7_75t_SL g144 ( 
.A(n_110),
.B(n_31),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_33),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_115),
.B(n_117),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_87),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_33),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_85),
.A2(n_73),
.B1(n_27),
.B2(n_28),
.Y(n_119)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_124),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_73),
.C(n_27),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_80),
.C(n_75),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_78),
.B(n_101),
.Y(n_123)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_102),
.B(n_22),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_35),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_22),
.Y(n_128)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_100),
.B1(n_88),
.B2(n_83),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_130),
.A2(n_135),
.B1(n_143),
.B2(n_144),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_119),
.C(n_108),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_141),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_125),
.A2(n_109),
.B1(n_122),
.B2(n_123),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_77),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_138),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_140),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_95),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_89),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_147),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_125),
.A2(n_86),
.B1(n_99),
.B2(n_98),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_99),
.B1(n_20),
.B2(n_18),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_150),
.B1(n_128),
.B2(n_117),
.Y(n_158)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_15),
.Y(n_148)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_121),
.A2(n_94),
.B1(n_15),
.B2(n_13),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

OAI32xp33_ASAP7_75t_L g153 ( 
.A1(n_136),
.A2(n_127),
.A3(n_114),
.B1(n_124),
.B2(n_116),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_149),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_107),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_154),
.A2(n_157),
.B(n_162),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_163),
.C(n_169),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_140),
.B(n_143),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_161),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_141),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_106),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_108),
.C(n_112),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_120),
.B1(n_111),
.B2(n_105),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_165),
.A2(n_156),
.B1(n_155),
.B2(n_132),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_139),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_166),
.B(n_146),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_131),
.A2(n_1),
.B(n_2),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_1),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_11),
.C(n_10),
.Y(n_169)
);

OAI322xp33_ASAP7_75t_L g171 ( 
.A1(n_152),
.A2(n_170),
.A3(n_153),
.B1(n_157),
.B2(n_162),
.C1(n_154),
.C2(n_163),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_177),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_159),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_178),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_167),
.B(n_158),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_134),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_156),
.C(n_165),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_146),
.Y(n_180)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_180),
.Y(n_198)
);

OA21x2_ASAP7_75t_SL g181 ( 
.A1(n_154),
.A2(n_147),
.B(n_150),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_184),
.Y(n_194)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_182),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_183),
.A2(n_186),
.B1(n_1),
.B2(n_2),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_185),
.A2(n_162),
.B1(n_169),
.B2(n_132),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_168),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_192),
.C(n_195),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_190),
.A2(n_183),
.B1(n_184),
.B2(n_5),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_173),
.C(n_177),
.Y(n_192)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_193),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_10),
.C(n_4),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g196 ( 
.A(n_182),
.Y(n_196)
);

INVx11_ASAP7_75t_L g201 ( 
.A(n_196),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_189),
.A2(n_175),
.B(n_174),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_199),
.B(n_4),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_179),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_203),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_178),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_175),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_207),
.C(n_195),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_188),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_3),
.C(n_4),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_196),
.Y(n_209)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_212),
.C(n_207),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_197),
.Y(n_211)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_211),
.Y(n_218)
);

AOI322xp5_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_191),
.A3(n_198),
.B1(n_188),
.B2(n_7),
.C1(n_3),
.C2(n_5),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_213),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_214),
.A2(n_200),
.B(n_206),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_215),
.B(n_205),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_208),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_220),
.Y(n_224)
);

O2A1O1Ixp33_ASAP7_75t_SL g225 ( 
.A1(n_221),
.A2(n_222),
.B(n_223),
.C(n_219),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_205),
.C(n_209),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_204),
.B1(n_5),
.B2(n_8),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_8),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_222),
.C(n_219),
.Y(n_226)
);

NOR2xp67_ASAP7_75t_SL g228 ( 
.A(n_226),
.B(n_227),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_8),
.Y(n_229)
);


endmodule