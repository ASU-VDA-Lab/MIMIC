module real_jpeg_7549_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_288;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_249;
wire n_286;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_285;
wire n_160;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_195;
wire n_61;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_228;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_240;
wire n_297;
wire n_55;
wire n_185;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_209;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_295;
wire n_202;
wire n_133;
wire n_213;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_0),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_0),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_0),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_0),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_0),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_0),
.B(n_248),
.Y(n_247)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_1),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_1),
.B(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_1),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g216 ( 
.A(n_1),
.B(n_217),
.Y(n_216)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_3),
.B(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_3),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_3),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_3),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_3),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_3),
.B(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_4),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_4),
.Y(n_238)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_6),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_6),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g171 ( 
.A(n_6),
.B(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_7),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_7),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_7),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_7),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_8),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g158 ( 
.A(n_8),
.Y(n_158)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_11),
.A2(n_28),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_11),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_11),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_11),
.B(n_49),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_11),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_11),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_11),
.B(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_12),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_12),
.Y(n_156)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_12),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_13),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_13),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_13),
.B(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_13),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_13),
.B(n_207),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_13),
.B(n_156),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_14),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_15),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_15),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_15),
.B(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_182),
.B1(n_296),
.B2(n_297),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_18),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_180),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_141),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_20),
.B(n_141),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_71),
.C(n_116),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_21),
.B(n_294),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_50),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_34),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_23),
.B(n_34),
.C(n_50),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B(n_32),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_25),
.B(n_223),
.Y(n_222)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_32),
.B(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_46),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_40),
.B1(n_41),
.B2(n_45),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_36),
.B(n_41),
.C(n_46),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_38),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_39),
.Y(n_225)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_63),
.C(n_66),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_51),
.A2(n_52),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_58),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_53),
.A2(n_58),
.B1(n_150),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_53),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_57),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_58),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_58),
.Y(n_150)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_63),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_70),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_71),
.B(n_116),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_90),
.C(n_106),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_72),
.B(n_287),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_84),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_74),
.B(n_81),
.C(n_84),
.Y(n_140)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_78),
.B(n_127),
.Y(n_147)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_89),
.Y(n_174)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_89),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_90),
.A2(n_106),
.B1(n_107),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_90),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_97),
.C(n_102),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_91),
.A2(n_92),
.B1(n_102),
.B2(n_103),
.Y(n_275)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_97),
.B(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_98),
.B(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_101),
.Y(n_192)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_105),
.Y(n_202)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_112),
.B2(n_113),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_136),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_137),
.C(n_140),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_124),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_118),
.B(n_125),
.C(n_135),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_130),
.B2(n_135),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_159),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_153),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_179),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_170),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx3_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.Y(n_170)
);

INVx4_ASAP7_75t_SL g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_182),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_291),
.B(n_295),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_277),
.B(n_290),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_263),
.B(n_276),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_230),
.B(n_262),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_220),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_187),
.B(n_220),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_203),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_188),
.B(n_204),
.C(n_214),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_193),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_189),
.B(n_194),
.C(n_199),
.Y(n_273)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_199),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_214),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_209),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_209),
.Y(n_221)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx8_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_214)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_216),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_216),
.B(n_218),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.C(n_226),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_222),
.A2(n_226),
.B1(n_227),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_222),
.Y(n_260)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_256),
.B(n_261),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_246),
.B(n_255),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_243),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_243),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_239),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_239),
.Y(n_257)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_258),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_265),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_272),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_273),
.C(n_274),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_271),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_269),
.C(n_271),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_289),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_289),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_286),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_283),
.C(n_286),
.Y(n_292)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_284),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_293),
.Y(n_295)
);


endmodule