module fake_jpeg_14481_n_579 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_579);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_579;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_13),
.B(n_4),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVxp33_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_12),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_55),
.B(n_69),
.Y(n_124)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_56),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_18),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_60),
.B(n_63),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_62),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_19),
.B(n_16),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_65),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_66),
.B(n_70),
.Y(n_152)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_29),
.B(n_16),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_29),
.B(n_30),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_74),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_75),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_30),
.B(n_15),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_76),
.B(n_79),
.Y(n_137)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_78),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_40),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_43),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_80),
.B(n_87),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_84),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_85),
.Y(n_168)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_40),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_20),
.B(n_15),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_91),
.B(n_98),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_21),
.B(n_14),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_92),
.B(n_93),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_40),
.Y(n_93)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_33),
.B(n_14),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_40),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_99),
.Y(n_119)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_38),
.B(n_0),
.Y(n_102)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_38),
.Y(n_103)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_104),
.Y(n_163)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

INVx11_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_27),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_106),
.Y(n_143)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_107),
.Y(n_167)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_20),
.Y(n_108)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_38),
.Y(n_109)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_109),
.Y(n_169)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_34),
.Y(n_110)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_57),
.A2(n_27),
.B1(n_45),
.B2(n_53),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_114),
.A2(n_88),
.B1(n_95),
.B2(n_97),
.Y(n_196)
);

AND2x4_ASAP7_75t_L g116 ( 
.A(n_71),
.B(n_77),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_116),
.B(n_104),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_94),
.A2(n_50),
.B1(n_31),
.B2(n_51),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_123),
.A2(n_153),
.B1(n_106),
.B2(n_72),
.Y(n_205)
);

BUFx2_ASAP7_75t_R g132 ( 
.A(n_56),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_132),
.B(n_6),
.Y(n_238)
);

INVx4_ASAP7_75t_SL g135 ( 
.A(n_108),
.Y(n_135)
);

INVx4_ASAP7_75t_SL g229 ( 
.A(n_135),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_31),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_61),
.Y(n_181)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_148),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_74),
.A2(n_44),
.B1(n_49),
.B2(n_53),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_149),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_236)
);

BUFx24_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

BUFx2_ASAP7_75t_SL g230 ( 
.A(n_151),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_81),
.A2(n_50),
.B1(n_51),
.B2(n_45),
.Y(n_153)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_73),
.Y(n_166)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_58),
.Y(n_171)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_171),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_67),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_172),
.B(n_173),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_78),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_84),
.Y(n_174)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_85),
.Y(n_175)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_175),
.Y(n_180)
);

INVx5_ASAP7_75t_SL g176 ( 
.A(n_61),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_176),
.Y(n_222)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_178),
.Y(n_243)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_179),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_181),
.B(n_183),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_124),
.B(n_47),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_182),
.B(n_184),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_155),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_164),
.B(n_152),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_130),
.Y(n_185)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_185),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_186),
.B(n_226),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_137),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_187),
.B(n_198),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_150),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_188),
.Y(n_271)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_189),
.Y(n_269)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_190),
.Y(n_275)
);

CKINVDCx12_ASAP7_75t_R g191 ( 
.A(n_131),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_191),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_193),
.Y(n_267)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_194),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_159),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g277 ( 
.A(n_195),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_196),
.A2(n_212),
.B1(n_234),
.B2(n_123),
.Y(n_242)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_117),
.Y(n_197)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_119),
.B(n_38),
.Y(n_198)
);

INVx11_ASAP7_75t_SL g200 ( 
.A(n_176),
.Y(n_200)
);

INVx11_ASAP7_75t_L g286 ( 
.A(n_200),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_116),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_201),
.B(n_204),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_202),
.Y(n_264)
);

BUFx12f_ASAP7_75t_L g203 ( 
.A(n_133),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_203),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_141),
.B(n_47),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_205),
.A2(n_206),
.B1(n_221),
.B2(n_239),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_129),
.A2(n_75),
.B1(n_47),
.B2(n_106),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_157),
.B(n_49),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_207),
.B(n_215),
.Y(n_261)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_129),
.Y(n_208)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_208),
.Y(n_256)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_209),
.Y(n_257)
);

BUFx24_ASAP7_75t_L g210 ( 
.A(n_131),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_210),
.Y(n_288)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_135),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_211),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_114),
.A2(n_134),
.B1(n_83),
.B2(n_167),
.Y(n_212)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_154),
.Y(n_213)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_213),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_140),
.B(n_47),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_216),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_116),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_217),
.B(n_218),
.Y(n_266)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_133),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_111),
.Y(n_219)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_219),
.Y(n_280)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_165),
.Y(n_220)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_220),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_160),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_151),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_223),
.B(n_225),
.Y(n_282)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_118),
.Y(n_225)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_165),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_161),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_227),
.B(n_232),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_112),
.B(n_44),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_231),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_113),
.B(n_121),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_122),
.B(n_103),
.Y(n_232)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_161),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_233),
.B(n_238),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_149),
.A2(n_62),
.B1(n_2),
.B2(n_3),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_144),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_235),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_236),
.A2(n_120),
.B1(n_7),
.B2(n_8),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_139),
.B(n_1),
.C(n_5),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_237),
.B(n_9),
.Y(n_293)
);

INVx11_ASAP7_75t_L g239 ( 
.A(n_151),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g240 ( 
.A(n_142),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_240),
.A2(n_159),
.B1(n_143),
.B2(n_168),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_186),
.A2(n_118),
.B1(n_125),
.B2(n_145),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_241),
.A2(n_281),
.B1(n_284),
.B2(n_291),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_242),
.A2(n_279),
.B1(n_290),
.B2(n_289),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_238),
.A2(n_153),
.B(n_163),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_245),
.A2(n_210),
.B(n_239),
.Y(n_305)
);

AOI32xp33_ASAP7_75t_L g249 ( 
.A1(n_205),
.A2(n_158),
.A3(n_159),
.B1(n_127),
.B2(n_128),
.Y(n_249)
);

NOR2x1_ASAP7_75t_L g341 ( 
.A(n_249),
.B(n_289),
.Y(n_341)
);

NAND2xp33_ASAP7_75t_SL g252 ( 
.A(n_222),
.B(n_136),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_252),
.A2(n_292),
.B(n_258),
.Y(n_335)
);

AND2x2_ASAP7_75t_SL g253 ( 
.A(n_199),
.B(n_115),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_253),
.B(n_229),
.C(n_211),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_156),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_254),
.B(n_273),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_192),
.B(n_156),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_274),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_177),
.B(n_142),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_283),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_234),
.A2(n_125),
.B1(n_168),
.B2(n_126),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_180),
.B(n_6),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_222),
.A2(n_208),
.B1(n_224),
.B2(n_209),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_206),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_179),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_291)
);

NAND2xp33_ASAP7_75t_SL g292 ( 
.A(n_220),
.B(n_9),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_293),
.B(n_195),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_225),
.A2(n_233),
.B1(n_227),
.B2(n_188),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_294),
.A2(n_295),
.B1(n_288),
.B2(n_291),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_178),
.A2(n_9),
.B1(n_10),
.B2(n_190),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_213),
.B(n_10),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_10),
.Y(n_306)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_268),
.Y(n_299)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_299),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_286),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_300),
.B(n_302),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_250),
.B(n_226),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_264),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_303),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_304),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_305),
.A2(n_320),
.B(n_333),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_306),
.B(n_314),
.Y(n_361)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_254),
.Y(n_307)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_307),
.Y(n_363)
);

BUFx12f_ASAP7_75t_L g308 ( 
.A(n_287),
.Y(n_308)
);

INVx6_ASAP7_75t_L g352 ( 
.A(n_308),
.Y(n_352)
);

A2O1A1Ixp33_ASAP7_75t_SL g309 ( 
.A1(n_260),
.A2(n_210),
.B(n_200),
.C(n_230),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_309),
.A2(n_320),
.B(n_330),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_286),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_310),
.B(n_312),
.Y(n_368)
);

INVx8_ASAP7_75t_L g311 ( 
.A(n_244),
.Y(n_311)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_311),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_255),
.B(n_229),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_262),
.B(n_261),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_313),
.B(n_325),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_246),
.B(n_202),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_275),
.Y(n_315)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_315),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_316),
.B(n_333),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_246),
.B(n_221),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_317),
.B(n_324),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_277),
.Y(n_318)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_318),
.Y(n_381)
);

OAI21xp33_ASAP7_75t_SL g319 ( 
.A1(n_245),
.A2(n_240),
.B(n_203),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_319),
.A2(n_335),
.B(n_341),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_266),
.A2(n_203),
.B(n_218),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_275),
.Y(n_321)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_321),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_270),
.B(n_218),
.C(n_240),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_322),
.B(n_327),
.C(n_285),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_323),
.A2(n_329),
.B1(n_340),
.B2(n_345),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_272),
.B(n_283),
.Y(n_324)
);

AND2x6_ASAP7_75t_L g325 ( 
.A(n_258),
.B(n_252),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_273),
.Y(n_326)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_326),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_258),
.B(n_276),
.C(n_293),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_257),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_328),
.B(n_331),
.Y(n_386)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_268),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_296),
.B(n_276),
.Y(n_331)
);

INVx13_ASAP7_75t_L g332 ( 
.A(n_263),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_332),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_276),
.B(n_278),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_253),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_334),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_281),
.A2(n_279),
.B1(n_294),
.B2(n_282),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_336),
.A2(n_298),
.B1(n_326),
.B2(n_307),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_267),
.B(n_253),
.Y(n_337)
);

MAJx2_ASAP7_75t_L g373 ( 
.A(n_337),
.B(n_304),
.C(n_335),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_247),
.B(n_280),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_338),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_339),
.A2(n_342),
.B1(n_256),
.B2(n_285),
.Y(n_349)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_277),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_289),
.A2(n_256),
.B1(n_288),
.B2(n_257),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_280),
.B(n_269),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_343),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_265),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_344),
.Y(n_380)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_248),
.Y(n_345)
);

CKINVDCx14_ASAP7_75t_R g346 ( 
.A(n_292),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_346),
.A2(n_259),
.B(n_251),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_347),
.B(n_369),
.C(n_384),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g412 ( 
.A1(n_349),
.A2(n_356),
.B1(n_357),
.B2(n_379),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_353),
.A2(n_355),
.B(n_354),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_305),
.A2(n_259),
.B(n_243),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_355),
.A2(n_364),
.B(n_358),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_336),
.A2(n_243),
.B1(n_271),
.B2(n_244),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_339),
.A2(n_271),
.B1(n_264),
.B2(n_269),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_360),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_341),
.A2(n_248),
.B(n_251),
.Y(n_364)
);

OAI22x1_ASAP7_75t_L g366 ( 
.A1(n_325),
.A2(n_265),
.B1(n_277),
.B2(n_287),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_366),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_327),
.B(n_277),
.C(n_322),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_372),
.A2(n_383),
.B1(n_363),
.B2(n_365),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_373),
.B(n_376),
.Y(n_404)
);

XOR2x2_ASAP7_75t_L g376 ( 
.A(n_324),
.B(n_331),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_377),
.A2(n_360),
.B(n_364),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_297),
.A2(n_317),
.B1(n_314),
.B2(n_301),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_301),
.B(n_297),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_330),
.A2(n_309),
.B1(n_315),
.B2(n_321),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_385),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_332),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_387),
.B(n_318),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_342),
.B(n_306),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_389),
.B(n_384),
.C(n_347),
.Y(n_420)
);

XOR2x2_ASAP7_75t_L g390 ( 
.A(n_348),
.B(n_345),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_390),
.B(n_425),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_381),
.Y(n_392)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_392),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_365),
.B(n_328),
.Y(n_394)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_394),
.Y(n_436)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_362),
.Y(n_396)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_396),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_397),
.A2(n_423),
.B(n_377),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_348),
.B(n_308),
.Y(n_398)
);

XNOR2x1_ASAP7_75t_L g452 ( 
.A(n_398),
.B(n_420),
.Y(n_452)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_352),
.Y(n_399)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_399),
.Y(n_449)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_362),
.Y(n_400)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_400),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_367),
.B(n_308),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_401),
.B(n_402),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_368),
.B(n_340),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_371),
.B(n_303),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_403),
.B(n_416),
.Y(n_429)
);

INVx13_ASAP7_75t_L g405 ( 
.A(n_388),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_405),
.Y(n_431)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_375),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g448 ( 
.A(n_406),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_407),
.Y(n_437)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_375),
.Y(n_408)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_408),
.Y(n_451)
);

AND2x6_ASAP7_75t_L g409 ( 
.A(n_378),
.B(n_358),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_409),
.A2(n_418),
.B(n_353),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_411),
.A2(n_357),
.B1(n_374),
.B2(n_370),
.Y(n_445)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_382),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_413),
.B(n_408),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_361),
.B(n_311),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_414),
.B(n_424),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_351),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_415),
.B(n_419),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_388),
.B(n_309),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_376),
.B(n_309),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_417),
.B(n_422),
.Y(n_444)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_382),
.Y(n_419)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_363),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_421),
.B(n_372),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_380),
.B(n_389),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_361),
.B(n_379),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_369),
.B(n_350),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_383),
.B(n_381),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_426),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_350),
.B(n_386),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_427),
.B(n_349),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_430),
.A2(n_404),
.B(n_427),
.Y(n_471)
);

NAND2xp33_ASAP7_75t_SL g486 ( 
.A(n_433),
.B(n_459),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_411),
.B(n_386),
.Y(n_434)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_434),
.Y(n_467)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_440),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_415),
.B(n_370),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_441),
.B(n_446),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_442),
.B(n_453),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_445),
.A2(n_458),
.B1(n_413),
.B2(n_398),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_414),
.B(n_359),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_412),
.A2(n_366),
.B1(n_373),
.B2(n_359),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_447),
.A2(n_393),
.B1(n_395),
.B2(n_410),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_394),
.B(n_352),
.Y(n_450)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_450),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_421),
.B(n_424),
.Y(n_453)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_453),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_406),
.B(n_419),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_454),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_405),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_460),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_393),
.A2(n_423),
.B1(n_395),
.B2(n_410),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_418),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_452),
.B(n_391),
.C(n_425),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_462),
.B(n_469),
.C(n_484),
.Y(n_503)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_455),
.Y(n_463)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_463),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_464),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_459),
.A2(n_397),
.B(n_409),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_465),
.B(n_472),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_437),
.A2(n_400),
.B1(n_396),
.B2(n_399),
.Y(n_468)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_468),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_391),
.C(n_420),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_470),
.B(n_446),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_471),
.B(n_488),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_428),
.B(n_390),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_434),
.A2(n_404),
.B1(n_440),
.B2(n_445),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_473),
.B(n_475),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_458),
.A2(n_430),
.B(n_433),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_437),
.A2(n_428),
.B1(n_432),
.B2(n_438),
.Y(n_477)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_477),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_429),
.A2(n_438),
.B(n_441),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_478),
.B(n_480),
.Y(n_490)
);

AO22x1_ASAP7_75t_L g479 ( 
.A1(n_436),
.A2(n_448),
.B1(n_451),
.B2(n_429),
.Y(n_479)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_479),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_444),
.B(n_431),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_455),
.Y(n_481)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_481),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_482),
.B(n_435),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_443),
.B(n_442),
.C(n_447),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_444),
.B(n_431),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_485),
.B(n_460),
.Y(n_511)
);

FAx1_ASAP7_75t_SL g488 ( 
.A(n_435),
.B(n_436),
.CI(n_454),
.CON(n_488),
.SN(n_488)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_492),
.B(n_494),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_484),
.B(n_450),
.Y(n_494)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_474),
.Y(n_499)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_499),
.Y(n_515)
);

BUFx12f_ASAP7_75t_L g500 ( 
.A(n_466),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_500),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_SL g519 ( 
.A(n_502),
.B(n_464),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_473),
.B(n_456),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_505),
.B(n_482),
.Y(n_517)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_474),
.Y(n_506)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_506),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_469),
.B(n_448),
.C(n_451),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_507),
.B(n_510),
.Y(n_522)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_461),
.Y(n_508)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_508),
.Y(n_526)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_461),
.Y(n_509)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_509),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_462),
.B(n_448),
.C(n_451),
.Y(n_510)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_511),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_471),
.B(n_449),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_512),
.B(n_479),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_492),
.B(n_488),
.Y(n_514)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_514),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_517),
.B(n_510),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_497),
.A2(n_470),
.B1(n_483),
.B2(n_476),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_518),
.A2(n_491),
.B1(n_531),
.B2(n_500),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_519),
.B(n_520),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_494),
.B(n_475),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_493),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_521),
.B(n_523),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_507),
.B(n_478),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_524),
.B(n_502),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_490),
.B(n_489),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_525),
.B(n_479),
.Y(n_543)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_500),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_530),
.B(n_498),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_496),
.B(n_488),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_531),
.Y(n_535)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_532),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_533),
.B(n_537),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_SL g536 ( 
.A1(n_522),
.A2(n_503),
.B(n_504),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_536),
.A2(n_521),
.B(n_528),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_513),
.B(n_512),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g551 ( 
.A(n_539),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_513),
.B(n_465),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_540),
.B(n_541),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_519),
.B(n_501),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_520),
.B(n_503),
.C(n_486),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_542),
.B(n_543),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_518),
.A2(n_476),
.B1(n_467),
.B2(n_487),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_544),
.B(n_547),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_546),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_529),
.B(n_449),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_L g566 ( 
.A1(n_553),
.A2(n_515),
.B(n_526),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_542),
.A2(n_528),
.B(n_524),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g565 ( 
.A1(n_555),
.A2(n_557),
.B(n_544),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_L g557 ( 
.A1(n_539),
.A2(n_514),
.B(n_516),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_533),
.B(n_483),
.C(n_487),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_558),
.B(n_559),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_538),
.B(n_527),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_552),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_560),
.A2(n_562),
.B(n_563),
.Y(n_567)
);

MAJx2_ASAP7_75t_L g561 ( 
.A(n_548),
.B(n_534),
.C(n_545),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_561),
.B(n_565),
.C(n_566),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_549),
.B(n_535),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_556),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_SL g568 ( 
.A1(n_564),
.A2(n_562),
.B(n_554),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_568),
.B(n_569),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_SL g569 ( 
.A1(n_560),
.A2(n_551),
.B(n_558),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_567),
.B(n_550),
.C(n_551),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_SL g574 ( 
.A1(n_572),
.A2(n_550),
.B(n_495),
.Y(n_574)
);

AOI322xp5_ASAP7_75t_L g573 ( 
.A1(n_571),
.A2(n_570),
.A3(n_557),
.B1(n_495),
.B2(n_463),
.C1(n_540),
.C2(n_439),
.Y(n_573)
);

OAI21x1_ASAP7_75t_L g575 ( 
.A1(n_573),
.A2(n_574),
.B(n_481),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_575),
.A2(n_439),
.B(n_457),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_576),
.B(n_457),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_577),
.B(n_537),
.C(n_467),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_578),
.B(n_541),
.Y(n_579)
);


endmodule