module fake_jpeg_18750_n_161 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_161);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_161;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

INVx8_ASAP7_75t_SL g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx4f_ASAP7_75t_SL g55 ( 
.A(n_1),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_3),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_12),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx11_ASAP7_75t_SL g65 ( 
.A(n_14),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_6),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_81),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_84),
.Y(n_88)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_78),
.A2(n_72),
.B1(n_56),
.B2(n_74),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_89),
.B1(n_94),
.B2(n_53),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_79),
.A2(n_48),
.B1(n_65),
.B2(n_57),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_61),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_93),
.B(n_64),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_71),
.B1(n_73),
.B2(n_75),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_92),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_47),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_87),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_55),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_2),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_59),
.Y(n_102)
);

FAx1_ASAP7_75t_SL g122 ( 
.A(n_102),
.B(n_53),
.CI(n_54),
.CON(n_122),
.SN(n_122)
);

AND2x4_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_73),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_108),
.B(n_96),
.Y(n_111)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_104),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_107),
.B1(n_0),
.B2(n_2),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_69),
.B1(n_75),
.B2(n_51),
.Y(n_107)
);

NAND2xp33_ASAP7_75t_SL g108 ( 
.A(n_86),
.B(n_62),
.Y(n_108)
);

AOI21xp33_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_119),
.B(n_122),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_63),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_113),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_98),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_114),
.A2(n_120),
.B(n_125),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_123),
.B1(n_4),
.B2(n_5),
.Y(n_127)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

NOR2xp67_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_0),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_66),
.B(n_50),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_67),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_122),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_52),
.B1(n_70),
.B2(n_32),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_131),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_4),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_115),
.Y(n_140)
);

AOI221xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_34),
.B1(n_45),
.B2(n_16),
.C(n_19),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_134),
.B(n_36),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_136),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_110),
.A2(n_35),
.B1(n_42),
.B2(n_20),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_137),
.A2(n_30),
.B1(n_40),
.B2(n_26),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_139),
.B(n_142),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

INVx3_ASAP7_75t_SL g141 ( 
.A(n_130),
.Y(n_141)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_147),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_140),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_144),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_138),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_147),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_154),
.B(n_143),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_155),
.A2(n_126),
.B(n_129),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_146),
.C(n_145),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_148),
.C(n_128),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_148),
.C(n_37),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_159),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_27),
.B(n_29),
.Y(n_161)
);


endmodule