module fake_jpeg_19240_n_38 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_38);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_38;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_0),
.Y(n_22)
);

O2A1O1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_23),
.B(n_25),
.C(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_0),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_20),
.B1(n_4),
.B2(n_5),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_1),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_26),
.B(n_28),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_27),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_25),
.A2(n_3),
.B1(n_8),
.B2(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_10),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_34),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_27),
.Y(n_34)
);

FAx1_ASAP7_75t_SL g36 ( 
.A(n_35),
.B(n_32),
.CI(n_12),
.CON(n_36),
.SN(n_36)
);

OAI211xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_11),
.B(n_13),
.C(n_15),
.Y(n_37)
);

BUFx24_ASAP7_75t_SL g38 ( 
.A(n_37),
.Y(n_38)
);


endmodule