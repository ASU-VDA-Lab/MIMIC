module fake_jpeg_26666_n_44 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_31;
wire n_17;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_0),
.B(n_4),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx6_ASAP7_75t_SL g10 ( 
.A(n_3),
.Y(n_10)
);

INVx11_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g13 ( 
.A(n_5),
.B(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

AND2x2_ASAP7_75t_SL g16 ( 
.A(n_1),
.B(n_2),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_22),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_19)
);

AOI21xp33_ASAP7_75t_L g29 ( 
.A1(n_19),
.A2(n_23),
.B(n_24),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx10_ASAP7_75t_R g30 ( 
.A(n_20),
.Y(n_30)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_16),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_26),
.C(n_9),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_29),
.C(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_16),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_37),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_13),
.B(n_18),
.Y(n_37)
);

INVxp33_ASAP7_75t_SL g39 ( 
.A(n_37),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_39),
.A2(n_25),
.B1(n_28),
.B2(n_21),
.Y(n_41)
);

AOI322xp5_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_13),
.A3(n_30),
.B1(n_31),
.B2(n_17),
.C1(n_16),
.C2(n_32),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_40),
.A2(n_41),
.B1(n_17),
.B2(n_13),
.Y(n_42)
);

AOI322xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_41),
.A3(n_17),
.B1(n_15),
.B2(n_9),
.C1(n_20),
.C2(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_15),
.Y(n_44)
);


endmodule