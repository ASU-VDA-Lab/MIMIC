module fake_jpeg_664_n_416 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_416);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_416;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_1),
.B(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_47),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_48),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g101 ( 
.A(n_49),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_50),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_67),
.Y(n_89)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_8),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_57),
.B(n_65),
.Y(n_108)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_8),
.C(n_13),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_42),
.C(n_30),
.Y(n_97)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_21),
.B(n_7),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_75),
.Y(n_110)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_80),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_77),
.Y(n_98)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_81),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_82),
.B(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_31),
.B(n_7),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_87),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_86),
.Y(n_125)
);

NAND2xp33_ASAP7_75t_SL g87 ( 
.A(n_15),
.B(n_6),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_51),
.A2(n_43),
.B1(n_24),
.B2(n_34),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_90),
.A2(n_94),
.B1(n_138),
.B2(n_125),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_60),
.A2(n_63),
.B1(n_41),
.B2(n_34),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_93),
.A2(n_102),
.B1(n_128),
.B2(n_135),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_45),
.A2(n_18),
.B1(n_42),
.B2(n_38),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_97),
.B(n_5),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_68),
.A2(n_41),
.B1(n_34),
.B2(n_15),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_16),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_106),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_16),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_56),
.B(n_24),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_19),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_38),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_117),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_29),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_58),
.A2(n_41),
.B1(n_15),
.B2(n_43),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_62),
.A2(n_48),
.B1(n_50),
.B2(n_46),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_130),
.A2(n_132),
.B1(n_0),
.B2(n_1),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_44),
.A2(n_36),
.B1(n_30),
.B2(n_29),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_86),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_125),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_66),
.A2(n_36),
.B1(n_26),
.B2(n_18),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_64),
.A2(n_26),
.B1(n_37),
.B2(n_19),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_19),
.B1(n_37),
.B2(n_75),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_139),
.A2(n_120),
.B1(n_136),
.B2(n_137),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_141),
.B(n_164),
.Y(n_191)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_142),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_101),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_143),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_37),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_144),
.B(n_154),
.Y(n_193)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_145),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_77),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_146),
.B(n_151),
.C(n_173),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_108),
.B(n_72),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_147),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_148),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_103),
.A2(n_71),
.B1(n_55),
.B2(n_49),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_150),
.A2(n_156),
.B1(n_158),
.B2(n_163),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_97),
.B(n_84),
.C(n_53),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_152),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_153),
.A2(n_177),
.B1(n_180),
.B2(n_156),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_89),
.B(n_0),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_99),
.B(n_0),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_155),
.B(n_161),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_90),
.A2(n_49),
.B1(n_1),
.B2(n_2),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_95),
.A2(n_47),
.B(n_9),
.C(n_10),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_158),
.B(n_163),
.Y(n_201)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_88),
.B(n_0),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_162),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_6),
.B(n_12),
.C(n_11),
.Y(n_163)
);

AO22x2_ASAP7_75t_SL g165 ( 
.A1(n_110),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_126),
.B(n_127),
.C(n_124),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_111),
.A2(n_5),
.B1(n_6),
.B2(n_10),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_166),
.A2(n_168),
.B1(n_178),
.B2(n_96),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_88),
.B(n_91),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_167),
.B(n_170),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_111),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_110),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_119),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_110),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_172),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_91),
.B(n_11),
.C(n_14),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_2),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_182),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_131),
.B(n_2),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_176),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_98),
.A2(n_3),
.B1(n_122),
.B2(n_137),
.Y(n_177)
);

INVx11_ASAP7_75t_L g178 ( 
.A(n_96),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_131),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_179),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_107),
.A2(n_3),
.B1(n_124),
.B2(n_109),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_104),
.Y(n_181)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_104),
.B(n_98),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_113),
.B(n_118),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_127),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_113),
.B(n_118),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_144),
.Y(n_198)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_100),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

INVx4_ASAP7_75t_SL g248 ( 
.A(n_187),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_189),
.A2(n_221),
.B1(n_224),
.B2(n_173),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_194),
.Y(n_233)
);

AND2x2_ASAP7_75t_SL g195 ( 
.A(n_141),
.B(n_100),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_195),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_197),
.B(n_198),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_176),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_203),
.A2(n_210),
.B1(n_211),
.B2(n_213),
.Y(n_227)
);

AOI32xp33_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_119),
.A3(n_126),
.B1(n_133),
.B2(n_116),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_183),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_175),
.A2(n_107),
.B1(n_109),
.B2(n_136),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_164),
.A2(n_120),
.B1(n_116),
.B2(n_121),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_147),
.A2(n_121),
.B1(n_133),
.B2(n_101),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_147),
.A2(n_160),
.B1(n_170),
.B2(n_172),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_216),
.A2(n_171),
.B1(n_151),
.B2(n_150),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_182),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_217),
.B(n_159),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_153),
.A2(n_96),
.B1(n_146),
.B2(n_171),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_167),
.B(n_176),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_223),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_221),
.A2(n_189),
.B1(n_217),
.B2(n_191),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_226),
.A2(n_231),
.B1(n_242),
.B2(n_246),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_228),
.B(n_245),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_229),
.B(n_202),
.Y(n_281)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_230),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_191),
.A2(n_161),
.B1(n_140),
.B2(n_149),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_213),
.A2(n_143),
.B1(n_169),
.B2(n_180),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_232),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_234),
.A2(n_238),
.B(n_249),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_206),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_235),
.B(n_254),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_208),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_236),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_216),
.A2(n_165),
.B1(n_174),
.B2(n_155),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_237),
.A2(n_204),
.B1(n_192),
.B2(n_209),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_201),
.A2(n_165),
.B(n_154),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_239),
.Y(n_283)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_240),
.Y(n_285)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_200),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_241),
.Y(n_269)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_186),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_244),
.Y(n_279)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_191),
.A2(n_165),
.B1(n_142),
.B2(n_152),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_222),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_252),
.Y(n_277)
);

A2O1A1O1Ixp25_ASAP7_75t_L g249 ( 
.A1(n_214),
.A2(n_181),
.B(n_185),
.C(n_145),
.D(n_157),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_148),
.C(n_152),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_229),
.C(n_226),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_219),
.B(n_178),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_253),
.B(n_260),
.Y(n_263)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_207),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_207),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_258),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_215),
.B(n_222),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_223),
.Y(n_284)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_209),
.A2(n_224),
.B1(n_195),
.B2(n_204),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_259),
.A2(n_197),
.B1(n_220),
.B2(n_192),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_219),
.B(n_193),
.Y(n_260)
);

AOI21xp33_ASAP7_75t_L g261 ( 
.A1(n_228),
.A2(n_201),
.B(n_197),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_261),
.A2(n_287),
.B(n_238),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_262),
.A2(n_265),
.B1(n_267),
.B2(n_286),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_237),
.A2(n_195),
.B1(n_212),
.B2(n_198),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_248),
.A2(n_195),
.B1(n_212),
.B2(n_198),
.Y(n_267)
);

AO21x1_ASAP7_75t_L g300 ( 
.A1(n_270),
.A2(n_289),
.B(n_227),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_250),
.C(n_256),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_199),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_278),
.B(n_284),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_236),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_280),
.B(n_290),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_231),
.Y(n_297)
);

OAI32xp33_ASAP7_75t_L g282 ( 
.A1(n_256),
.A2(n_223),
.A3(n_193),
.B1(n_187),
.B2(n_205),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_282),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_248),
.A2(n_220),
.B1(n_187),
.B2(n_211),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_259),
.A2(n_196),
.B(n_188),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_247),
.B(n_210),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_288),
.B(n_258),
.Y(n_306)
);

AND2x6_ASAP7_75t_L g289 ( 
.A(n_249),
.B(n_196),
.Y(n_289)
);

OA22x2_ASAP7_75t_L g290 ( 
.A1(n_248),
.A2(n_203),
.B1(n_225),
.B2(n_208),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_233),
.A2(n_190),
.B(n_199),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_291),
.A2(n_233),
.B(n_246),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_292),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_293),
.B(n_298),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_287),
.A2(n_251),
.B(n_243),
.Y(n_294)
);

NOR2xp67_ASAP7_75t_SL g332 ( 
.A(n_294),
.B(n_275),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_273),
.A2(n_227),
.B1(n_251),
.B2(n_257),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_296),
.B(n_301),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_297),
.B(n_303),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_245),
.C(n_244),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_275),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_299),
.B(n_271),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_300),
.B(n_306),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_291),
.A2(n_240),
.B(n_241),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_302),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_230),
.C(n_239),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_277),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_304),
.B(n_305),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_277),
.B(n_255),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_270),
.B(n_225),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_312),
.Y(n_322)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_274),
.Y(n_308)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_308),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_265),
.A2(n_273),
.B1(n_262),
.B2(n_266),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_309),
.A2(n_314),
.B1(n_315),
.B2(n_290),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_266),
.B(n_264),
.C(n_263),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_266),
.A2(n_288),
.B1(n_268),
.B2(n_282),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_313),
.A2(n_290),
.B1(n_271),
.B2(n_283),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_286),
.A2(n_267),
.B1(n_263),
.B2(n_289),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_289),
.A2(n_274),
.B1(n_269),
.B2(n_279),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_264),
.A2(n_290),
.B1(n_269),
.B2(n_279),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_290),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_319),
.A2(n_321),
.B1(n_338),
.B2(n_329),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_321),
.A2(n_340),
.B1(n_310),
.B2(n_302),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_276),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_326),
.B(n_303),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_310),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_335),
.Y(n_355)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_329),
.Y(n_341)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_308),
.Y(n_330)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_330),
.Y(n_350)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_299),
.Y(n_331)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_331),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_332),
.A2(n_294),
.B(n_292),
.Y(n_343)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_311),
.Y(n_333)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_333),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_305),
.B(n_311),
.Y(n_334)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_334),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_310),
.Y(n_335)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_336),
.Y(n_345)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_317),
.Y(n_338)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_338),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_309),
.A2(n_283),
.B1(n_285),
.B2(n_280),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_343),
.A2(n_339),
.B(n_332),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_344),
.A2(n_349),
.B1(n_358),
.B2(n_315),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_328),
.B(n_293),
.C(n_298),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_346),
.B(n_357),
.C(n_359),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_334),
.Y(n_347)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_347),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_351),
.B(n_352),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_328),
.B(n_296),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_324),
.B(n_297),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_354),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_324),
.B(n_307),
.C(n_304),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_319),
.A2(n_316),
.B1(n_313),
.B2(n_295),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_322),
.B(n_295),
.C(n_316),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_346),
.B(n_337),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_360),
.B(n_362),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_357),
.B(n_337),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_365),
.A2(n_301),
.B(n_348),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_366),
.B(n_369),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_359),
.B(n_314),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_367),
.B(n_370),
.Y(n_384)
);

HAxp5_ASAP7_75t_SL g368 ( 
.A(n_343),
.B(n_320),
.CON(n_368),
.SN(n_368)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_368),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_342),
.B(n_300),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_358),
.A2(n_320),
.B1(n_318),
.B2(n_333),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_341),
.A2(n_340),
.B1(n_325),
.B2(n_318),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_371),
.A2(n_374),
.B1(n_349),
.B2(n_355),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_342),
.B(n_300),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_345),
.C(n_344),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_341),
.A2(n_325),
.B1(n_335),
.B2(n_327),
.Y(n_374)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_375),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_365),
.A2(n_355),
.B(n_348),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_377),
.B(n_378),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_364),
.B(n_345),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_379),
.B(n_380),
.Y(n_387)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_361),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_374),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_383),
.Y(n_393)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_371),
.Y(n_383)
);

NOR2xp67_ASAP7_75t_SL g392 ( 
.A(n_386),
.B(n_367),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_380),
.B(n_323),
.Y(n_388)
);

OAI21x1_ASAP7_75t_L g402 ( 
.A1(n_388),
.A2(n_390),
.B(n_392),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_376),
.B(n_363),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_389),
.B(n_394),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_377),
.B(n_330),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_376),
.B(n_373),
.C(n_360),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_384),
.A2(n_370),
.B1(n_366),
.B2(n_323),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_396),
.B(n_331),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_397),
.B(n_400),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_387),
.B(n_386),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_399),
.B(n_403),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_391),
.B(n_373),
.C(n_362),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_395),
.A2(n_381),
.B(n_379),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_401),
.A2(n_385),
.B(n_353),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_393),
.B(n_372),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_399),
.A2(n_390),
.B1(n_356),
.B2(n_388),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_404),
.A2(n_406),
.B1(n_407),
.B2(n_350),
.Y(n_411)
);

AOI211xp5_ASAP7_75t_SL g406 ( 
.A1(n_402),
.A2(n_368),
.B(n_369),
.C(n_385),
.Y(n_406)
);

XNOR2x2_ASAP7_75t_SL g409 ( 
.A(n_405),
.B(n_398),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_409),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_408),
.A2(n_400),
.B(n_336),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_410),
.A2(n_411),
.B(n_406),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_413),
.B(n_285),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_414),
.B(n_412),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_415),
.B(n_278),
.Y(n_416)
);


endmodule