module fake_ariane_443_n_105 (n_8, n_7, n_1, n_6, n_13, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_16, n_5, n_12, n_15, n_10, n_105);

input n_8;
input n_7;
input n_1;
input n_6;
input n_13;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_16;
input n_5;
input n_12;
input n_15;
input n_10;

output n_105;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_19;
wire n_40;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_72;
wire n_44;
wire n_30;
wire n_82;
wire n_42;
wire n_31;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_102;
wire n_22;
wire n_81;
wire n_87;
wire n_43;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_35;
wire n_54;
wire n_25;

CKINVDCx5p33_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVxp67_ASAP7_75t_SL g26 ( 
.A(n_1),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVxp67_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NAND2xp33_ASAP7_75t_SL g45 ( 
.A(n_19),
.B(n_3),
.Y(n_45)
);

CKINVDCx6p67_ASAP7_75t_R g46 ( 
.A(n_28),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_26),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

AND2x4_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_21),
.Y(n_51)
);

OAI221xp5_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_26),
.B1(n_27),
.B2(n_34),
.C(n_21),
.Y(n_52)
);

AO22x2_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_53)
);

AND2x4_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_36),
.Y(n_54)
);

AO22x2_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_46),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_52),
.A2(n_33),
.B1(n_24),
.B2(n_47),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_48),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_31),
.B(n_36),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_60),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_53),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_54),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

AND2x4_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_54),
.Y(n_70)
);

AO21x2_ASAP7_75t_L g71 ( 
.A1(n_67),
.A2(n_61),
.B(n_39),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_46),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_53),
.B1(n_55),
.B2(n_58),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_69),
.A2(n_68),
.B(n_66),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_73),
.B(n_72),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_70),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_78),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_55),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_63),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_81),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_83),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_82),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_34),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_90),
.B(n_84),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_25),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_25),
.C(n_44),
.Y(n_97)
);

OAI221xp5_ASAP7_75t_L g98 ( 
.A1(n_92),
.A2(n_45),
.B1(n_44),
.B2(n_43),
.C(n_50),
.Y(n_98)
);

NOR3xp33_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_43),
.C(n_51),
.Y(n_99)
);

AOI221xp5_ASAP7_75t_L g100 ( 
.A1(n_98),
.A2(n_55),
.B1(n_53),
.B2(n_93),
.C(n_95),
.Y(n_100)
);

AOI222xp33_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_96),
.B1(n_97),
.B2(n_55),
.C1(n_51),
.C2(n_99),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_75),
.B1(n_66),
.B2(n_65),
.Y(n_102)
);

OAI211xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_5),
.B(n_7),
.C(n_9),
.Y(n_103)
);

OAI222xp33_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_9),
.B1(n_10),
.B2(n_71),
.C1(n_14),
.C2(n_12),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_71),
.B1(n_16),
.B2(n_18),
.Y(n_105)
);


endmodule