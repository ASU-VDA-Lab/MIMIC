module fake_jpeg_3010_n_222 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_222);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_222;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_25),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_21),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_38),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_26),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_10),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx8_ASAP7_75t_SL g75 ( 
.A(n_13),
.Y(n_75)
);

BUFx16f_ASAP7_75t_L g76 ( 
.A(n_8),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_82),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_84),
.Y(n_91)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_68),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_90),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_83),
.B(n_77),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_88),
.B(n_66),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_81),
.A2(n_57),
.B1(n_53),
.B2(n_75),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_63),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_84),
.A2(n_57),
.B1(n_53),
.B2(n_70),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_93),
.A2(n_95),
.B1(n_96),
.B2(n_56),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_69),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_94),
.B(n_54),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_70),
.B1(n_69),
.B2(n_64),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_79),
.A2(n_59),
.B1(n_73),
.B2(n_55),
.Y(n_96)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_56),
.B(n_61),
.C(n_65),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_100),
.B(n_103),
.Y(n_127)
);

OA22x2_ASAP7_75t_SL g101 ( 
.A1(n_88),
.A2(n_74),
.B1(n_71),
.B2(n_62),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_101),
.Y(n_123)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_91),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_60),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_115),
.Y(n_119)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_111),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_68),
.B1(n_72),
.B2(n_60),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_109),
.A2(n_74),
.B1(n_71),
.B2(n_2),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_97),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_50),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_51),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_66),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_121),
.B(n_122),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_63),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_107),
.C(n_100),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_117),
.C(n_49),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_61),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_4),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_114),
.A2(n_98),
.B1(n_92),
.B2(n_72),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_120),
.B1(n_131),
.B2(n_123),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_92),
.B(n_62),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_7),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_32),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_133),
.A2(n_136),
.B1(n_5),
.B2(n_6),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_0),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_135),
.B(n_137),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_101),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_3),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_140),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_146),
.C(n_140),
.Y(n_171)
);

NOR2x1_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_4),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_144),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_147),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_46),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_120),
.A2(n_45),
.B1(n_43),
.B2(n_41),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_126),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_149),
.Y(n_172)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_40),
.B(n_33),
.Y(n_150)
);

NAND3xp33_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_27),
.C(n_24),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_134),
.A2(n_31),
.B(n_29),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_151),
.A2(n_23),
.B(n_9),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_153),
.B(n_164),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_163),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_5),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_156),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_158),
.Y(n_178)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_161),
.Y(n_183)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_124),
.B(n_7),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_171),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_142),
.A2(n_130),
.B(n_136),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_166),
.A2(n_174),
.B(n_175),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_16),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_158),
.A2(n_133),
.B1(n_140),
.B2(n_10),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_151),
.B1(n_146),
.B2(n_159),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_143),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_11),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_181),
.C(n_18),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_156),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_182),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_12),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

XNOR2x1_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_153),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_193),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_186),
.A2(n_191),
.B1(n_174),
.B2(n_187),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_167),
.A2(n_14),
.B(n_15),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_192),
.Y(n_201)
);

OAI321xp33_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_14),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.C(n_18),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_17),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_194),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_181),
.C(n_165),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_182),
.B(n_19),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_177),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_198),
.A2(n_170),
.B1(n_178),
.B2(n_169),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_203),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_171),
.C(n_180),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_195),
.C(n_176),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_202),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_185),
.B(n_172),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_190),
.Y(n_204)
);

INVx11_ASAP7_75t_L g206 ( 
.A(n_204),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_207),
.A2(n_209),
.B1(n_211),
.B2(n_204),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_188),
.C(n_193),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_213),
.Y(n_215)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_206),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_206),
.A2(n_197),
.B1(n_208),
.B2(n_209),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_214),
.A2(n_197),
.B1(n_210),
.B2(n_201),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_216),
.B(n_214),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_217),
.B(n_216),
.Y(n_218)
);

A2O1A1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_218),
.A2(n_215),
.B(n_207),
.C(n_173),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_219),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_220),
.A2(n_210),
.B1(n_20),
.B2(n_22),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_19),
.Y(n_222)
);


endmodule