module fake_jpeg_8656_n_118 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_118);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_118;

wire n_117;
wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_22),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx5_ASAP7_75t_SL g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_14),
.B1(n_17),
.B2(n_15),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_31),
.A2(n_35),
.B1(n_17),
.B2(n_11),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_22),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_22),
.A2(n_17),
.B1(n_14),
.B2(n_18),
.Y(n_35)
);

NAND3xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_0),
.C(n_1),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_16),
.B(n_11),
.C(n_19),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_26),
.B(n_23),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_20),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_40),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_18),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_47),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_20),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_44),
.Y(n_58)
);

INVxp67_ASAP7_75t_SL g61 ( 
.A(n_43),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_15),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_14),
.B1(n_16),
.B2(n_10),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_19),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_48),
.Y(n_59)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_49),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_27),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_18),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_56),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_49),
.B1(n_41),
.B2(n_45),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_10),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_60),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_12),
.B(n_22),
.C(n_3),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_45),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_60),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_63),
.B(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2x1p5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_45),
.Y(n_67)
);

AOI21x1_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_63),
.B(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_70),
.B(n_54),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_52),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_74),
.B(n_78),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_67),
.C(n_48),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_81),
.A2(n_67),
.B(n_69),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_39),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_91),
.C(n_1),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_81),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_88),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_76),
.Y(n_89)
);

BUFx24_ASAP7_75t_SL g92 ( 
.A(n_89),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_47),
.B1(n_32),
.B2(n_24),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_90),
.A2(n_77),
.B1(n_82),
.B2(n_80),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_36),
.C(n_34),
.Y(n_91)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

OA21x2_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_86),
.B(n_8),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_88),
.A2(n_6),
.B1(n_8),
.B2(n_7),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_97),
.A2(n_7),
.B1(n_5),
.B2(n_87),
.Y(n_102)
);

OAI31xp33_ASAP7_75t_L g100 ( 
.A1(n_94),
.A2(n_84),
.A3(n_83),
.B(n_85),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_100),
.A2(n_101),
.B(n_92),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_2),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_95),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_108),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_105),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_99),
.B(n_96),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_107),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_98),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_110),
.A2(n_109),
.B(n_111),
.Y(n_112)
);

AOI211xp5_ASAP7_75t_L g115 ( 
.A1(n_112),
.A2(n_113),
.B(n_4),
.C(n_36),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_111),
.B(n_107),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_3),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_114),
.Y(n_116)
);

AO21x1_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_115),
.B(n_4),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_24),
.Y(n_118)
);


endmodule