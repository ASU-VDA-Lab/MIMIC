module fake_jpeg_1052_n_159 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_159);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_48),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_1),
.Y(n_67)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_62),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_46),
.Y(n_71)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVxp67_ASAP7_75t_SL g91 ( 
.A(n_64),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_49),
.B1(n_51),
.B2(n_46),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_51),
.B1(n_53),
.B2(n_45),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_67),
.B(n_69),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_56),
.Y(n_69)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_56),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_75),
.B(n_52),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_79),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_66),
.A2(n_49),
.B1(n_55),
.B2(n_45),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_86),
.B1(n_6),
.B2(n_8),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_55),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_42),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_9),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_42),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_43),
.B1(n_41),
.B2(n_53),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_2),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_88),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_17),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_50),
.B(n_53),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_2),
.B(n_3),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_89),
.A2(n_65),
.B1(n_68),
.B2(n_64),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_98),
.B1(n_100),
.B2(n_105),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_85),
.A2(n_74),
.B1(n_68),
.B2(n_4),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_99),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_82),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_106),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_74),
.C(n_16),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_11),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_81),
.A2(n_15),
.B1(n_38),
.B2(n_37),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_102),
.B(n_14),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_10),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_26),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_113),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_88),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_11),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_122),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_101),
.A2(n_91),
.B1(n_12),
.B2(n_13),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_112),
.B1(n_116),
.B2(n_118),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_40),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_118),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_119),
.A2(n_33),
.B1(n_36),
.B2(n_117),
.Y(n_135)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_93),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_125),
.Y(n_134)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_98),
.A2(n_19),
.B(n_20),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_109),
.A2(n_22),
.B(n_25),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_133),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_29),
.B(n_32),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_135),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_115),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_137),
.B(n_112),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_139),
.A2(n_110),
.B1(n_127),
.B2(n_138),
.Y(n_142)
);

OA21x2_ASAP7_75t_SL g148 ( 
.A1(n_141),
.A2(n_134),
.B(n_136),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_133),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_139),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_144),
.C(n_146),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_134),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_148),
.Y(n_151)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_147),
.C(n_149),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_152),
.A2(n_150),
.B(n_140),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

NOR2x1p5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_141),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_145),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_131),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_132),
.Y(n_159)
);


endmodule