module fake_jpeg_23305_n_272 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_272);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_20),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_32),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_25),
.B(n_12),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_1),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_16),
.Y(n_43)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_44),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_43),
.B(n_37),
.Y(n_67)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_24),
.B1(n_18),
.B2(n_27),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_48),
.B1(n_30),
.B2(n_35),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_32),
.A2(n_24),
.B1(n_18),
.B2(n_14),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_32),
.A2(n_24),
.B1(n_18),
.B2(n_22),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_51),
.B1(n_21),
.B2(n_23),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_32),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_53),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_31),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_SL g78 ( 
.A(n_55),
.B(n_72),
.C(n_42),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_36),
.B(n_35),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_70),
.B(n_73),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_58),
.A2(n_19),
.B1(n_46),
.B2(n_39),
.Y(n_88)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_62),
.Y(n_90)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_31),
.B1(n_33),
.B2(n_29),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_42),
.B1(n_31),
.B2(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_34),
.Y(n_66)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_49),
.B(n_25),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_40),
.B(n_30),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_19),
.B1(n_17),
.B2(n_13),
.Y(n_89)
);

NAND2x1_ASAP7_75t_SL g72 ( 
.A(n_42),
.B(n_31),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_40),
.B(n_36),
.Y(n_73)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_81),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_82),
.B(n_93),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_79),
.A2(n_88),
.B1(n_69),
.B2(n_60),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_45),
.B1(n_48),
.B2(n_36),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_85),
.B1(n_87),
.B2(n_89),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_57),
.A2(n_26),
.B(n_53),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_53),
.C(n_47),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_86),
.C(n_71),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_59),
.A2(n_39),
.B1(n_41),
.B2(n_46),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_33),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_58),
.A2(n_39),
.B1(n_41),
.B2(n_46),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_55),
.A2(n_33),
.B(n_29),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_64),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_55),
.B(n_63),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_96),
.A2(n_109),
.B(n_110),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_104),
.C(n_79),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_77),
.B(n_91),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_100),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_77),
.B(n_62),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_88),
.B1(n_69),
.B2(n_72),
.Y(n_123)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_102),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_103),
.B(n_105),
.Y(n_115)
);

MAJx2_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_55),
.C(n_64),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_90),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_75),
.A2(n_58),
.B(n_72),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_72),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_92),
.B(n_67),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_111),
.B(n_12),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_91),
.B(n_66),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_75),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_126),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_94),
.B(n_74),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_119),
.A2(n_135),
.B(n_33),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_109),
.A2(n_89),
.B1(n_82),
.B2(n_74),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_120),
.A2(n_122),
.B1(n_110),
.B2(n_111),
.Y(n_143)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_134),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_114),
.A2(n_80),
.B1(n_87),
.B2(n_79),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_124),
.B1(n_129),
.B2(n_61),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_79),
.B1(n_92),
.B2(n_61),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_79),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_104),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_130),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_133),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_68),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_69),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_99),
.A2(n_61),
.B(n_56),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_136),
.B(n_11),
.Y(n_144)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_140),
.Y(n_161)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_116),
.B(n_106),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_145),
.B(n_151),
.Y(n_163)
);

OAI32xp33_ASAP7_75t_L g142 ( 
.A1(n_120),
.A2(n_105),
.A3(n_113),
.B1(n_110),
.B2(n_112),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_144),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_143),
.A2(n_148),
.B1(n_153),
.B2(n_118),
.Y(n_165)
);

OA21x2_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_132),
.B(n_124),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_149),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_117),
.B(n_102),
.Y(n_147)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_122),
.A2(n_128),
.B1(n_115),
.B2(n_126),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_154),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_133),
.B(n_97),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_97),
.B1(n_60),
.B2(n_61),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_61),
.Y(n_156)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_54),
.B1(n_52),
.B2(n_17),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_127),
.B(n_11),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_144),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_60),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_29),
.Y(n_169)
);

BUFx4f_ASAP7_75t_SL g162 ( 
.A(n_154),
.Y(n_162)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_165),
.B(n_138),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_143),
.A2(n_54),
.B1(n_52),
.B2(n_29),
.Y(n_167)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_177),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_54),
.B1(n_52),
.B2(n_17),
.Y(n_170)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_15),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_176),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_152),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_173),
.A2(n_137),
.B1(n_140),
.B2(n_146),
.Y(n_187)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_15),
.C(n_20),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_15),
.C(n_20),
.Y(n_177)
);

INVxp33_ASAP7_75t_SL g178 ( 
.A(n_145),
.Y(n_178)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_20),
.C(n_13),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_153),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_182),
.Y(n_186)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

XNOR2x1_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_148),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_184),
.B(n_167),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_185),
.A2(n_187),
.B(n_177),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_SL g190 ( 
.A1(n_163),
.A2(n_145),
.B(n_160),
.C(n_147),
.Y(n_190)
);

A2O1A1Ixp33_ASAP7_75t_SL g208 ( 
.A1(n_190),
.A2(n_180),
.B(n_176),
.C(n_172),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_162),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_191),
.A2(n_193),
.B(n_195),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_192),
.Y(n_202)
);

NOR3xp33_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_142),
.C(n_145),
.Y(n_193)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_152),
.B(n_138),
.C(n_141),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_169),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_158),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_171),
.Y(n_207)
);

NAND3xp33_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_168),
.C(n_161),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_203),
.A2(n_9),
.B(n_4),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_204),
.B(n_205),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_199),
.A2(n_179),
.B1(n_174),
.B2(n_171),
.Y(n_206)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_208),
.A2(n_212),
.B(n_190),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_198),
.B(n_138),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_10),
.C(n_9),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_187),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_213),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_1),
.C(n_2),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_197),
.C(n_183),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_194),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_215),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_195),
.B(n_11),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_217),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_186),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_196),
.B(n_9),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_10),
.Y(n_223)
);

AOI21xp33_ASAP7_75t_L g219 ( 
.A1(n_203),
.A2(n_193),
.B(n_190),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_219),
.A2(n_224),
.B(n_227),
.Y(n_234)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

BUFx24_ASAP7_75t_SL g225 ( 
.A(n_211),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_208),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_228),
.A2(n_215),
.B(n_208),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_2),
.C(n_3),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_214),
.C(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_232),
.Y(n_237)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_235),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_230),
.B(n_209),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_220),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_205),
.C(n_202),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_6),
.C(n_7),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_208),
.B1(n_4),
.B2(n_5),
.Y(n_240)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_242),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_3),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_5),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_244),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_226),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_247),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_221),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_251),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_244),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_237),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_254),
.A2(n_253),
.B(n_245),
.Y(n_260)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_256),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_249),
.B(n_233),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_259),
.Y(n_263)
);

NOR2x1_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_238),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_L g265 ( 
.A1(n_258),
.A2(n_6),
.B(n_7),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_6),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_261),
.A2(n_254),
.B(n_7),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_262),
.A2(n_264),
.B(n_265),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_266),
.A2(n_255),
.B(n_258),
.Y(n_267)
);

INVxp33_ASAP7_75t_L g269 ( 
.A(n_267),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_269),
.A2(n_263),
.B(n_268),
.Y(n_270)
);

AO21x1_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_6),
.B(n_7),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_8),
.Y(n_272)
);


endmodule