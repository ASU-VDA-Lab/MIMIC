module fake_jpeg_11104_n_439 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_439);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_439;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_50),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_16),
.B(n_25),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_75),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_54),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_55),
.Y(n_140)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_89),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_60),
.Y(n_117)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_16),
.B(n_7),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_64),
.B(n_69),
.Y(n_120)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_22),
.B(n_7),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx6_ASAP7_75t_SL g100 ( 
.A(n_74),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_22),
.B(n_7),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_15),
.Y(n_81)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_25),
.B(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_83),
.B(n_85),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_26),
.B(n_7),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_88),
.Y(n_107)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_17),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_26),
.B(n_6),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx6_ASAP7_75t_SL g101 ( 
.A(n_90),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_29),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_73),
.A2(n_34),
.B1(n_17),
.B2(n_33),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_104),
.A2(n_111),
.B1(n_128),
.B2(n_143),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_56),
.A2(n_42),
.B1(n_38),
.B2(n_39),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_49),
.B(n_42),
.C(n_38),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_113),
.B(n_122),
.Y(n_168)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_37),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_118),
.B(n_121),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_74),
.B(n_37),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_76),
.A2(n_42),
.B1(n_38),
.B2(n_28),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_41),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_127),
.B(n_139),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_52),
.A2(n_34),
.B1(n_33),
.B2(n_28),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_61),
.A2(n_39),
.B1(n_23),
.B2(n_28),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_132),
.A2(n_39),
.B1(n_59),
.B2(n_57),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_50),
.B(n_36),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_52),
.B(n_36),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_68),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_66),
.A2(n_71),
.B1(n_46),
.B2(n_48),
.Y(n_143)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

BUFx2_ASAP7_75t_SL g217 ( 
.A(n_145),
.Y(n_217)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_146),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_147),
.B(n_153),
.Y(n_202)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_148),
.Y(n_198)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_53),
.B(n_65),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_149),
.B(n_159),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_103),
.B(n_138),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_150),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_151),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_92),
.B(n_31),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_152),
.B(n_154),
.Y(n_206)
);

OAI32xp33_ASAP7_75t_L g153 ( 
.A1(n_120),
.A2(n_81),
.A3(n_54),
.B1(n_55),
.B2(n_70),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_93),
.B(n_31),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_136),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_157),
.B(n_158),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_100),
.Y(n_158)
);

INVx4_ASAP7_75t_SL g159 ( 
.A(n_101),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_101),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_160),
.B(n_167),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_109),
.B(n_94),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_161),
.B(n_166),
.Y(n_214)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_95),
.Y(n_163)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_132),
.A2(n_33),
.B1(n_45),
.B2(n_44),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_164),
.A2(n_184),
.B1(n_186),
.B2(n_191),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_99),
.B(n_45),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_117),
.B(n_98),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_144),
.Y(n_170)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_105),
.Y(n_171)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_172),
.Y(n_226)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_97),
.Y(n_173)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_173),
.Y(n_204)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_174),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_107),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_175),
.Y(n_222)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_178),
.A2(n_131),
.B1(n_102),
.B2(n_140),
.Y(n_210)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_119),
.Y(n_179)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_111),
.A2(n_91),
.B1(n_87),
.B2(n_84),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_182),
.A2(n_192),
.B1(n_155),
.B2(n_149),
.Y(n_223)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_108),
.Y(n_183)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_124),
.A2(n_44),
.B1(n_40),
.B2(n_27),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_98),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_185),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_96),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_188),
.Y(n_218)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_135),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_189),
.B(n_190),
.Y(n_221)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_102),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_96),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_104),
.A2(n_79),
.B1(n_78),
.B2(n_77),
.Y(n_192)
);

AND2x2_ASAP7_75t_SL g194 ( 
.A(n_162),
.B(n_113),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_194),
.B(n_209),
.C(n_216),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_162),
.A2(n_143),
.B1(n_128),
.B2(n_72),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_196),
.A2(n_210),
.B1(n_228),
.B2(n_232),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_168),
.B(n_161),
.C(n_152),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_168),
.B(n_107),
.C(n_129),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_154),
.A2(n_106),
.B(n_40),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_27),
.C(n_145),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_223),
.A2(n_227),
.B1(n_30),
.B2(n_165),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_166),
.A2(n_110),
.B(n_126),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_133),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_181),
.A2(n_106),
.B1(n_112),
.B2(n_68),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_153),
.A2(n_131),
.B1(n_115),
.B2(n_133),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_169),
.A2(n_115),
.B1(n_137),
.B2(n_140),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_163),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_233),
.B(n_234),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_173),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_235),
.A2(n_250),
.B(n_227),
.Y(n_272)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_236),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_196),
.A2(n_183),
.B1(n_189),
.B2(n_188),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_237),
.A2(n_266),
.B1(n_267),
.B2(n_211),
.Y(n_280)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_238),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_170),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_239),
.B(n_244),
.Y(n_279)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_212),
.Y(n_240)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_240),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_202),
.A2(n_137),
.B1(n_170),
.B2(n_171),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_241),
.A2(n_261),
.B1(n_210),
.B2(n_229),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_146),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_243),
.B(n_245),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_218),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_148),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_206),
.B(n_176),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_246),
.B(n_249),
.Y(n_288)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_224),
.Y(n_247)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_247),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_206),
.B(n_172),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_203),
.B(n_165),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_251),
.B(n_254),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_209),
.B(n_216),
.C(n_194),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_255),
.Y(n_271)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_199),
.Y(n_253)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_218),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_194),
.B(n_174),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_215),
.B(n_159),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_256),
.B(n_268),
.Y(n_297)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_199),
.Y(n_257)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_257),
.Y(n_298)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_204),
.Y(n_258)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_258),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_223),
.A2(n_180),
.B1(n_177),
.B2(n_190),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_259),
.A2(n_263),
.B1(n_217),
.B2(n_213),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_229),
.A2(n_191),
.B1(n_186),
.B2(n_151),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_260),
.A2(n_208),
.B1(n_212),
.B2(n_197),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_225),
.A2(n_39),
.B1(n_23),
.B2(n_110),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_221),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_262),
.B(n_265),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_229),
.A2(n_126),
.B1(n_30),
.B2(n_35),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_211),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_264),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_195),
.Y(n_265)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_224),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_204),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_270),
.B(n_272),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_241),
.A2(n_232),
.B1(n_219),
.B2(n_213),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_273),
.A2(n_277),
.B1(n_268),
.B2(n_240),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_235),
.A2(n_244),
.B1(n_254),
.B2(n_261),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_280),
.A2(n_195),
.B1(n_201),
.B2(n_198),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_281),
.A2(n_286),
.B1(n_290),
.B2(n_293),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_256),
.A2(n_215),
.B(n_231),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_282),
.A2(n_295),
.B(n_205),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_242),
.B(n_193),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_284),
.B(n_201),
.C(n_198),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_248),
.A2(n_193),
.B1(n_221),
.B2(n_207),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_248),
.A2(n_259),
.B1(n_262),
.B2(n_243),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_255),
.B(n_231),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_291),
.B(n_8),
.Y(n_326)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_292),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_245),
.A2(n_249),
.B1(n_246),
.B2(n_252),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_242),
.A2(n_263),
.B1(n_250),
.B2(n_258),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_300),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_236),
.A2(n_238),
.B(n_257),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_253),
.A2(n_207),
.B1(n_205),
.B2(n_208),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_301),
.B(n_302),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_277),
.A2(n_247),
.B1(n_264),
.B2(n_266),
.Y(n_302)
);

AOI21x1_ASAP7_75t_L g336 ( 
.A1(n_303),
.A2(n_272),
.B(n_282),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_310),
.C(n_316),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_274),
.B(n_265),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_307),
.B(n_313),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_308),
.B(n_317),
.Y(n_333)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_275),
.Y(n_309)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_309),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_271),
.B(n_197),
.C(n_226),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_274),
.B(n_230),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_279),
.B(n_230),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_314),
.B(n_327),
.Y(n_341)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_275),
.Y(n_315)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_315),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_271),
.B(n_226),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_296),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_297),
.B(n_30),
.Y(n_318)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_318),
.Y(n_351)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_276),
.Y(n_319)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_319),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_284),
.B(n_0),
.C(n_1),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_320),
.B(n_325),
.C(n_285),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_288),
.B(n_1),
.Y(n_321)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_321),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_288),
.B(n_1),
.Y(n_322)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_322),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_287),
.B(n_1),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_323),
.B(n_324),
.Y(n_349)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_276),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_293),
.B(n_2),
.C(n_3),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_326),
.B(n_297),
.Y(n_344)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_285),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_273),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_328),
.A2(n_322),
.B1(n_323),
.B2(n_306),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_311),
.A2(n_280),
.B1(n_287),
.B2(n_270),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_329),
.A2(n_348),
.B1(n_302),
.B2(n_303),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_291),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_334),
.B(n_345),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_336),
.A2(n_328),
.B(n_327),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_317),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_339),
.B(n_340),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_310),
.B(n_294),
.C(n_296),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_342),
.B(n_312),
.C(n_320),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_344),
.B(n_308),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_304),
.B(n_289),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_SL g346 ( 
.A(n_304),
.B(n_290),
.C(n_281),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_346),
.B(n_352),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_311),
.A2(n_286),
.B1(n_299),
.B2(n_298),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_305),
.B(n_295),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_350),
.B(n_318),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_321),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_301),
.Y(n_354)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_354),
.Y(n_375)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_335),
.Y(n_355)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_355),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_366),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_349),
.B(n_333),
.Y(n_357)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_357),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_333),
.A2(n_306),
.B1(n_312),
.B2(n_325),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_358),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_359),
.B(n_368),
.C(n_373),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_330),
.B(n_326),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_362),
.B(n_364),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_365),
.A2(n_351),
.B(n_341),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_332),
.A2(n_324),
.B1(n_319),
.B2(n_315),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_349),
.B(n_337),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_367),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_330),
.B(n_309),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_335),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_369),
.B(n_371),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_329),
.A2(n_348),
.B1(n_332),
.B2(n_336),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_370),
.B(n_345),
.Y(n_386)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_338),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_372),
.B(n_374),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_342),
.B(n_299),
.C(n_298),
.Y(n_373)
);

NAND3xp33_ASAP7_75t_L g374 ( 
.A(n_331),
.B(n_283),
.C(n_300),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_368),
.B(n_350),
.C(n_334),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_379),
.B(n_344),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_354),
.A2(n_343),
.B1(n_337),
.B2(n_346),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_382),
.A2(n_384),
.B1(n_278),
.B2(n_269),
.Y(n_402)
);

OA22x2_ASAP7_75t_L g384 ( 
.A1(n_370),
.A2(n_343),
.B1(n_347),
.B2(n_278),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_385),
.B(n_386),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_363),
.B(n_340),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_387),
.B(n_361),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_381),
.A2(n_356),
.B1(n_357),
.B2(n_367),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_392),
.A2(n_375),
.B1(n_388),
.B2(n_380),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_378),
.B(n_373),
.C(n_359),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_393),
.B(n_395),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_390),
.B(n_360),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_394),
.B(n_397),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_379),
.C(n_390),
.Y(n_395)
);

OR2x2_ASAP7_75t_L g404 ( 
.A(n_396),
.B(n_398),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_382),
.B(n_360),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_385),
.B(n_362),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_386),
.B(n_364),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_399),
.B(n_400),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_377),
.B(n_372),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_377),
.B(n_365),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_401),
.B(n_403),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_402),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_391),
.A2(n_381),
.B1(n_375),
.B2(n_389),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_406),
.B(n_411),
.Y(n_420)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_407),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_391),
.A2(n_384),
.B1(n_383),
.B2(n_269),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_401),
.A2(n_384),
.B1(n_376),
.B2(n_283),
.Y(n_412)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_412),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_400),
.A2(n_384),
.B1(n_3),
.B2(n_5),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_414),
.B(n_410),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_408),
.B(n_397),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_415),
.B(n_420),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_405),
.B(n_393),
.C(n_395),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_417),
.B(n_418),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_409),
.B(n_408),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_419),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_404),
.B(n_394),
.C(n_6),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_421),
.A2(n_422),
.B(n_404),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_409),
.B(n_2),
.C(n_14),
.Y(n_422)
);

INVx11_ASAP7_75t_L g425 ( 
.A(n_417),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_425),
.A2(n_413),
.B(n_8),
.Y(n_432)
);

NOR2xp67_ASAP7_75t_L g427 ( 
.A(n_415),
.B(n_410),
.Y(n_427)
);

A2O1A1O1Ixp25_ASAP7_75t_L g431 ( 
.A1(n_427),
.A2(n_429),
.B(n_416),
.C(n_413),
.D(n_10),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_428),
.B(n_422),
.C(n_423),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_430),
.A2(n_431),
.B(n_426),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_432),
.B(n_6),
.Y(n_433)
);

OAI21xp33_ASAP7_75t_L g435 ( 
.A1(n_433),
.A2(n_434),
.B(n_424),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_435),
.B(n_10),
.C(n_11),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_436),
.A2(n_13),
.B(n_14),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_437),
.A2(n_13),
.B(n_14),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_438),
.A2(n_13),
.B(n_380),
.Y(n_439)
);


endmodule