module fake_jpeg_18985_n_318 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_8),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_31),
.Y(n_50)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_19),
.B(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_40),
.A2(n_30),
.B1(n_29),
.B2(n_27),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_52),
.B1(n_40),
.B2(n_42),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_30),
.B1(n_31),
.B2(n_27),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_53),
.B1(n_57),
.B2(n_34),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_22),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_30),
.B1(n_29),
.B2(n_33),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_36),
.B1(n_34),
.B2(n_42),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_29),
.B1(n_18),
.B2(n_16),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_34),
.B1(n_40),
.B2(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_35),
.A2(n_18),
.B1(n_28),
.B2(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_59),
.B(n_61),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_60),
.A2(n_47),
.B1(n_39),
.B2(n_37),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_62),
.B(n_66),
.Y(n_118)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_35),
.B(n_24),
.C(n_19),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_64),
.A2(n_74),
.B(n_68),
.C(n_70),
.Y(n_117)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_53),
.B(n_20),
.Y(n_66)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_57),
.A2(n_24),
.B1(n_20),
.B2(n_21),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_34),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_69),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_34),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_75),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_22),
.B(n_21),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_71),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_72),
.A2(n_73),
.B1(n_47),
.B2(n_39),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_91),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_56),
.B(n_42),
.Y(n_75)
);

NAND2x1_ASAP7_75t_SL g76 ( 
.A(n_52),
.B(n_40),
.Y(n_76)
);

NOR2x1_ASAP7_75t_R g108 ( 
.A(n_76),
.B(n_82),
.Y(n_108)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_48),
.A2(n_25),
.B1(n_18),
.B2(n_32),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_32),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_83),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_43),
.A2(n_25),
.B1(n_18),
.B2(n_17),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_54),
.B(n_39),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_89),
.Y(n_122)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_86),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_46),
.A2(n_0),
.B(n_1),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_32),
.B(n_25),
.C(n_23),
.Y(n_97)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_46),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_90),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_93),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_124),
.B(n_82),
.Y(n_125)
);

OAI32xp33_ASAP7_75t_L g101 ( 
.A1(n_66),
.A2(n_58),
.A3(n_32),
.B1(n_17),
.B2(n_23),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_115),
.Y(n_141)
);

AND2x6_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_17),
.Y(n_107)
);

OAI221xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_117),
.B1(n_76),
.B2(n_91),
.C(n_79),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_62),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_85),
.B1(n_86),
.B2(n_80),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_119),
.A2(n_120),
.B1(n_69),
.B2(n_60),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_72),
.A2(n_83),
.B1(n_87),
.B2(n_71),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_38),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_148),
.Y(n_157)
);

NOR2x1_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_69),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_126),
.A2(n_98),
.B(n_111),
.Y(n_165)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_128),
.A2(n_139),
.B1(n_145),
.B2(n_108),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_115),
.B(n_89),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_130),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_81),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_132),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_102),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_102),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_134),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_114),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_88),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_135),
.B(n_140),
.Y(n_174)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_137),
.B(n_144),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_138),
.A2(n_146),
.B1(n_97),
.B2(n_111),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_76),
.B1(n_93),
.B2(n_92),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_99),
.B(n_92),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_95),
.B(n_77),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_143),
.B(n_149),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_99),
.B(n_37),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_112),
.A2(n_84),
.B1(n_39),
.B2(n_37),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_107),
.A2(n_37),
.B1(n_39),
.B2(n_84),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_103),
.B(n_63),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_96),
.Y(n_181)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_118),
.B(n_12),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_67),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_151),
.A2(n_124),
.B(n_106),
.Y(n_163)
);

INVxp67_ASAP7_75t_SL g152 ( 
.A(n_96),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_154),
.A2(n_159),
.B1(n_105),
.B2(n_109),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_155),
.A2(n_105),
.B1(n_109),
.B2(n_90),
.Y(n_202)
);

AOI322xp5_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_121),
.A3(n_117),
.B1(n_113),
.B2(n_110),
.C1(n_101),
.C2(n_124),
.Y(n_156)
);

MAJx2_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_171),
.C(n_134),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_163),
.B(n_165),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_136),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_162),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_128),
.A2(n_121),
.B1(n_116),
.B2(n_106),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_129),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_170),
.C(n_182),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_142),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_130),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_164),
.B(n_176),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_165),
.A2(n_173),
.B(n_67),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_123),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_126),
.B(n_15),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_131),
.A2(n_98),
.B(n_100),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_135),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_132),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_181),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_123),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_138),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_183),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_100),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_184),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_169),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_191),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_125),
.B(n_139),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_189),
.A2(n_190),
.B(n_199),
.Y(n_228)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_183),
.A2(n_144),
.B1(n_151),
.B2(n_146),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_192),
.A2(n_202),
.B1(n_215),
.B2(n_162),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_176),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_198),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_171),
.B(n_151),
.Y(n_194)
);

XNOR2x2_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_153),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_160),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_133),
.B(n_145),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_208),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_96),
.C(n_63),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_211),
.C(n_178),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_161),
.B(n_105),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_210),
.Y(n_234)
);

BUFx12f_ASAP7_75t_SL g206 ( 
.A(n_157),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_206),
.A2(n_179),
.B(n_172),
.Y(n_216)
);

NOR3xp33_ASAP7_75t_L g208 ( 
.A(n_164),
.B(n_137),
.C(n_11),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_172),
.A2(n_11),
.B(n_15),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_209),
.A2(n_212),
.B(n_153),
.Y(n_231)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_37),
.C(n_38),
.Y(n_211)
);

BUFx12_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_167),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_214),
.B(n_158),
.Y(n_220)
);

AO22x1_ASAP7_75t_SL g215 ( 
.A1(n_159),
.A2(n_38),
.B1(n_28),
.B2(n_26),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_216),
.A2(n_213),
.B(n_192),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_217),
.B(n_199),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_218),
.A2(n_203),
.B1(n_185),
.B2(n_215),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_154),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_221),
.Y(n_250)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_174),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_207),
.B(n_177),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_186),
.Y(n_241)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_188),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_174),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_237),
.Y(n_256)
);

MAJx2_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_194),
.C(n_212),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_231),
.A2(n_7),
.B1(n_13),
.B2(n_10),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_236),
.C(n_238),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_155),
.C(n_178),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_180),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_189),
.B(n_17),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_245),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_241),
.Y(n_262)
);

AO22x1_ASAP7_75t_L g242 ( 
.A1(n_234),
.A2(n_193),
.B1(n_205),
.B2(n_188),
.Y(n_242)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_242),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_224),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_251),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_244),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_247),
.A2(n_229),
.B1(n_225),
.B2(n_233),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_201),
.Y(n_248)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_222),
.A2(n_209),
.B1(n_200),
.B2(n_215),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_249),
.A2(n_257),
.B1(n_6),
.B2(n_10),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

A2O1A1O1Ixp25_ASAP7_75t_L g253 ( 
.A1(n_230),
.A2(n_211),
.B(n_213),
.C(n_9),
.D(n_12),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_231),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_226),
.B(n_8),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_254),
.A2(n_255),
.B1(n_236),
.B2(n_228),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_218),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_271),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_261),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_232),
.C(n_221),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_266),
.C(n_274),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_255),
.A2(n_228),
.B1(n_237),
.B2(n_219),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_5),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_217),
.C(n_238),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_251),
.A2(n_253),
.B1(n_246),
.B2(n_240),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_270),
.A2(n_256),
.B(n_247),
.Y(n_277)
);

XOR2x2_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_6),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_273),
.B(n_7),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_38),
.C(n_28),
.Y(n_274)
);

OAI221xp5_ASAP7_75t_L g275 ( 
.A1(n_270),
.A2(n_248),
.B1(n_256),
.B2(n_250),
.C(n_252),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_282),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g276 ( 
.A(n_262),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_279),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_0),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_5),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_281),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_269),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_9),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_285),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_0),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_259),
.B(n_26),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_274),
.C(n_258),
.Y(n_294)
);

NOR2xp67_ASAP7_75t_L g288 ( 
.A(n_286),
.B(n_271),
.Y(n_288)
);

NOR2xp67_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_1),
.Y(n_299)
);

NOR2x1_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_258),
.Y(n_290)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_290),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_263),
.C(n_266),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_38),
.Y(n_300)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_294),
.Y(n_305)
);

NOR2xp67_ASAP7_75t_SL g295 ( 
.A(n_284),
.B(n_272),
.Y(n_295)
);

OAI21x1_ASAP7_75t_L g304 ( 
.A1(n_295),
.A2(n_2),
.B(n_3),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_296),
.B(n_1),
.Y(n_301)
);

AOI21x1_ASAP7_75t_L g298 ( 
.A1(n_289),
.A2(n_278),
.B(n_2),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_301),
.Y(n_307)
);

AOI21x1_ASAP7_75t_L g310 ( 
.A1(n_299),
.A2(n_304),
.B(n_301),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_300),
.A2(n_38),
.B(n_4),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_38),
.C(n_3),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_297),
.C(n_38),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_2),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_296),
.Y(n_308)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_308),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_312),
.C(n_4),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_310),
.A2(n_311),
.B(n_305),
.Y(n_314)
);

MAJx2_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_290),
.C(n_292),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_314),
.B(n_315),
.C(n_307),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_313),
.B(n_308),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_317),
.Y(n_318)
);


endmodule