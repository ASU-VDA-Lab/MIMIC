module fake_jpeg_334_n_445 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_445);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_445;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_SL g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_54),
.Y(n_133)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_55),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_56),
.Y(n_136)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_28),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_58),
.B(n_66),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_59),
.Y(n_160)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_21),
.B(n_10),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_61),
.B(n_75),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_62),
.Y(n_171)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

BUFx16f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_64),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_25),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_49),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_68),
.Y(n_182)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

OR2x2_ASAP7_75t_SL g70 ( 
.A(n_22),
.B(n_9),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_70),
.B(n_83),
.Y(n_129)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_73),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_74),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_21),
.B(n_9),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_30),
.B(n_11),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_78),
.B(n_88),
.Y(n_138)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_82),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_35),
.Y(n_82)
);

NAND2xp33_ASAP7_75t_SL g83 ( 
.A(n_46),
.B(n_0),
.Y(n_83)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_22),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_86),
.A2(n_27),
.B1(n_47),
.B2(n_42),
.Y(n_174)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_87),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_20),
.B(n_12),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_35),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_90),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_35),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_91),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_11),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_93),
.B(n_99),
.Y(n_147)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

BUFx10_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_30),
.B(n_13),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_24),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_103),
.Y(n_131)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_24),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_24),
.Y(n_105)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_106),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_19),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_108),
.Y(n_168)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_23),
.Y(n_109)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_109),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_32),
.B(n_13),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_110),
.B(n_16),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_44),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_112),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_19),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_94),
.A2(n_53),
.B1(n_40),
.B2(n_26),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_142),
.A2(n_97),
.B1(n_80),
.B2(n_77),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_143),
.B(n_74),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_101),
.A2(n_36),
.B1(n_31),
.B2(n_18),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g217 ( 
.A1(n_148),
.A2(n_170),
.B1(n_178),
.B2(n_95),
.Y(n_217)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_149),
.Y(n_194)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_54),
.Y(n_153)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_153),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_63),
.B(n_32),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_154),
.B(n_155),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_60),
.B(n_53),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_64),
.B(n_40),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_156),
.B(n_159),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_64),
.B(n_36),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_65),
.Y(n_161)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_161),
.Y(n_229)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_69),
.Y(n_162)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_162),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_163),
.B(n_177),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_87),
.B(n_31),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_165),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_79),
.B(n_18),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_91),
.B(n_45),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_169),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_73),
.B(n_45),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_56),
.A2(n_27),
.B1(n_47),
.B2(n_42),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_92),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_183),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_174),
.A2(n_95),
.B1(n_102),
.B2(n_98),
.Y(n_201)
);

AND2x2_ASAP7_75t_SL g176 ( 
.A(n_70),
.B(n_23),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_176),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_83),
.B(n_34),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_68),
.A2(n_71),
.B1(n_84),
.B2(n_106),
.Y(n_178)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_96),
.Y(n_181)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_105),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_108),
.Y(n_184)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_184),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_52),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_186),
.B(n_191),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_118),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_187),
.B(n_198),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_188),
.B(n_189),
.Y(n_264)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_138),
.A2(n_86),
.A3(n_34),
.B1(n_52),
.B2(n_39),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_125),
.Y(n_190)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_190),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_129),
.B(n_39),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_192),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_146),
.Y(n_196)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_196),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_122),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_134),
.B(n_62),
.C(n_104),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_200),
.B(n_216),
.C(n_223),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_201),
.A2(n_235),
.B1(n_178),
.B2(n_124),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_128),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_202),
.B(n_204),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_136),
.Y(n_203)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_203),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_131),
.Y(n_204)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_133),
.Y(n_205)
);

NAND2xp33_ASAP7_75t_SL g258 ( 
.A(n_205),
.B(n_208),
.Y(n_258)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_132),
.Y(n_206)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_206),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_145),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_207),
.B(n_212),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_117),
.Y(n_208)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_125),
.Y(n_209)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_209),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_211),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_127),
.B(n_67),
.Y(n_212)
);

OR2x4_ASAP7_75t_L g214 ( 
.A(n_129),
.B(n_147),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_225),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_115),
.Y(n_215)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_215),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_107),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_217),
.A2(n_219),
.B1(n_237),
.B2(n_238),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_218),
.A2(n_136),
.B1(n_171),
.B2(n_160),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_120),
.A2(n_74),
.B1(n_107),
.B2(n_59),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_141),
.B(n_167),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_220),
.B(n_226),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_119),
.B(n_76),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_221),
.B(n_230),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_148),
.A2(n_57),
.B(n_72),
.Y(n_223)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_224),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_113),
.B(n_14),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g226 ( 
.A(n_132),
.Y(n_226)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_114),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_227),
.Y(n_268)
);

A2O1A1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_143),
.A2(n_57),
.B(n_72),
.C(n_14),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_L g263 ( 
.A1(n_228),
.A2(n_241),
.B(n_123),
.C(n_130),
.Y(n_263)
);

AO22x1_ASAP7_75t_SL g230 ( 
.A1(n_121),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_139),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_233),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_170),
.A2(n_3),
.B1(n_6),
.B2(n_157),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_113),
.B(n_133),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_236),
.B(n_239),
.Y(n_283)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_158),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_168),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_126),
.B(n_6),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_151),
.B(n_115),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_123),
.Y(n_254)
);

A2O1A1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_140),
.A2(n_182),
.B(n_173),
.C(n_116),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_114),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_242),
.A2(n_209),
.B1(n_196),
.B2(n_206),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_151),
.B(n_182),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_243),
.A2(n_152),
.B1(n_220),
.B2(n_192),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_244),
.A2(n_250),
.B1(n_279),
.B2(n_286),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_217),
.A2(n_194),
.B1(n_191),
.B2(n_201),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_245),
.A2(n_248),
.B1(n_251),
.B2(n_252),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_214),
.A2(n_144),
.B1(n_124),
.B2(n_135),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_185),
.A2(n_137),
.B1(n_150),
.B2(n_135),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_221),
.A2(n_160),
.B1(n_171),
.B2(n_180),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_254),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_263),
.A2(n_271),
.B1(n_279),
.B2(n_264),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_186),
.B(n_199),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_266),
.B(n_282),
.C(n_257),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_239),
.A2(n_180),
.B1(n_144),
.B2(n_130),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_269),
.A2(n_276),
.B1(n_278),
.B2(n_285),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_200),
.A2(n_228),
.B1(n_189),
.B2(n_193),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_217),
.A2(n_152),
.B1(n_211),
.B2(n_230),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_277),
.A2(n_280),
.B1(n_226),
.B2(n_254),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_217),
.A2(n_241),
.B1(n_188),
.B2(n_195),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_188),
.A2(n_223),
.B1(n_230),
.B2(n_243),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_229),
.A2(n_238),
.B1(n_237),
.B2(n_231),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_213),
.B(n_232),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_210),
.B(n_197),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_287),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_216),
.A2(n_231),
.B1(n_197),
.B2(n_240),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_224),
.A2(n_203),
.B1(n_227),
.B2(n_216),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_240),
.A2(n_190),
.B1(n_234),
.B2(n_222),
.Y(n_287)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_288),
.Y(n_289)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_285),
.Y(n_292)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_292),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_260),
.B(n_282),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_293),
.B(n_302),
.Y(n_337)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_294),
.Y(n_339)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_265),
.Y(n_296)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_296),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_242),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_306),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_263),
.A2(n_205),
.B(n_206),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_298),
.A2(n_313),
.B(n_316),
.Y(n_341)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_299),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_301),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_266),
.B(n_226),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_265),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_303),
.B(n_304),
.Y(n_334)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_287),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_259),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_257),
.B(n_264),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_307),
.B(n_252),
.C(n_274),
.Y(n_325)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_249),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_308),
.B(n_309),
.Y(n_342)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_249),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_261),
.B(n_270),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_310),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_311),
.B(n_321),
.Y(n_335)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_255),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_312),
.B(n_315),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_281),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_314),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_259),
.B(n_264),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_284),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_278),
.A2(n_276),
.B(n_258),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_317),
.A2(n_320),
.B(n_313),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_247),
.A2(n_267),
.B(n_246),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_318),
.A2(n_298),
.B(n_317),
.Y(n_323)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_255),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_319),
.A2(n_312),
.B1(n_309),
.B2(n_308),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_247),
.A2(n_250),
.B1(n_268),
.B2(n_246),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_275),
.B(n_253),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_253),
.B(n_275),
.Y(n_322)
);

MAJx2_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_256),
.C(n_315),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_323),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_269),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_324),
.B(n_328),
.C(n_338),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_325),
.B(n_319),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_274),
.Y(n_328)
);

AO22x1_ASAP7_75t_L g329 ( 
.A1(n_300),
.A2(n_255),
.B1(n_251),
.B2(n_262),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_329),
.B(n_346),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_290),
.A2(n_273),
.B1(n_262),
.B2(n_256),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_330),
.A2(n_329),
.B1(n_347),
.B2(n_339),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_336),
.B(n_296),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_295),
.B(n_318),
.C(n_311),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_343),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_294),
.A2(n_300),
.B(n_304),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_344),
.Y(n_363)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_345),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_320),
.A2(n_295),
.B(n_291),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_297),
.B(n_291),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_349),
.B(n_324),
.C(n_325),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_344),
.A2(n_290),
.B1(n_292),
.B2(n_316),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_351),
.A2(n_353),
.B1(n_365),
.B2(n_329),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_323),
.A2(n_305),
.B1(n_289),
.B2(n_321),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_342),
.Y(n_354)
);

CKINVDCx14_ASAP7_75t_R g382 ( 
.A(n_354),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_357),
.B(n_370),
.Y(n_377)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_340),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_358),
.Y(n_389)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_340),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_359),
.A2(n_367),
.B1(n_368),
.B2(n_371),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_327),
.B(n_303),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_360),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_327),
.B(n_301),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_362),
.A2(n_366),
.B(n_326),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_364),
.B(n_335),
.C(n_336),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_333),
.A2(n_289),
.B1(n_343),
.B2(n_347),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_345),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_339),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_331),
.B(n_334),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_369),
.A2(n_326),
.B1(n_354),
.B2(n_350),
.Y(n_388)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_333),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_363),
.A2(n_331),
.B1(n_346),
.B2(n_332),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_372),
.A2(n_361),
.B1(n_386),
.B2(n_378),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_370),
.B(n_338),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_373),
.B(n_374),
.C(n_376),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_355),
.B(n_335),
.C(n_328),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_356),
.A2(n_341),
.B(n_332),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_378),
.B(n_352),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_355),
.B(n_349),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_379),
.B(n_386),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_364),
.B(n_341),
.C(n_348),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_380),
.B(n_383),
.C(n_385),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_337),
.Y(n_383)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_384),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_356),
.B(n_348),
.C(n_337),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_361),
.B(n_330),
.Y(n_386)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_387),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_388),
.B(n_351),
.Y(n_391)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_391),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_385),
.B(n_359),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_392),
.B(n_400),
.Y(n_408)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_389),
.Y(n_394)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_394),
.Y(n_409)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_389),
.Y(n_396)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_396),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_398),
.B(n_401),
.Y(n_413)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_389),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_381),
.B(n_367),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_402),
.A2(n_403),
.B1(n_350),
.B2(n_383),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_382),
.B(n_358),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_390),
.A2(n_384),
.B1(n_363),
.B2(n_372),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_404),
.A2(n_390),
.B1(n_353),
.B2(n_375),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_395),
.B(n_376),
.C(n_379),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_406),
.B(n_407),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_395),
.B(n_373),
.C(n_380),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_399),
.B(n_377),
.C(n_374),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_410),
.B(n_412),
.C(n_397),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_411),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_399),
.B(n_377),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_415),
.B(n_421),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_406),
.B(n_397),
.C(n_402),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_417),
.B(n_419),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_408),
.B(n_393),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_409),
.Y(n_420)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_420),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_413),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_413),
.B(n_391),
.Y(n_422)
);

INVxp33_ASAP7_75t_L g426 ( 
.A(n_422),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_423),
.A2(n_416),
.B1(n_368),
.B2(n_352),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_416),
.A2(n_405),
.B(n_404),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_424),
.A2(n_396),
.B(n_365),
.Y(n_435)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_425),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_418),
.B(n_407),
.C(n_410),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_427),
.B(n_417),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_431),
.B(n_435),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_426),
.A2(n_423),
.B1(n_414),
.B2(n_394),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_432),
.B(n_433),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_424),
.B(n_412),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_434),
.A2(n_428),
.B(n_430),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_438),
.A2(n_426),
.B(n_437),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_439),
.B(n_440),
.C(n_427),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_436),
.Y(n_440)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_441),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_442),
.A2(n_435),
.B1(n_429),
.B2(n_433),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_443),
.B(n_425),
.C(n_415),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_444),
.B(n_371),
.Y(n_445)
);


endmodule