module fake_aes_7638_n_30 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_30);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_7), .Y(n_10) );
NOR2xp33_ASAP7_75t_R g11 ( .A(n_2), .B(n_8), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_3), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_3), .Y(n_14) );
A2O1A1Ixp33_ASAP7_75t_L g15 ( .A1(n_12), .A2(n_0), .B(n_1), .C(n_2), .Y(n_15) );
AOI21xp5_ASAP7_75t_L g16 ( .A1(n_12), .A2(n_0), .B(n_1), .Y(n_16) );
AOI21xp5_ASAP7_75t_L g17 ( .A1(n_12), .A2(n_0), .B(n_1), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_15), .B(n_10), .Y(n_18) );
OAI22xp5_ASAP7_75t_L g19 ( .A1(n_16), .A2(n_13), .B1(n_10), .B2(n_14), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
OR2x2_ASAP7_75t_L g21 ( .A(n_18), .B(n_4), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_18), .B(n_17), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_22), .B(n_19), .Y(n_23) );
AOI222xp33_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_20), .B1(n_22), .B2(n_21), .C1(n_11), .C2(n_5), .Y(n_24) );
AOI221xp5_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_22), .B1(n_21), .B2(n_11), .C(n_8), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
BUFx2_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
BUFx2_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
OAI22xp5_ASAP7_75t_SL g29 ( .A1(n_26), .A2(n_23), .B1(n_6), .B2(n_7), .Y(n_29) );
AOI22xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_27), .B1(n_28), .B2(n_9), .Y(n_30) );
endmodule