module fake_jpeg_4942_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_47),
.Y(n_67)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_44),
.Y(n_60)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_29),
.B1(n_32),
.B2(n_28),
.Y(n_65)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_27),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_49),
.B(n_52),
.Y(n_94)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_54),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_27),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_32),
.B1(n_29),
.B2(n_31),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_53),
.A2(n_23),
.B1(n_19),
.B2(n_20),
.Y(n_86)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx5_ASAP7_75t_SL g95 ( 
.A(n_56),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_20),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_63),
.Y(n_92)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_39),
.B(n_32),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_29),
.B1(n_23),
.B2(n_33),
.Y(n_80)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_18),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_71),
.Y(n_93)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_43),
.B1(n_29),
.B2(n_41),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_77),
.A2(n_98),
.B1(n_59),
.B2(n_71),
.Y(n_101)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_88),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_87),
.B1(n_90),
.B2(n_64),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_46),
.B1(n_40),
.B2(n_31),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_86),
.B1(n_89),
.B2(n_91),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_74),
.A2(n_23),
.B1(n_19),
.B2(n_21),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

AO22x2_ASAP7_75t_L g89 ( 
.A1(n_49),
.A2(n_46),
.B1(n_40),
.B2(n_38),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_74),
.A2(n_21),
.B1(n_33),
.B2(n_17),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_49),
.A2(n_17),
.B1(n_18),
.B2(n_21),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_67),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_97),
.B(n_39),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_56),
.A2(n_33),
.B1(n_46),
.B2(n_40),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_99),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_67),
.B(n_57),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_100),
.A2(n_113),
.B(n_78),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_114),
.B1(n_118),
.B2(n_83),
.Y(n_134)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_103),
.B(n_106),
.Y(n_152)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_105),
.Y(n_146)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_107),
.A2(n_81),
.B1(n_75),
.B2(n_78),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_57),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_121),
.Y(n_130)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_111),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_77),
.A2(n_52),
.B(n_73),
.C(n_62),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_79),
.A2(n_72),
.B1(n_64),
.B2(n_52),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_112),
.A2(n_120),
.B1(n_122),
.B2(n_126),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_60),
.B(n_58),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_66),
.B1(n_54),
.B2(n_51),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_119),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_73),
.B1(n_50),
.B2(n_25),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_98),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_55),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_92),
.B(n_48),
.Y(n_123)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_96),
.C(n_39),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_92),
.B(n_48),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_128),
.Y(n_138)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_127),
.Y(n_129)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_133),
.B(n_135),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_136),
.B1(n_143),
.B2(n_155),
.Y(n_159)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_94),
.B1(n_92),
.B2(n_82),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_137),
.A2(n_145),
.B1(n_149),
.B2(n_129),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_94),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_142),
.Y(n_163)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_140),
.B(n_141),
.Y(n_158)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_122),
.A2(n_91),
.B1(n_82),
.B2(n_75),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_126),
.A2(n_81),
.B1(n_82),
.B2(n_75),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_144),
.A2(n_150),
.B(n_30),
.Y(n_185)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_121),
.B(n_39),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_147),
.A2(n_106),
.B(n_73),
.Y(n_172)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_96),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_156),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_103),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_111),
.A2(n_88),
.B1(n_99),
.B2(n_81),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_113),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_160),
.A2(n_172),
.B(n_138),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_142),
.B1(n_132),
.B2(n_102),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_161),
.A2(n_165),
.B1(n_171),
.B2(n_177),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_128),
.B1(n_118),
.B2(n_123),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_162),
.A2(n_180),
.B1(n_184),
.B2(n_141),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_156),
.A2(n_125),
.B1(n_109),
.B2(n_102),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_167),
.Y(n_188)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_100),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_175),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_155),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_169),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_157),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_174),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_108),
.B1(n_124),
.B2(n_116),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_131),
.A2(n_120),
.B1(n_34),
.B2(n_30),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_SL g199 ( 
.A1(n_173),
.A2(n_185),
.B(n_147),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_146),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_146),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_76),
.Y(n_176)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_136),
.A2(n_76),
.B1(n_38),
.B2(n_50),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_178),
.B(n_186),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_55),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_26),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_154),
.A2(n_38),
.B1(n_25),
.B2(n_34),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_30),
.C(n_26),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_140),
.B1(n_133),
.B2(n_129),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_138),
.A2(n_25),
.B1(n_30),
.B2(n_103),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_187),
.A2(n_194),
.B(n_199),
.Y(n_236)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_193),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_182),
.Y(n_190)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_190),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_153),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_207),
.C(n_208),
.Y(n_225)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

OA21x2_ASAP7_75t_L g194 ( 
.A1(n_170),
.A2(n_147),
.B(n_144),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_198),
.A2(n_200),
.B1(n_159),
.B2(n_178),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_162),
.A2(n_131),
.B1(n_147),
.B2(n_139),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_201),
.A2(n_206),
.B1(n_172),
.B2(n_173),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_202),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_182),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_204),
.B(n_175),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_169),
.A2(n_137),
.B1(n_149),
.B2(n_30),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_26),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_179),
.Y(n_209)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_176),
.Y(n_217)
);

INVxp33_ASAP7_75t_SL g211 ( 
.A(n_158),
.Y(n_211)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_26),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_186),
.C(n_174),
.Y(n_227)
);

AOI32xp33_ASAP7_75t_L g213 ( 
.A1(n_185),
.A2(n_16),
.A3(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_213),
.B(n_177),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_159),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_214),
.Y(n_215)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_216),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_217),
.B(n_227),
.C(n_232),
.Y(n_260)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_218),
.B(n_219),
.Y(n_245)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_221),
.A2(n_222),
.B1(n_203),
.B2(n_194),
.Y(n_250)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_223),
.B(n_234),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_168),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_228),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_166),
.Y(n_226)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_226),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_201),
.B(n_163),
.Y(n_228)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_229),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_197),
.A2(n_165),
.B1(n_161),
.B2(n_160),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_231),
.A2(n_239),
.B(n_209),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_165),
.C(n_163),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_164),
.Y(n_233)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_164),
.C(n_184),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_3),
.C(n_4),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_187),
.A2(n_180),
.B(n_158),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_16),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_210),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_235),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_242),
.B(n_257),
.Y(n_280)
);

NOR2x1_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_193),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_243),
.A2(n_244),
.B(n_259),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_215),
.A2(n_205),
.B1(n_198),
.B2(n_194),
.Y(n_244)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_247),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_203),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_264),
.C(n_265),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_250),
.A2(n_236),
.B1(n_240),
.B2(n_6),
.Y(n_274)
);

MAJx2_ASAP7_75t_L g278 ( 
.A(n_252),
.B(n_4),
.C(n_5),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_190),
.Y(n_254)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_254),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_227),
.B(n_189),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_256),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_238),
.B(n_202),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_220),
.Y(n_257)
);

OA21x2_ASAP7_75t_L g259 ( 
.A1(n_230),
.A2(n_0),
.B(n_2),
.Y(n_259)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_226),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_263),
.A2(n_241),
.B(n_237),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_225),
.B(n_3),
.C(n_4),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_243),
.A2(n_222),
.B1(n_241),
.B2(n_237),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_267),
.A2(n_273),
.B1(n_259),
.B2(n_247),
.Y(n_296)
);

NOR3xp33_ASAP7_75t_SL g268 ( 
.A(n_252),
.B(n_216),
.C(n_228),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_274),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_225),
.C(n_232),
.Y(n_270)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_283),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_251),
.A2(n_231),
.B1(n_236),
.B2(n_217),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_248),
.C(n_254),
.Y(n_275)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_4),
.C(n_5),
.Y(n_277)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_277),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_264),
.Y(n_285)
);

NOR2xp67_ASAP7_75t_SL g279 ( 
.A(n_242),
.B(n_11),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_282),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_261),
.B(n_11),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_281),
.B(n_245),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_6),
.C(n_7),
.Y(n_282)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_282),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_246),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_286),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_249),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_291),
.C(n_266),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_250),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_267),
.A2(n_253),
.B1(n_257),
.B2(n_262),
.Y(n_293)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_293),
.Y(n_309)
);

FAx1_ASAP7_75t_SL g294 ( 
.A(n_268),
.B(n_244),
.CI(n_265),
.CON(n_294),
.SN(n_294)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_295),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_296),
.A2(n_298),
.B(n_278),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_284),
.A2(n_276),
.B1(n_269),
.B2(n_272),
.Y(n_297)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_297),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_276),
.A2(n_259),
.B1(n_7),
.B2(n_8),
.Y(n_298)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_302),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_280),
.B(n_270),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_303),
.A2(n_308),
.B(n_312),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_307),
.C(n_310),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_300),
.B(n_266),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_313),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_277),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_6),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_288),
.C(n_291),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_292),
.A2(n_11),
.B(n_15),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_296),
.A2(n_10),
.B(n_15),
.Y(n_313)
);

AOI21xp33_ASAP7_75t_L g314 ( 
.A1(n_294),
.A2(n_12),
.B(n_14),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_314),
.A2(n_299),
.B1(n_294),
.B2(n_286),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_298),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_322),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_321),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_285),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_310),
.C(n_311),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_14),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_324),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_6),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_307),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_328),
.A2(n_329),
.B(n_330),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_16),
.Y(n_329)
);

XNOR2x1_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_322),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_7),
.Y(n_331)
);

OAI21x1_ASAP7_75t_L g333 ( 
.A1(n_331),
.A2(n_318),
.B(n_9),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_316),
.B(n_7),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_332),
.B(n_8),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_337),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_326),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_334),
.A2(n_336),
.B(n_330),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_319),
.Y(n_336)
);

MAJx2_ASAP7_75t_L g340 ( 
.A(n_338),
.B(n_335),
.C(n_327),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_339),
.C(n_8),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_8),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_9),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_9),
.Y(n_344)
);


endmodule