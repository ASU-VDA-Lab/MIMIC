module fake_aes_10811_n_880 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_92, n_11, n_223, n_25, n_30, n_59, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_880);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_880;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_878;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_567;
wire n_809;
wire n_580;
wire n_502;
wire n_543;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_230;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_876;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_466;
wire n_302;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_716;
wire n_653;
wire n_260;
wire n_806;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_573;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_837;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_68), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_193), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_144), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_169), .Y(n_231) );
CKINVDCx16_ASAP7_75t_R g232 ( .A(n_5), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_183), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_105), .Y(n_234) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_48), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_170), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_94), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_143), .Y(n_238) );
BUFx5_ASAP7_75t_L g239 ( .A(n_158), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_134), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_0), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_76), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_139), .Y(n_243) );
BUFx10_ASAP7_75t_L g244 ( .A(n_173), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_128), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_4), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_75), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_168), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_8), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_200), .Y(n_250) );
CKINVDCx16_ASAP7_75t_R g251 ( .A(n_204), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_214), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_30), .Y(n_253) );
BUFx3_ASAP7_75t_L g254 ( .A(n_26), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_163), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_41), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_28), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_12), .Y(n_258) );
BUFx2_ASAP7_75t_SL g259 ( .A(n_137), .Y(n_259) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_125), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_127), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_151), .Y(n_262) );
CKINVDCx14_ASAP7_75t_R g263 ( .A(n_51), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_153), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_58), .Y(n_265) );
BUFx3_ASAP7_75t_L g266 ( .A(n_55), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_10), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_218), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_62), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_100), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_123), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_101), .Y(n_272) );
INVx1_ASAP7_75t_SL g273 ( .A(n_161), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_208), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_219), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_25), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_224), .Y(n_277) );
CKINVDCx20_ASAP7_75t_R g278 ( .A(n_138), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_164), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_56), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_199), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_15), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_201), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_179), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_132), .Y(n_285) );
INVx1_ASAP7_75t_SL g286 ( .A(n_82), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_102), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_42), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_135), .B(n_14), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_43), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_186), .Y(n_291) );
BUFx3_ASAP7_75t_L g292 ( .A(n_145), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_37), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_83), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_74), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_180), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_87), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_97), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_67), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_57), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_178), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_22), .Y(n_302) );
CKINVDCx20_ASAP7_75t_R g303 ( .A(n_203), .Y(n_303) );
INVxp67_ASAP7_75t_L g304 ( .A(n_90), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_120), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_33), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_24), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_162), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_60), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_160), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_209), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_78), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_21), .Y(n_313) );
CKINVDCx20_ASAP7_75t_R g314 ( .A(n_202), .Y(n_314) );
CKINVDCx16_ASAP7_75t_R g315 ( .A(n_194), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_19), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_177), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_133), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_49), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_181), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_53), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_166), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_140), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_79), .Y(n_324) );
CKINVDCx20_ASAP7_75t_R g325 ( .A(n_99), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_206), .Y(n_326) );
BUFx3_ASAP7_75t_L g327 ( .A(n_216), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_225), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_98), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_148), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_89), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_187), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_159), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_131), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_107), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_44), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_12), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_205), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_220), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_189), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_232), .A2(n_315), .B1(n_251), .B2(n_337), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_235), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_253), .B(n_0), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_253), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_287), .B(n_1), .Y(n_345) );
BUFx2_ASAP7_75t_L g346 ( .A(n_316), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_244), .Y(n_347) );
INVx5_ASAP7_75t_L g348 ( .A(n_235), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_287), .Y(n_349) );
BUFx3_ASAP7_75t_L g350 ( .A(n_254), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_326), .Y(n_351) );
INVx6_ASAP7_75t_L g352 ( .A(n_244), .Y(n_352) );
INVx2_ASAP7_75t_SL g353 ( .A(n_326), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_239), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_239), .Y(n_355) );
INVx2_ASAP7_75t_SL g356 ( .A(n_318), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_249), .Y(n_357) );
BUFx8_ASAP7_75t_SL g358 ( .A(n_267), .Y(n_358) );
INVx6_ASAP7_75t_L g359 ( .A(n_239), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_239), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_241), .Y(n_361) );
INVx6_ASAP7_75t_L g362 ( .A(n_239), .Y(n_362) );
BUFx8_ASAP7_75t_SL g363 ( .A(n_278), .Y(n_363) );
BUFx12f_ASAP7_75t_L g364 ( .A(n_228), .Y(n_364) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_235), .Y(n_365) );
OAI22xp5_ASAP7_75t_SL g366 ( .A1(n_246), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_263), .B(n_5), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_263), .Y(n_368) );
INVx5_ASAP7_75t_L g369 ( .A(n_235), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_353), .B(n_282), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_353), .B(n_304), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_354), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_357), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_347), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_354), .Y(n_375) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_342), .Y(n_376) );
INVx8_ASAP7_75t_L g377 ( .A(n_368), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_343), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_355), .Y(n_379) );
NOR2x1p5_ASAP7_75t_L g380 ( .A(n_347), .B(n_258), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_352), .B(n_304), .Y(n_381) );
BUFx2_ASAP7_75t_L g382 ( .A(n_361), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_345), .Y(n_383) );
INVx4_ASAP7_75t_L g384 ( .A(n_359), .Y(n_384) );
INVx3_ASAP7_75t_L g385 ( .A(n_355), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_344), .B(n_231), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_360), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_360), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_347), .B(n_239), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_367), .Y(n_390) );
INVxp33_ASAP7_75t_L g391 ( .A(n_367), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_359), .Y(n_392) );
AOI21x1_ASAP7_75t_L g393 ( .A1(n_349), .A2(n_230), .B(n_229), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_351), .B(n_234), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_346), .B(n_289), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_359), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_356), .B(n_259), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_356), .B(n_266), .Y(n_398) );
INVx3_ASAP7_75t_L g399 ( .A(n_362), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_371), .B(n_368), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_391), .B(n_350), .Y(n_401) );
INVx6_ASAP7_75t_L g402 ( .A(n_380), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_385), .Y(n_403) );
BUFx3_ASAP7_75t_L g404 ( .A(n_382), .Y(n_404) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_378), .B(n_364), .Y(n_405) );
OAI22xp33_ASAP7_75t_SL g406 ( .A1(n_390), .A2(n_362), .B1(n_236), .B2(n_238), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_370), .B(n_341), .Y(n_407) );
INVx3_ASAP7_75t_L g408 ( .A(n_374), .Y(n_408) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_383), .B(n_364), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_370), .B(n_386), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_373), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_394), .B(n_352), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_374), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_391), .B(n_350), .Y(n_414) );
INVx2_ASAP7_75t_SL g415 ( .A(n_395), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_398), .B(n_352), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_385), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_397), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_397), .B(n_273), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_398), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_395), .A2(n_366), .B1(n_314), .B2(n_303), .C(n_325), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_381), .B(n_286), .Y(n_422) );
NOR3xp33_ASAP7_75t_L g423 ( .A(n_389), .B(n_393), .C(n_243), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_389), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_377), .B(n_237), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_372), .B(n_233), .Y(n_426) );
AND2x6_ASAP7_75t_L g427 ( .A(n_392), .B(n_247), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_372), .B(n_375), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_385), .Y(n_429) );
NAND2xp5_ASAP7_75t_SL g430 ( .A(n_384), .B(n_240), .Y(n_430) );
BUFx5_ASAP7_75t_L g431 ( .A(n_396), .Y(n_431) );
O2A1O1Ixp33_ASAP7_75t_SL g432 ( .A1(n_428), .A2(n_379), .B(n_387), .C(n_375), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_420), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_418), .B(n_377), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_410), .B(n_384), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_401), .B(n_384), .Y(n_436) );
BUFx4f_ASAP7_75t_L g437 ( .A(n_402), .Y(n_437) );
AOI21xp5_ASAP7_75t_L g438 ( .A1(n_428), .A2(n_387), .B(n_379), .Y(n_438) );
BUFx4f_ASAP7_75t_L g439 ( .A(n_402), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g440 ( .A1(n_424), .A2(n_388), .B(n_399), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_407), .A2(n_388), .B1(n_399), .B2(n_265), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_401), .B(n_399), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_404), .B(n_242), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_414), .B(n_245), .Y(n_444) );
OAI21xp5_ASAP7_75t_L g445 ( .A1(n_423), .A2(n_268), .B(n_248), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_415), .B(n_363), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_414), .B(n_250), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_411), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_419), .B(n_252), .Y(n_449) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_408), .Y(n_450) );
INVx4_ASAP7_75t_L g451 ( .A(n_408), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_400), .B(n_255), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_405), .B(n_358), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_412), .A2(n_271), .B(n_269), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_406), .B(n_256), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_416), .B(n_257), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_425), .B(n_261), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_406), .B(n_274), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_403), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_413), .A2(n_285), .B(n_277), .Y(n_460) );
CKINVDCx5p33_ASAP7_75t_R g461 ( .A(n_409), .Y(n_461) );
AOI21x1_ASAP7_75t_L g462 ( .A1(n_426), .A2(n_290), .B(n_288), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_417), .A2(n_294), .B(n_291), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_427), .A2(n_334), .B1(n_320), .B2(n_322), .Y(n_464) );
AND2x4_ASAP7_75t_L g465 ( .A(n_430), .B(n_296), .Y(n_465) );
NAND2x1p5_ASAP7_75t_L g466 ( .A(n_437), .B(n_358), .Y(n_466) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_450), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_448), .B(n_421), .Y(n_468) );
AND2x4_ASAP7_75t_L g469 ( .A(n_433), .B(n_426), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_459), .Y(n_470) );
OAI21xp5_ASAP7_75t_L g471 ( .A1(n_438), .A2(n_429), .B(n_422), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_441), .B(n_427), .Y(n_472) );
OAI21x1_ASAP7_75t_L g473 ( .A1(n_440), .A2(n_300), .B(n_298), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_450), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_432), .A2(n_306), .B(n_305), .Y(n_475) );
BUFx2_ASAP7_75t_L g476 ( .A(n_446), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_434), .B(n_427), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_445), .A2(n_324), .B(n_307), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_437), .Y(n_479) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_450), .Y(n_480) );
AO21x2_ASAP7_75t_L g481 ( .A1(n_445), .A2(n_330), .B(n_328), .Y(n_481) );
BUFx10_ASAP7_75t_L g482 ( .A(n_453), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_462), .Y(n_483) );
INVxp67_ASAP7_75t_L g484 ( .A(n_455), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_461), .B(n_431), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_436), .A2(n_340), .B(n_338), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_452), .A2(n_270), .B(n_262), .Y(n_487) );
OAI21x1_ASAP7_75t_L g488 ( .A1(n_463), .A2(n_297), .B(n_283), .Y(n_488) );
NAND2x1p5_ASAP7_75t_L g489 ( .A(n_439), .B(n_292), .Y(n_489) );
INVx4_ASAP7_75t_L g490 ( .A(n_451), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_457), .B(n_427), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_444), .A2(n_310), .B(n_308), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_442), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_458), .B(n_465), .Y(n_494) );
OAI21x1_ASAP7_75t_L g495 ( .A1(n_460), .A2(n_323), .B(n_313), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_447), .A2(n_339), .B(n_329), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_435), .Y(n_497) );
AO31x2_ASAP7_75t_L g498 ( .A1(n_458), .A2(n_431), .A3(n_342), .B(n_365), .Y(n_498) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_451), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_454), .A2(n_272), .B(n_264), .Y(n_500) );
NAND3xp33_ASAP7_75t_L g501 ( .A(n_464), .B(n_365), .C(n_342), .Y(n_501) );
OAI21x1_ASAP7_75t_L g502 ( .A1(n_456), .A2(n_431), .B(n_312), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_443), .B(n_6), .Y(n_503) );
OAI21x1_ASAP7_75t_L g504 ( .A1(n_449), .A2(n_431), .B(n_312), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_468), .B(n_465), .Y(n_505) );
BUFx3_ASAP7_75t_L g506 ( .A(n_466), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_468), .B(n_439), .Y(n_507) );
OAI21x1_ASAP7_75t_L g508 ( .A1(n_502), .A2(n_312), .B(n_260), .Y(n_508) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_471), .A2(n_369), .B(n_348), .Y(n_509) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_471), .A2(n_369), .B(n_348), .Y(n_510) );
OAI21x1_ASAP7_75t_SL g511 ( .A1(n_494), .A2(n_6), .B(n_7), .Y(n_511) );
INVx3_ASAP7_75t_SL g512 ( .A(n_482), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_483), .A2(n_369), .B(n_348), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_476), .B(n_7), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_470), .Y(n_515) );
OAI21x1_ASAP7_75t_L g516 ( .A1(n_473), .A2(n_260), .B(n_342), .Y(n_516) );
OAI21xp5_ASAP7_75t_L g517 ( .A1(n_478), .A2(n_486), .B(n_497), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_470), .Y(n_518) );
OAI21x1_ASAP7_75t_L g519 ( .A1(n_488), .A2(n_260), .B(n_365), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_469), .Y(n_520) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_475), .A2(n_276), .B(n_275), .Y(n_521) );
AOI222xp33_ASAP7_75t_L g522 ( .A1(n_469), .A2(n_293), .B1(n_327), .B2(n_260), .C1(n_333), .C2(n_331), .Y(n_522) );
OAI21x1_ASAP7_75t_SL g523 ( .A1(n_490), .A2(n_8), .B(n_9), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_484), .B(n_279), .Y(n_524) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_495), .A2(n_369), .B(n_348), .Y(n_525) );
OAI21x1_ASAP7_75t_L g526 ( .A1(n_474), .A2(n_365), .B(n_27), .Y(n_526) );
INVx2_ASAP7_75t_SL g527 ( .A(n_479), .Y(n_527) );
AND2x4_ASAP7_75t_L g528 ( .A(n_490), .B(n_9), .Y(n_528) );
INVx3_ASAP7_75t_L g529 ( .A(n_499), .Y(n_529) );
AO31x2_ASAP7_75t_L g530 ( .A1(n_492), .A2(n_376), .A3(n_11), .B(n_13), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_489), .B(n_10), .Y(n_531) );
OAI21x1_ASAP7_75t_L g532 ( .A1(n_496), .A2(n_29), .B(n_23), .Y(n_532) );
AO21x2_ASAP7_75t_L g533 ( .A1(n_481), .A2(n_376), .B(n_32), .Y(n_533) );
INVx4_ASAP7_75t_L g534 ( .A(n_499), .Y(n_534) );
OAI21x1_ASAP7_75t_L g535 ( .A1(n_501), .A2(n_34), .B(n_31), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_482), .B(n_280), .Y(n_536) );
INVx3_ASAP7_75t_L g537 ( .A(n_499), .Y(n_537) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_481), .A2(n_376), .B(n_36), .Y(n_538) );
OAI21x1_ASAP7_75t_L g539 ( .A1(n_501), .A2(n_38), .B(n_35), .Y(n_539) );
BUFx3_ASAP7_75t_L g540 ( .A(n_467), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_493), .Y(n_541) );
NOR2xp33_ASAP7_75t_R g542 ( .A(n_485), .B(n_11), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_498), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_491), .B(n_281), .Y(n_544) );
NAND2x1p5_ASAP7_75t_L g545 ( .A(n_467), .B(n_13), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_503), .Y(n_546) );
AO21x2_ASAP7_75t_L g547 ( .A1(n_487), .A2(n_376), .B(n_130), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_472), .A2(n_311), .B(n_335), .C(n_332), .Y(n_548) );
OAI21x1_ASAP7_75t_L g549 ( .A1(n_477), .A2(n_126), .B(n_227), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_480), .B(n_14), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_498), .Y(n_551) );
AO21x2_ASAP7_75t_L g552 ( .A1(n_498), .A2(n_124), .B(n_226), .Y(n_552) );
OA21x2_ASAP7_75t_L g553 ( .A1(n_500), .A2(n_336), .B(n_321), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_480), .B(n_15), .Y(n_554) );
OA332x1_ASAP7_75t_L g555 ( .A1(n_480), .A2(n_16), .A3(n_17), .B1(n_18), .B2(n_19), .B3(n_20), .C1(n_319), .C2(n_317), .Y(n_555) );
OAI21x1_ASAP7_75t_L g556 ( .A1(n_504), .A2(n_121), .B(n_223), .Y(n_556) );
CKINVDCx5p33_ASAP7_75t_R g557 ( .A(n_479), .Y(n_557) );
OAI21x1_ASAP7_75t_L g558 ( .A1(n_504), .A2(n_119), .B(n_222), .Y(n_558) );
OAI21x1_ASAP7_75t_SL g559 ( .A1(n_494), .A2(n_16), .B(n_17), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_468), .B(n_18), .Y(n_560) );
INVx6_ASAP7_75t_L g561 ( .A(n_482), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_515), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_541), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_507), .B(n_20), .Y(n_564) );
BUFx2_ASAP7_75t_L g565 ( .A(n_534), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_543), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_514), .B(n_309), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_551), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_518), .Y(n_569) );
INVx3_ASAP7_75t_L g570 ( .A(n_534), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_505), .A2(n_546), .B1(n_520), .B2(n_542), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_528), .B(n_284), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_528), .Y(n_573) );
OAI21xp5_ASAP7_75t_L g574 ( .A1(n_517), .A2(n_301), .B(n_299), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_508), .Y(n_575) );
OA21x2_ASAP7_75t_L g576 ( .A1(n_509), .A2(n_295), .B(n_302), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_560), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_560), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_505), .B(n_39), .Y(n_579) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_550), .Y(n_580) );
AO21x1_ASAP7_75t_L g581 ( .A1(n_545), .A2(n_40), .B(n_45), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_531), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_517), .A2(n_46), .B1(n_47), .B2(n_50), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_511), .A2(n_52), .B1(n_54), .B2(n_59), .Y(n_584) );
OA21x2_ASAP7_75t_L g585 ( .A1(n_509), .A2(n_61), .B(n_63), .Y(n_585) );
CKINVDCx11_ASAP7_75t_R g586 ( .A(n_512), .Y(n_586) );
AOI22xp33_ASAP7_75t_SL g587 ( .A1(n_523), .A2(n_64), .B1(n_65), .B2(n_66), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_550), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_554), .Y(n_589) );
BUFx2_ASAP7_75t_L g590 ( .A(n_529), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_559), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_561), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_545), .Y(n_593) );
INVx3_ASAP7_75t_L g594 ( .A(n_529), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_530), .Y(n_595) );
NAND2x1p5_ASAP7_75t_L g596 ( .A(n_537), .B(n_69), .Y(n_596) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_537), .Y(n_597) );
BUFx2_ASAP7_75t_L g598 ( .A(n_561), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_530), .Y(n_599) );
NAND2xp33_ASAP7_75t_SL g600 ( .A(n_555), .B(n_70), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_522), .B(n_71), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_522), .A2(n_72), .B1(n_73), .B2(n_77), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_544), .A2(n_80), .B1(n_81), .B2(n_84), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_527), .Y(n_604) );
BUFx2_ASAP7_75t_L g605 ( .A(n_557), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_553), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_553), .Y(n_607) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_540), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_521), .A2(n_85), .B1(n_86), .B2(n_88), .Y(n_609) );
OAI22xp33_ASAP7_75t_L g610 ( .A1(n_506), .A2(n_91), .B1(n_92), .B2(n_93), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_519), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_556), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_532), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_558), .Y(n_614) );
AO21x2_ASAP7_75t_L g615 ( .A1(n_510), .A2(n_95), .B(n_96), .Y(n_615) );
BUFx2_ASAP7_75t_L g616 ( .A(n_521), .Y(n_616) );
AO222x2_ASAP7_75t_L g617 ( .A1(n_536), .A2(n_221), .B1(n_104), .B2(n_106), .C1(n_108), .C2(n_109), .Y(n_617) );
CKINVDCx11_ASAP7_75t_R g618 ( .A(n_524), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_552), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_548), .B(n_103), .Y(n_620) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_510), .Y(n_621) );
AOI21xp33_ASAP7_75t_L g622 ( .A1(n_525), .A2(n_547), .B(n_538), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_549), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_516), .Y(n_624) );
AND2x4_ASAP7_75t_L g625 ( .A(n_525), .B(n_110), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_526), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_533), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_535), .Y(n_628) );
BUFx6f_ASAP7_75t_L g629 ( .A(n_539), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_533), .Y(n_630) );
OAI21x1_ASAP7_75t_L g631 ( .A1(n_513), .A2(n_111), .B(n_112), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_538), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_505), .A2(n_113), .B1(n_114), .B2(n_115), .Y(n_633) );
CKINVDCx5p33_ASAP7_75t_R g634 ( .A(n_506), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_541), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_541), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_541), .Y(n_637) );
INVx3_ASAP7_75t_L g638 ( .A(n_534), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_541), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_568), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_568), .Y(n_641) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_566), .Y(n_642) );
CKINVDCx10_ASAP7_75t_R g643 ( .A(n_586), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_582), .B(n_116), .Y(n_644) );
AND2x4_ASAP7_75t_L g645 ( .A(n_588), .B(n_117), .Y(n_645) );
OR2x6_ASAP7_75t_L g646 ( .A(n_625), .B(n_118), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_563), .Y(n_647) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_566), .Y(n_648) );
INVx2_ASAP7_75t_SL g649 ( .A(n_634), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_635), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_600), .A2(n_122), .B1(n_129), .B2(n_136), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_564), .B(n_141), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_636), .B(n_142), .Y(n_653) );
NOR2x1_ASAP7_75t_L g654 ( .A(n_570), .B(n_638), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_637), .B(n_639), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_562), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_617), .B(n_146), .Y(n_657) );
OR2x2_ASAP7_75t_L g658 ( .A(n_569), .B(n_147), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_604), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_573), .Y(n_660) );
AND2x4_ASAP7_75t_L g661 ( .A(n_580), .B(n_149), .Y(n_661) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_597), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_589), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_565), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_572), .B(n_150), .Y(n_665) );
OAI21xp5_ASAP7_75t_SL g666 ( .A1(n_571), .A2(n_152), .B(n_154), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_598), .B(n_155), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_608), .B(n_156), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_586), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_595), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_577), .B(n_217), .Y(n_671) );
AND2x4_ASAP7_75t_L g672 ( .A(n_593), .B(n_157), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_578), .B(n_215), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_608), .B(n_165), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_571), .B(n_167), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_599), .Y(n_676) );
BUFx3_ASAP7_75t_L g677 ( .A(n_570), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_638), .B(n_171), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_567), .B(n_601), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_600), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_592), .B(n_172), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_605), .B(n_590), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_597), .B(n_174), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_579), .B(n_175), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_594), .B(n_176), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_617), .A2(n_182), .B1(n_184), .B2(n_185), .Y(n_686) );
INVx2_ASAP7_75t_SL g687 ( .A(n_594), .Y(n_687) );
BUFx12f_ASAP7_75t_L g688 ( .A(n_618), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_618), .B(n_602), .Y(n_689) );
CKINVDCx5p33_ASAP7_75t_R g690 ( .A(n_603), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_602), .A2(n_188), .B1(n_190), .B2(n_191), .Y(n_691) );
AND2x2_ASAP7_75t_L g692 ( .A(n_574), .B(n_192), .Y(n_692) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_621), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_606), .B(n_195), .Y(n_694) );
BUFx2_ASAP7_75t_L g695 ( .A(n_596), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_607), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_575), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_591), .B(n_196), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_620), .B(n_197), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_576), .B(n_198), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_575), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_596), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_611), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_616), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_576), .B(n_207), .Y(n_705) );
INVx2_ASAP7_75t_SL g706 ( .A(n_625), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_581), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_621), .A2(n_210), .B1(n_211), .B2(n_212), .Y(n_708) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_619), .Y(n_709) );
INVx2_ASAP7_75t_SL g710 ( .A(n_576), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_587), .B(n_213), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_631), .Y(n_712) );
OR2x2_ASAP7_75t_L g713 ( .A(n_610), .B(n_584), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_610), .B(n_633), .Y(n_714) );
BUFx2_ASAP7_75t_L g715 ( .A(n_615), .Y(n_715) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_623), .Y(n_716) );
INVxp67_ASAP7_75t_L g717 ( .A(n_615), .Y(n_717) );
INVx3_ASAP7_75t_L g718 ( .A(n_585), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_611), .Y(n_719) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_642), .Y(n_720) );
BUFx2_ASAP7_75t_L g721 ( .A(n_677), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_647), .Y(n_722) );
INVx2_ASAP7_75t_SL g723 ( .A(n_643), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_650), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_682), .B(n_628), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_659), .B(n_584), .Y(n_726) );
AOI221xp5_ASAP7_75t_L g727 ( .A1(n_657), .A2(n_609), .B1(n_583), .B2(n_622), .C(n_613), .Y(n_727) );
NOR2xp67_ASAP7_75t_L g728 ( .A(n_688), .B(n_609), .Y(n_728) );
BUFx6f_ASAP7_75t_L g729 ( .A(n_677), .Y(n_729) );
AND2x4_ASAP7_75t_L g730 ( .A(n_706), .B(n_632), .Y(n_730) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_642), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_663), .B(n_585), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_686), .A2(n_583), .B1(n_612), .B2(n_614), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_686), .A2(n_612), .B1(n_614), .B2(n_624), .Y(n_734) );
NOR2x1p5_ASAP7_75t_L g735 ( .A(n_688), .B(n_629), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_657), .A2(n_629), .B1(n_627), .B2(n_630), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_664), .B(n_627), .Y(n_737) );
BUFx4f_ASAP7_75t_L g738 ( .A(n_646), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_655), .B(n_630), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_656), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_660), .Y(n_741) );
AND2x2_ASAP7_75t_SL g742 ( .A(n_695), .B(n_632), .Y(n_742) );
NOR2xp33_ASAP7_75t_SL g743 ( .A(n_669), .B(n_624), .Y(n_743) );
INVx2_ASAP7_75t_SL g744 ( .A(n_649), .Y(n_744) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_648), .Y(n_745) );
BUFx3_ASAP7_75t_L g746 ( .A(n_687), .Y(n_746) );
INVxp67_ASAP7_75t_SL g747 ( .A(n_648), .Y(n_747) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_662), .Y(n_748) );
BUFx2_ASAP7_75t_L g749 ( .A(n_654), .Y(n_749) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_662), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_689), .A2(n_626), .B1(n_629), .B2(n_679), .Y(n_751) );
INVxp33_ASAP7_75t_SL g752 ( .A(n_665), .Y(n_752) );
OR2x2_ASAP7_75t_L g753 ( .A(n_640), .B(n_641), .Y(n_753) );
AND2x2_ASAP7_75t_L g754 ( .A(n_706), .B(n_674), .Y(n_754) );
AND2x4_ASAP7_75t_L g755 ( .A(n_693), .B(n_676), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_696), .Y(n_756) );
AND2x2_ASAP7_75t_L g757 ( .A(n_668), .B(n_652), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_693), .B(n_683), .Y(n_758) );
BUFx2_ASAP7_75t_L g759 ( .A(n_646), .Y(n_759) );
AOI22xp33_ASAP7_75t_SL g760 ( .A1(n_713), .A2(n_714), .B1(n_646), .B2(n_690), .Y(n_760) );
OR2x2_ASAP7_75t_L g761 ( .A(n_658), .B(n_676), .Y(n_761) );
OR2x2_ASAP7_75t_L g762 ( .A(n_670), .B(n_704), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_670), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_644), .B(n_661), .Y(n_764) );
AND2x2_ASAP7_75t_L g765 ( .A(n_661), .B(n_678), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_709), .B(n_716), .Y(n_766) );
OR2x2_ASAP7_75t_L g767 ( .A(n_709), .B(n_716), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_661), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_702), .Y(n_769) );
OAI222xp33_ASAP7_75t_L g770 ( .A1(n_690), .A2(n_710), .B1(n_714), .B2(n_680), .C1(n_675), .C2(n_707), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_651), .A2(n_666), .B1(n_711), .B2(n_672), .Y(n_771) );
AND2x2_ASAP7_75t_L g772 ( .A(n_667), .B(n_645), .Y(n_772) );
OR2x2_ASAP7_75t_L g773 ( .A(n_720), .B(n_697), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_763), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_756), .Y(n_775) );
AOI221xp5_ASAP7_75t_L g776 ( .A1(n_760), .A2(n_651), .B1(n_671), .B2(n_673), .C(n_653), .Y(n_776) );
INVx2_ASAP7_75t_SL g777 ( .A(n_746), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_754), .B(n_698), .Y(n_778) );
AND2x4_ASAP7_75t_L g779 ( .A(n_735), .B(n_701), .Y(n_779) );
AND2x4_ASAP7_75t_L g780 ( .A(n_721), .B(n_701), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_725), .B(n_645), .Y(n_781) );
AND2x4_ASAP7_75t_SL g782 ( .A(n_729), .B(n_681), .Y(n_782) );
BUFx3_ASAP7_75t_L g783 ( .A(n_746), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_722), .B(n_645), .Y(n_784) );
AND2x2_ASAP7_75t_L g785 ( .A(n_758), .B(n_672), .Y(n_785) );
OR2x2_ASAP7_75t_L g786 ( .A(n_720), .B(n_697), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_731), .Y(n_787) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_731), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_724), .Y(n_789) );
OR2x2_ASAP7_75t_L g790 ( .A(n_745), .B(n_719), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_741), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_760), .B(n_703), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_740), .Y(n_793) );
OR2x2_ASAP7_75t_L g794 ( .A(n_745), .B(n_672), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_762), .Y(n_795) );
AND2x2_ASAP7_75t_L g796 ( .A(n_751), .B(n_715), .Y(n_796) );
AND2x4_ASAP7_75t_L g797 ( .A(n_759), .B(n_712), .Y(n_797) );
INVx2_ASAP7_75t_L g798 ( .A(n_753), .Y(n_798) );
NOR2xp33_ASAP7_75t_L g799 ( .A(n_752), .B(n_699), .Y(n_799) );
AND2x4_ASAP7_75t_L g800 ( .A(n_747), .B(n_718), .Y(n_800) );
INVxp33_ASAP7_75t_L g801 ( .A(n_738), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_726), .B(n_694), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_739), .B(n_705), .Y(n_803) );
NAND2xp67_ASAP7_75t_L g804 ( .A(n_772), .B(n_764), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_769), .B(n_700), .Y(n_805) );
OR2x2_ASAP7_75t_L g806 ( .A(n_767), .B(n_766), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_748), .Y(n_807) );
NAND2x1p5_ASAP7_75t_L g808 ( .A(n_738), .B(n_684), .Y(n_808) );
BUFx2_ASAP7_75t_SL g809 ( .A(n_723), .Y(n_809) );
AND2x4_ASAP7_75t_L g810 ( .A(n_747), .B(n_718), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_748), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_750), .Y(n_812) );
AND2x2_ASAP7_75t_L g813 ( .A(n_751), .B(n_717), .Y(n_813) );
NOR2xp33_ASAP7_75t_L g814 ( .A(n_804), .B(n_770), .Y(n_814) );
INVxp67_ASAP7_75t_L g815 ( .A(n_783), .Y(n_815) );
OR2x2_ASAP7_75t_L g816 ( .A(n_806), .B(n_750), .Y(n_816) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_788), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_775), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_795), .B(n_736), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_807), .B(n_736), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_775), .Y(n_821) );
OAI21xp5_ASAP7_75t_L g822 ( .A1(n_801), .A2(n_728), .B(n_770), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_811), .B(n_755), .Y(n_823) );
INVx2_ASAP7_75t_L g824 ( .A(n_773), .Y(n_824) );
AND2x2_ASAP7_75t_L g825 ( .A(n_781), .B(n_742), .Y(n_825) );
AND2x2_ASAP7_75t_L g826 ( .A(n_785), .B(n_742), .Y(n_826) );
AND2x2_ASAP7_75t_L g827 ( .A(n_798), .B(n_749), .Y(n_827) );
NAND2x1_ASAP7_75t_SL g828 ( .A(n_797), .B(n_765), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_777), .B(n_744), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_786), .Y(n_830) );
INVxp67_ASAP7_75t_L g831 ( .A(n_797), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_789), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_790), .Y(n_833) );
AND2x2_ASAP7_75t_L g834 ( .A(n_778), .B(n_755), .Y(n_834) );
NOR2xp33_ASAP7_75t_L g835 ( .A(n_791), .B(n_757), .Y(n_835) );
INVx2_ASAP7_75t_L g836 ( .A(n_774), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_793), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_817), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_817), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_836), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_816), .Y(n_841) );
OAI22xp33_ASAP7_75t_SL g842 ( .A1(n_815), .A2(n_808), .B1(n_743), .B2(n_799), .Y(n_842) );
AOI22xp5_ASAP7_75t_L g843 ( .A1(n_814), .A2(n_792), .B1(n_734), .B2(n_771), .Y(n_843) );
A2O1A1Ixp33_ASAP7_75t_L g844 ( .A1(n_814), .A2(n_809), .B(n_771), .C(n_782), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_819), .B(n_812), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_818), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_824), .B(n_787), .Y(n_847) );
NAND4xp25_ASAP7_75t_L g848 ( .A(n_822), .B(n_727), .C(n_776), .D(n_734), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g849 ( .A1(n_835), .A2(n_802), .B1(n_803), .B2(n_796), .Y(n_849) );
NAND2x1_ASAP7_75t_L g850 ( .A(n_829), .B(n_810), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_835), .A2(n_813), .B1(n_768), .B2(n_727), .Y(n_851) );
AOI31xp33_ASAP7_75t_L g852 ( .A1(n_844), .A2(n_829), .A3(n_831), .B(n_733), .Y(n_852) );
XOR2xp5_ASAP7_75t_L g853 ( .A(n_842), .B(n_827), .Y(n_853) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_848), .A2(n_843), .B1(n_851), .B2(n_849), .Y(n_854) );
OA21x2_ASAP7_75t_L g855 ( .A1(n_838), .A2(n_820), .B(n_832), .Y(n_855) );
XOR2x2_ASAP7_75t_L g856 ( .A(n_850), .B(n_828), .Y(n_856) );
NOR3xp33_ASAP7_75t_L g857 ( .A(n_839), .B(n_733), .C(n_691), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_846), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_841), .B(n_834), .Y(n_859) );
INVx3_ASAP7_75t_L g860 ( .A(n_856), .Y(n_860) );
OAI311xp33_ASAP7_75t_L g861 ( .A1(n_854), .A2(n_845), .A3(n_847), .B1(n_823), .C1(n_794), .Y(n_861) );
OAI221xp5_ASAP7_75t_SL g862 ( .A1(n_853), .A2(n_825), .B1(n_826), .B2(n_784), .C(n_805), .Y(n_862) );
NOR2xp33_ASAP7_75t_L g863 ( .A(n_852), .B(n_830), .Y(n_863) );
OAI322xp33_ASAP7_75t_L g864 ( .A1(n_858), .A2(n_821), .A3(n_837), .B1(n_833), .B2(n_840), .C1(n_793), .C2(n_836), .Y(n_864) );
NAND3xp33_ASAP7_75t_L g865 ( .A(n_863), .B(n_855), .C(n_857), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_864), .Y(n_866) );
NOR4xp25_ASAP7_75t_L g867 ( .A(n_860), .B(n_859), .C(n_855), .D(n_692), .Y(n_867) );
NOR3xp33_ASAP7_75t_L g868 ( .A(n_865), .B(n_862), .C(n_685), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_866), .Y(n_869) );
NOR3xp33_ASAP7_75t_SL g870 ( .A(n_869), .B(n_861), .C(n_867), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_870), .B(n_868), .Y(n_871) );
NAND2x1p5_ASAP7_75t_SL g872 ( .A(n_871), .B(n_708), .Y(n_872) );
AOI22xp5_ASAP7_75t_L g873 ( .A1(n_872), .A2(n_729), .B1(n_800), .B2(n_779), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_873), .Y(n_874) );
HB1xp67_ASAP7_75t_L g875 ( .A(n_874), .Y(n_875) );
XOR2xp5_ASAP7_75t_L g876 ( .A(n_875), .B(n_779), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_876), .Y(n_877) );
AND2x2_ASAP7_75t_L g878 ( .A(n_877), .B(n_780), .Y(n_878) );
OR2x6_ASAP7_75t_L g879 ( .A(n_878), .B(n_730), .Y(n_879) );
AOI211xp5_ASAP7_75t_L g880 ( .A1(n_879), .A2(n_732), .B(n_737), .C(n_761), .Y(n_880) );
endmodule