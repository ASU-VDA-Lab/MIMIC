module fake_netlist_6_182_n_1725 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1725);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1725;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_13),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_101),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_146),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_114),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_118),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_86),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_151),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_12),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_92),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_77),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_78),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_84),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_115),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_124),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_24),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_25),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_105),
.Y(n_173)
);

INVxp67_ASAP7_75t_SL g174 ( 
.A(n_127),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_1),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_60),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_119),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_120),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_113),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_58),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g181 ( 
.A(n_3),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_6),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_14),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_111),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_31),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_102),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_27),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_57),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_71),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_64),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_149),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_18),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_108),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_141),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_70),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_95),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_82),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_126),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_88),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_52),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_73),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_144),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_7),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_85),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_42),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_139),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_51),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_23),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_18),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_22),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_27),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_121),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_152),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_43),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_94),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_21),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_28),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_87),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_13),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_97),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_90),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_53),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_34),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_9),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_39),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_5),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g229 ( 
.A(n_72),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_122),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_68),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_130),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_42),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_15),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_30),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_25),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_49),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_62),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_5),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_74),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_137),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_28),
.Y(n_242)
);

BUFx8_ASAP7_75t_SL g243 ( 
.A(n_3),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_49),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_15),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_145),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_45),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_10),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_44),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_96),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_123),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_154),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_65),
.Y(n_253)
);

INVxp67_ASAP7_75t_SL g254 ( 
.A(n_155),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_44),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_32),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_4),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_36),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_134),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_24),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_19),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_80),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_104),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_54),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_59),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_66),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_107),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_30),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_21),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_98),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_39),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_103),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_55),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_32),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_35),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_106),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_133),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_46),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_135),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_45),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_148),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_75),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_129),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_131),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_91),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_31),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_138),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_8),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_69),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_43),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_76),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_50),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_40),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_0),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_116),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_8),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_6),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_147),
.Y(n_298)
);

BUFx10_ASAP7_75t_L g299 ( 
.A(n_48),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_4),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_125),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_38),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_79),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_67),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_12),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_83),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_23),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_47),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_19),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_167),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_191),
.Y(n_311)
);

NOR2xp67_ASAP7_75t_L g312 ( 
.A(n_239),
.B(n_0),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_176),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_243),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_195),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_198),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_181),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_214),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_200),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_184),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_181),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_169),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_220),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_177),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_219),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_253),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_181),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_181),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_285),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_215),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_295),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_181),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_181),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_205),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_217),
.Y(n_335)
);

INVxp33_ASAP7_75t_SL g336 ( 
.A(n_156),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_222),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_275),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_181),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_177),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_197),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_181),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_163),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_230),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_163),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_197),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_213),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_183),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_267),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_267),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_183),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_232),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_204),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_240),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_156),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_241),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_246),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_204),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_233),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_267),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_250),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_251),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_233),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_296),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_252),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_259),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_262),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_296),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_263),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_302),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_302),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_265),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_305),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_239),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_305),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_213),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_182),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_299),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_270),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_157),
.Y(n_380)
);

BUFx8_ASAP7_75t_L g381 ( 
.A(n_376),
.Y(n_381)
);

OAI21x1_ASAP7_75t_L g382 ( 
.A1(n_317),
.A2(n_196),
.B(n_164),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_355),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_317),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_321),
.B(n_190),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_349),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_312),
.B(n_229),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_349),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_377),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_349),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_347),
.B(n_190),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_321),
.B(n_238),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_350),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_376),
.B(n_244),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_350),
.Y(n_395)
);

BUFx8_ASAP7_75t_L g396 ( 
.A(n_322),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_350),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_310),
.B(n_235),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_360),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_360),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_327),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_360),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_327),
.B(n_238),
.Y(n_403)
);

OA21x2_ASAP7_75t_L g404 ( 
.A1(n_328),
.A2(n_172),
.B(n_171),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_328),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_332),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_332),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_333),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_333),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_339),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_339),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_342),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_342),
.B(n_196),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_343),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_324),
.B(n_244),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_343),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_345),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_345),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_348),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_348),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_351),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_351),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_353),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_353),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_338),
.A2(n_290),
.B1(n_236),
.B2(n_237),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_358),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_358),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_312),
.B(n_320),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_380),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_320),
.B(n_229),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_325),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_359),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_359),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_363),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_363),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_364),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_340),
.B(n_157),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_364),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_341),
.B(n_158),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_346),
.B(n_158),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_368),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_368),
.B(n_159),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_370),
.B(n_159),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_370),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_371),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_391),
.B(n_415),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_383),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_384),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_384),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_437),
.B(n_315),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_391),
.B(n_407),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_396),
.B(n_316),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_437),
.B(n_319),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_398),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_396),
.B(n_334),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_407),
.Y(n_456)
);

NAND2xp33_ASAP7_75t_L g457 ( 
.A(n_391),
.B(n_267),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_408),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_408),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_409),
.Y(n_460)
);

INVx8_ASAP7_75t_L g461 ( 
.A(n_385),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_335),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_409),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_404),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_383),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_384),
.Y(n_466)
);

AND2x6_ASAP7_75t_L g467 ( 
.A(n_385),
.B(n_267),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_411),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_384),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_R g470 ( 
.A(n_429),
.B(n_336),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_411),
.B(n_352),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_415),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_412),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_389),
.Y(n_474)
);

OAI22xp33_ASAP7_75t_L g475 ( 
.A1(n_431),
.A2(n_311),
.B1(n_318),
.B2(n_338),
.Y(n_475)
);

INVxp33_ASAP7_75t_L g476 ( 
.A(n_398),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_412),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_415),
.B(n_356),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_401),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_401),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_401),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_401),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_410),
.Y(n_483)
);

NAND2x1p5_ASAP7_75t_L g484 ( 
.A(n_404),
.B(n_161),
.Y(n_484)
);

INVx5_ASAP7_75t_L g485 ( 
.A(n_405),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_439),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_440),
.B(n_357),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_410),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_404),
.Y(n_489)
);

OR2x6_ASAP7_75t_L g490 ( 
.A(n_428),
.B(n_218),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_385),
.B(n_371),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_410),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_404),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_404),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_440),
.B(n_361),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_385),
.B(n_362),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_385),
.B(n_365),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_410),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_392),
.B(n_369),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_386),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_386),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_392),
.B(n_373),
.Y(n_502)
);

AND2x2_ASAP7_75t_SL g503 ( 
.A(n_404),
.B(n_306),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_396),
.B(n_372),
.Y(n_504)
);

NAND3xp33_ASAP7_75t_SL g505 ( 
.A(n_425),
.B(n_331),
.C(n_330),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_386),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_396),
.B(n_379),
.Y(n_507)
);

NAND3xp33_ASAP7_75t_L g508 ( 
.A(n_389),
.B(n_378),
.C(n_374),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_395),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_395),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_413),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_395),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_392),
.B(n_224),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_396),
.Y(n_514)
);

INVx4_ASAP7_75t_L g515 ( 
.A(n_405),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_402),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_392),
.B(n_264),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_402),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_392),
.B(n_291),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_405),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_398),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_403),
.B(n_373),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_428),
.B(n_337),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_403),
.B(n_375),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_405),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_405),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_403),
.B(n_375),
.Y(n_527)
);

OAI21xp33_ASAP7_75t_SL g528 ( 
.A1(n_387),
.A2(n_187),
.B(n_175),
.Y(n_528)
);

NOR2x1p5_ASAP7_75t_L g529 ( 
.A(n_394),
.B(n_314),
.Y(n_529)
);

OAI22xp33_ASAP7_75t_L g530 ( 
.A1(n_431),
.A2(n_256),
.B1(n_309),
.B2(n_192),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_413),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_430),
.A2(n_344),
.B1(n_367),
.B2(n_366),
.Y(n_532)
);

OR2x6_ASAP7_75t_L g533 ( 
.A(n_430),
.B(n_209),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_413),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_413),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_387),
.B(n_354),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_429),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_405),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_403),
.B(n_374),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_405),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_405),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_431),
.B(n_313),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_402),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_403),
.Y(n_544)
);

AND2x6_ASAP7_75t_L g545 ( 
.A(n_413),
.B(n_306),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_R g546 ( 
.A(n_429),
.B(n_160),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_406),
.B(n_174),
.Y(n_547)
);

INVxp33_ASAP7_75t_L g548 ( 
.A(n_425),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_406),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_406),
.B(n_254),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_381),
.B(n_442),
.Y(n_551)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_442),
.B(n_211),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_406),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_406),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_406),
.B(n_166),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_443),
.B(n_414),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_406),
.Y(n_557)
);

OAI22xp33_ASAP7_75t_L g558 ( 
.A1(n_443),
.A2(n_271),
.B1(n_206),
.B2(n_210),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_406),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_418),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_394),
.Y(n_561)
);

INVxp33_ASAP7_75t_L g562 ( 
.A(n_394),
.Y(n_562)
);

AND2x6_ASAP7_75t_L g563 ( 
.A(n_390),
.B(n_306),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_414),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_382),
.A2(n_234),
.B1(n_228),
.B2(n_227),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_417),
.B(n_180),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_419),
.B(n_323),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_390),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_381),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_418),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_381),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_418),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_417),
.B(n_188),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_382),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_381),
.B(n_229),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_419),
.B(n_420),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_420),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_381),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_390),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_418),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_390),
.Y(n_581)
);

INVx5_ASAP7_75t_L g582 ( 
.A(n_390),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_421),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_421),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_382),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_427),
.Y(n_586)
);

AND2x6_ASAP7_75t_L g587 ( 
.A(n_390),
.B(n_306),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_417),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_427),
.B(n_193),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_432),
.Y(n_590)
);

BUFx10_ASAP7_75t_L g591 ( 
.A(n_432),
.Y(n_591)
);

AND2x6_ASAP7_75t_L g592 ( 
.A(n_390),
.B(n_306),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_421),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_486),
.B(n_417),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_561),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_588),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_464),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_552),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_588),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_446),
.B(n_326),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_464),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_531),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_486),
.B(n_417),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_450),
.B(n_435),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_453),
.A2(n_487),
.B1(n_462),
.B2(n_446),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_562),
.B(n_160),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_556),
.B(n_435),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_556),
.B(n_435),
.Y(n_608)
);

A2O1A1Ixp33_ASAP7_75t_L g609 ( 
.A1(n_472),
.A2(n_287),
.B(n_199),
.C(n_201),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_472),
.B(n_162),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_468),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_531),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_470),
.Y(n_613)
);

NOR2xp67_ASAP7_75t_L g614 ( 
.A(n_536),
.B(n_433),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_468),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_544),
.B(n_194),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_544),
.B(n_435),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_451),
.B(n_435),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_534),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_562),
.B(n_162),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_534),
.Y(n_621)
);

INVxp33_ASAP7_75t_L g622 ( 
.A(n_447),
.Y(n_622)
);

OAI21xp5_ASAP7_75t_L g623 ( 
.A1(n_489),
.A2(n_400),
.B(n_388),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_522),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g625 ( 
.A(n_447),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_495),
.B(n_438),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_478),
.B(n_165),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_465),
.B(n_329),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_473),
.B(n_477),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_473),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_511),
.A2(n_203),
.B1(n_266),
.B2(n_281),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_477),
.B(n_438),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_456),
.B(n_438),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_535),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_493),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_458),
.B(n_438),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_465),
.B(n_299),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_471),
.B(n_165),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_461),
.Y(n_639)
);

INVx6_ASAP7_75t_L g640 ( 
.A(n_591),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_503),
.A2(n_231),
.B1(n_207),
.B2(n_208),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_591),
.B(n_539),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_459),
.B(n_438),
.Y(n_643)
);

AOI221x1_ASAP7_75t_L g644 ( 
.A1(n_574),
.A2(n_202),
.B1(n_212),
.B2(n_223),
.C(n_388),
.Y(n_644)
);

INVxp33_ASAP7_75t_L g645 ( 
.A(n_474),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_460),
.B(n_416),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_496),
.A2(n_276),
.B1(n_189),
.B2(n_186),
.Y(n_647)
);

O2A1O1Ixp33_ASAP7_75t_L g648 ( 
.A1(n_494),
.A2(n_225),
.B(n_245),
.C(n_247),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_474),
.B(n_299),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_490),
.A2(n_168),
.B1(n_170),
.B2(n_173),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_497),
.A2(n_277),
.B1(n_189),
.B2(n_186),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g652 ( 
.A(n_537),
.Y(n_652)
);

NAND3xp33_ASAP7_75t_L g653 ( 
.A(n_567),
.B(n_242),
.C(n_216),
.Y(n_653)
);

NOR3xp33_ASAP7_75t_L g654 ( 
.A(n_505),
.B(n_248),
.C(n_268),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_564),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_475),
.B(n_499),
.Y(n_656)
);

INVxp33_ASAP7_75t_L g657 ( 
.A(n_542),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_577),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_463),
.B(n_416),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_586),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_490),
.A2(n_298),
.B1(n_170),
.B2(n_173),
.Y(n_661)
);

NOR2x1p5_ASAP7_75t_L g662 ( 
.A(n_514),
.B(n_182),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_R g663 ( 
.A(n_514),
.B(n_168),
.Y(n_663)
);

A2O1A1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_552),
.A2(n_422),
.B(n_421),
.C(n_423),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_537),
.Y(n_665)
);

NOR2x1p5_ASAP7_75t_L g666 ( 
.A(n_508),
.B(n_185),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_539),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_503),
.B(n_416),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_484),
.B(n_178),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_SL g670 ( 
.A1(n_548),
.A2(n_294),
.B1(n_308),
.B2(n_307),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_522),
.B(n_416),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_L g672 ( 
.A1(n_574),
.A2(n_399),
.B(n_400),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_522),
.B(n_416),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_491),
.B(n_416),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_491),
.B(n_416),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_502),
.B(n_524),
.Y(n_676)
);

A2O1A1Ixp33_ASAP7_75t_L g677 ( 
.A1(n_513),
.A2(n_423),
.B(n_422),
.C(n_424),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_484),
.B(n_178),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_593),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_502),
.B(n_416),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_591),
.B(n_179),
.Y(n_681)
);

INVxp33_ASAP7_75t_L g682 ( 
.A(n_476),
.Y(n_682)
);

NAND2x1p5_ASAP7_75t_L g683 ( 
.A(n_569),
.B(n_433),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_593),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_524),
.B(n_422),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_560),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_558),
.B(n_179),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_517),
.B(n_272),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_461),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_484),
.B(n_272),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_527),
.B(n_422),
.Y(n_691)
);

AO22x2_ASAP7_75t_L g692 ( 
.A1(n_551),
.A2(n_280),
.B1(n_257),
.B2(n_278),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_527),
.B(n_423),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_490),
.B(n_273),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_590),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_560),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_519),
.B(n_273),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_457),
.B(n_423),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_530),
.B(n_276),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_533),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_533),
.B(n_277),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_457),
.B(n_424),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_576),
.B(n_424),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_570),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_570),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_589),
.B(n_585),
.Y(n_706)
);

A2O1A1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_585),
.A2(n_426),
.B(n_424),
.C(n_436),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_461),
.B(n_426),
.Y(n_708)
);

INVx8_ASAP7_75t_L g709 ( 
.A(n_533),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_547),
.B(n_279),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_589),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_565),
.A2(n_286),
.B1(n_249),
.B2(n_399),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_569),
.B(n_279),
.Y(n_713)
);

OR2x6_ASAP7_75t_L g714 ( 
.A(n_533),
.B(n_441),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_461),
.B(n_426),
.Y(n_715)
);

O2A1O1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_566),
.A2(n_445),
.B(n_444),
.C(n_434),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_526),
.B(n_426),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_526),
.B(n_436),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_526),
.B(n_436),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_572),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_572),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_589),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_500),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_529),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_548),
.A2(n_436),
.B1(n_284),
.B2(n_434),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_538),
.B(n_434),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_575),
.B(n_578),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_523),
.B(n_282),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_550),
.B(n_282),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_580),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_580),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_538),
.B(n_549),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_578),
.B(n_283),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_546),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_532),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_538),
.B(n_390),
.Y(n_736)
);

NOR2xp67_ASAP7_75t_L g737 ( 
.A(n_452),
.B(n_444),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_549),
.B(n_393),
.Y(n_738)
);

INVxp67_ASAP7_75t_SL g739 ( 
.A(n_525),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_528),
.B(n_283),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_549),
.B(n_393),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_583),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_554),
.B(n_445),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_467),
.A2(n_284),
.B1(n_274),
.B2(n_308),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_455),
.B(n_289),
.Y(n_745)
);

INVx5_ASAP7_75t_R g746 ( 
.A(n_476),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_554),
.B(n_553),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_583),
.Y(n_748)
);

OAI22xp33_ASAP7_75t_L g749 ( 
.A1(n_504),
.A2(n_185),
.B1(n_288),
.B2(n_307),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_555),
.B(n_289),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_525),
.B(n_304),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_525),
.B(n_304),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_525),
.B(n_303),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_525),
.B(n_303),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_541),
.B(n_301),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_584),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_554),
.B(n_397),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_584),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_557),
.B(n_397),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_507),
.B(n_301),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_L g761 ( 
.A(n_467),
.B(n_298),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_454),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_480),
.Y(n_763)
);

BUFx6f_ASAP7_75t_SL g764 ( 
.A(n_467),
.Y(n_764)
);

NOR2xp67_ASAP7_75t_L g765 ( 
.A(n_653),
.B(n_573),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_634),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_605),
.B(n_656),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_706),
.B(n_541),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_634),
.Y(n_769)
);

AND2x6_ASAP7_75t_SL g770 ( 
.A(n_746),
.B(n_521),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_598),
.B(n_571),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_639),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_602),
.Y(n_773)
);

OR2x2_ASAP7_75t_SL g774 ( 
.A(n_735),
.B(n_571),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_656),
.B(n_480),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_623),
.A2(n_515),
.B(n_540),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_611),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_612),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_638),
.B(n_481),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_625),
.B(n_559),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_641),
.A2(n_481),
.B1(n_488),
.B2(n_479),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_708),
.A2(n_515),
.B(n_540),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_639),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_619),
.Y(n_784)
);

A2O1A1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_694),
.A2(n_488),
.B(n_274),
.C(n_288),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_SL g786 ( 
.A1(n_694),
.A2(n_292),
.B1(n_293),
.B2(n_300),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_600),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_638),
.B(n_448),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_715),
.A2(n_540),
.B(n_515),
.Y(n_789)
);

OR2x2_ASAP7_75t_L g790 ( 
.A(n_595),
.B(n_292),
.Y(n_790)
);

OAI21xp5_ASAP7_75t_L g791 ( 
.A1(n_668),
.A2(n_448),
.B(n_449),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_627),
.B(n_449),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_615),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_637),
.B(n_293),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_627),
.B(n_466),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_635),
.A2(n_467),
.B1(n_545),
.B2(n_469),
.Y(n_796)
);

HB1xp67_ASAP7_75t_L g797 ( 
.A(n_596),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_599),
.B(n_520),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_607),
.B(n_466),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_621),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_672),
.A2(n_520),
.B(n_541),
.Y(n_801)
);

O2A1O1Ixp5_ASAP7_75t_L g802 ( 
.A1(n_707),
.A2(n_498),
.B(n_483),
.C(n_469),
.Y(n_802)
);

A2O1A1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_608),
.A2(n_297),
.B(n_300),
.C(n_482),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_604),
.A2(n_520),
.B(n_541),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_649),
.B(n_297),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_626),
.A2(n_541),
.B(n_485),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_674),
.A2(n_485),
.B(n_568),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_675),
.A2(n_485),
.B(n_568),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_680),
.A2(n_485),
.B(n_568),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_618),
.A2(n_485),
.B(n_579),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_640),
.Y(n_811)
);

OAI21xp5_ASAP7_75t_L g812 ( 
.A1(n_597),
.A2(n_498),
.B(n_483),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_706),
.B(n_579),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_739),
.A2(n_581),
.B(n_579),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_615),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_706),
.B(n_581),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_671),
.A2(n_581),
.B(n_482),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_657),
.B(n_479),
.Y(n_818)
);

NAND2xp33_ASAP7_75t_R g819 ( 
.A(n_762),
.B(n_221),
.Y(n_819)
);

OAI21x1_ASAP7_75t_L g820 ( 
.A1(n_736),
.A2(n_492),
.B(n_518),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_597),
.B(n_601),
.Y(n_821)
);

OAI21xp5_ASAP7_75t_L g822 ( 
.A1(n_601),
.A2(n_676),
.B(n_669),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_630),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_701),
.A2(n_492),
.B(n_260),
.C(n_258),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_614),
.B(n_467),
.Y(n_825)
);

AOI21x1_ASAP7_75t_L g826 ( 
.A1(n_594),
.A2(n_510),
.B(n_506),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_603),
.B(n_467),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_697),
.B(n_509),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_667),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_673),
.A2(n_582),
.B(n_518),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_697),
.B(n_629),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_630),
.B(n_506),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_635),
.B(n_509),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_743),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_685),
.A2(n_693),
.B(n_691),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_655),
.B(n_501),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_732),
.A2(n_582),
.B(n_543),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_658),
.B(n_501),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_617),
.A2(n_703),
.B(n_747),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_743),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_660),
.B(n_510),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_679),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_692),
.A2(n_545),
.B1(n_284),
.B2(n_587),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_695),
.B(n_512),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_711),
.B(n_512),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_738),
.A2(n_582),
.B(n_500),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_722),
.B(n_516),
.Y(n_847)
);

INVxp67_ASAP7_75t_L g848 ( 
.A(n_606),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_606),
.B(n_516),
.Y(n_849)
);

AOI21x1_ASAP7_75t_L g850 ( 
.A1(n_632),
.A2(n_543),
.B(n_582),
.Y(n_850)
);

A2O1A1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_701),
.A2(n_226),
.B(n_255),
.C(n_261),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_620),
.B(n_545),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_669),
.A2(n_545),
.B(n_587),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_679),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_SL g855 ( 
.A(n_613),
.B(n_269),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_622),
.B(n_645),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_624),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_620),
.B(n_545),
.Y(n_858)
);

INVx6_ASAP7_75t_L g859 ( 
.A(n_640),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_710),
.B(n_592),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_729),
.B(n_592),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_727),
.B(n_582),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_628),
.B(n_1),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_666),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_741),
.A2(n_757),
.B(n_690),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_763),
.B(n_592),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_678),
.A2(n_397),
.B(n_393),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_678),
.A2(n_397),
.B(n_393),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_642),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_728),
.B(n_592),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_684),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_690),
.A2(n_397),
.B(n_393),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_639),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_684),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_728),
.B(n_587),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_723),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_616),
.B(n_587),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_734),
.B(n_2),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_616),
.B(n_725),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_723),
.B(n_686),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_686),
.B(n_587),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_639),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_677),
.A2(n_587),
.B(n_563),
.Y(n_883)
);

OAI21xp33_ASAP7_75t_L g884 ( 
.A1(n_760),
.A2(n_661),
.B(n_650),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_726),
.A2(n_397),
.B(n_393),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_696),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_717),
.A2(n_718),
.B(n_719),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_665),
.Y(n_888)
);

AOI21x1_ASAP7_75t_L g889 ( 
.A1(n_646),
.A2(n_563),
.B(n_397),
.Y(n_889)
);

INVxp67_ASAP7_75t_L g890 ( 
.A(n_610),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_689),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_696),
.B(n_563),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_737),
.B(n_143),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_698),
.A2(n_397),
.B(n_393),
.Y(n_894)
);

AND2x6_ASAP7_75t_L g895 ( 
.A(n_727),
.B(n_393),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_702),
.A2(n_563),
.B(n_142),
.Y(n_896)
);

INVxp67_ASAP7_75t_L g897 ( 
.A(n_740),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_704),
.B(n_563),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_704),
.B(n_563),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_705),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_714),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_705),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_720),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_720),
.B(n_9),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_721),
.Y(n_905)
);

AO21x1_ASAP7_75t_L g906 ( 
.A1(n_751),
.A2(n_10),
.B(n_11),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_731),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_731),
.B(n_11),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_640),
.B(n_16),
.Y(n_909)
);

O2A1O1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_699),
.A2(n_17),
.B(n_20),
.C(n_22),
.Y(n_910)
);

O2A1O1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_687),
.A2(n_17),
.B(n_20),
.C(n_26),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_700),
.B(n_26),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_664),
.A2(n_643),
.B(n_633),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_759),
.A2(n_61),
.B(n_136),
.Y(n_914)
);

A2O1A1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_760),
.A2(n_29),
.B(n_33),
.C(n_34),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_727),
.B(n_56),
.Y(n_916)
);

AOI21xp33_ASAP7_75t_L g917 ( 
.A1(n_749),
.A2(n_29),
.B(n_33),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_742),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_742),
.Y(n_919)
);

OR2x2_ASAP7_75t_SL g920 ( 
.A(n_670),
.B(n_35),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_748),
.B(n_36),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_748),
.B(n_758),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_756),
.B(n_37),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_636),
.A2(n_89),
.B(n_132),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_756),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_758),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_659),
.A2(n_81),
.B(n_128),
.Y(n_927)
);

OAI321xp33_ASAP7_75t_L g928 ( 
.A1(n_740),
.A2(n_37),
.A3(n_38),
.B1(n_40),
.B2(n_41),
.C(n_46),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_730),
.B(n_692),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_692),
.B(n_41),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_750),
.B(n_688),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_689),
.A2(n_99),
.B(n_112),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_681),
.B(n_47),
.Y(n_933)
);

INVx4_ASAP7_75t_L g934 ( 
.A(n_689),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_652),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_750),
.B(n_48),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_648),
.A2(n_50),
.B(n_63),
.C(n_93),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_644),
.A2(n_752),
.B(n_753),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_689),
.B(n_100),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_716),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_744),
.A2(n_109),
.B1(n_110),
.B2(n_140),
.Y(n_941)
);

AOI21x1_ASAP7_75t_L g942 ( 
.A1(n_753),
.A2(n_754),
.B(n_755),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_754),
.B(n_755),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_631),
.B(n_647),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_793),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_772),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_787),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_767),
.A2(n_917),
.B(n_897),
.C(n_884),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_793),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_R g950 ( 
.A(n_888),
.B(n_724),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_769),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_R g952 ( 
.A(n_819),
.B(n_709),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_772),
.Y(n_953)
);

INVx3_ASAP7_75t_SL g954 ( 
.A(n_935),
.Y(n_954)
);

O2A1O1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_897),
.A2(n_745),
.B(n_651),
.C(n_713),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_815),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_848),
.B(n_709),
.Y(n_957)
);

NAND2x1p5_ASAP7_75t_L g958 ( 
.A(n_934),
.B(n_733),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_831),
.B(n_714),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_776),
.A2(n_835),
.B(n_801),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_772),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_L g962 ( 
.A1(n_944),
.A2(n_709),
.B1(n_654),
.B2(n_714),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_839),
.A2(n_683),
.B(n_761),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_848),
.B(n_712),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_941),
.A2(n_683),
.B1(n_764),
.B2(n_662),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_770),
.Y(n_966)
);

INVx4_ASAP7_75t_L g967 ( 
.A(n_772),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_775),
.B(n_779),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_782),
.A2(n_609),
.B(n_764),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_901),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_941),
.A2(n_663),
.B1(n_682),
.B2(n_786),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_856),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_856),
.B(n_890),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_789),
.A2(n_804),
.B(n_822),
.Y(n_974)
);

BUFx4f_ASAP7_75t_L g975 ( 
.A(n_859),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_821),
.A2(n_663),
.B(n_799),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_901),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_851),
.A2(n_785),
.B(n_915),
.C(n_824),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_821),
.A2(n_795),
.B(n_792),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_783),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_788),
.A2(n_865),
.B(n_816),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_794),
.B(n_805),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_771),
.Y(n_983)
);

INVx5_ASAP7_75t_L g984 ( 
.A(n_783),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_863),
.B(n_797),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_864),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_783),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_811),
.B(n_869),
.Y(n_988)
);

OAI22x1_ASAP7_75t_L g989 ( 
.A1(n_890),
.A2(n_869),
.B1(n_878),
.B2(n_912),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_813),
.A2(n_816),
.B(n_828),
.Y(n_990)
);

INVx4_ASAP7_75t_L g991 ( 
.A(n_783),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_823),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_855),
.B(n_829),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_829),
.B(n_797),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_813),
.A2(n_768),
.B(n_887),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_818),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_768),
.A2(n_875),
.B(n_870),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_777),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_873),
.Y(n_999)
);

INVx1_ASAP7_75t_SL g1000 ( 
.A(n_790),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_879),
.A2(n_943),
.B(n_931),
.C(n_938),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_851),
.A2(n_818),
.B(n_824),
.C(n_936),
.Y(n_1002)
);

BUFx12f_ASAP7_75t_L g1003 ( 
.A(n_774),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_786),
.B(n_933),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_857),
.B(n_834),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_791),
.A2(n_806),
.B(n_849),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_902),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_827),
.A2(n_833),
.B(n_913),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_814),
.A2(n_825),
.B(n_858),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_902),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_859),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_857),
.B(n_840),
.Y(n_1012)
);

O2A1O1Ixp5_ASAP7_75t_SL g1013 ( 
.A1(n_940),
.A2(n_939),
.B(n_916),
.C(n_929),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_773),
.B(n_778),
.Y(n_1014)
);

OAI221xp5_ASAP7_75t_L g1015 ( 
.A1(n_785),
.A2(n_819),
.B1(n_912),
.B2(n_930),
.C(n_915),
.Y(n_1015)
);

AOI21x1_ASAP7_75t_L g1016 ( 
.A1(n_850),
.A2(n_826),
.B(n_942),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_SL g1017 ( 
.A(n_934),
.B(n_873),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_873),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_843),
.A2(n_800),
.B1(n_784),
.B2(n_796),
.Y(n_1019)
);

INVx4_ASAP7_75t_L g1020 ( 
.A(n_873),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_766),
.B(n_918),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_918),
.B(n_919),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_919),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_882),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_842),
.Y(n_1025)
);

INVx5_ASAP7_75t_L g1026 ( 
.A(n_882),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_874),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_780),
.B(n_798),
.Y(n_1028)
);

NOR2xp67_ASAP7_75t_SL g1029 ( 
.A(n_928),
.B(n_882),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_852),
.A2(n_880),
.B(n_812),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_854),
.B(n_871),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_811),
.B(n_882),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_886),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_900),
.Y(n_1034)
);

NAND2xp33_ASAP7_75t_L g1035 ( 
.A(n_891),
.B(n_895),
.Y(n_1035)
);

OAI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_802),
.A2(n_803),
.B(n_817),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_802),
.A2(n_803),
.B(n_883),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_922),
.A2(n_862),
.B(n_810),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_780),
.B(n_859),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_765),
.A2(n_910),
.B(n_798),
.C(n_911),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_862),
.A2(n_832),
.B(n_809),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_891),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_860),
.A2(n_861),
.B(n_893),
.C(n_937),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_903),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_904),
.A2(n_923),
.B(n_921),
.C(n_908),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_905),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_925),
.B(n_926),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_891),
.B(n_909),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_907),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_891),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_876),
.B(n_838),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_893),
.B(n_876),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_836),
.B(n_844),
.Y(n_1053)
);

AO32x2_ASAP7_75t_L g1054 ( 
.A1(n_781),
.A2(n_906),
.A3(n_843),
.B1(n_820),
.B2(n_895),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_841),
.B(n_847),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_845),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_807),
.A2(n_808),
.B(n_853),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_881),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_939),
.A2(n_877),
.B(n_866),
.C(n_899),
.Y(n_1059)
);

BUFx2_ASAP7_75t_SL g1060 ( 
.A(n_895),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_892),
.A2(n_898),
.B(n_896),
.C(n_924),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_895),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_932),
.A2(n_927),
.B(n_914),
.C(n_830),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_920),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_867),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_894),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_837),
.A2(n_846),
.B(n_868),
.Y(n_1067)
);

NOR2x1_ASAP7_75t_L g1068 ( 
.A(n_872),
.B(n_885),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_889),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_811),
.B(n_901),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_811),
.B(n_901),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_848),
.B(n_605),
.Y(n_1072)
);

O2A1O1Ixp5_ASAP7_75t_L g1073 ( 
.A1(n_938),
.A2(n_551),
.B(n_831),
.C(n_767),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_776),
.A2(n_461),
.B(n_835),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_831),
.B(n_605),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_835),
.A2(n_767),
.B(n_839),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_772),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_848),
.B(n_605),
.Y(n_1078)
);

BUFx12f_ASAP7_75t_L g1079 ( 
.A(n_888),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_776),
.A2(n_461),
.B(n_835),
.Y(n_1080)
);

OAI22x1_ASAP7_75t_L g1081 ( 
.A1(n_890),
.A2(n_735),
.B1(n_425),
.B2(n_605),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_767),
.A2(n_917),
.B(n_897),
.C(n_884),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_848),
.B(n_605),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_884),
.A2(n_767),
.B1(n_605),
.B2(n_944),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_787),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_888),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_971),
.A2(n_1083),
.B(n_1072),
.C(n_1082),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1014),
.Y(n_1088)
);

AOI221x1_ASAP7_75t_L g1089 ( 
.A1(n_989),
.A2(n_971),
.B1(n_1040),
.B2(n_960),
.C(n_1002),
.Y(n_1089)
);

INVx4_ASAP7_75t_SL g1090 ( 
.A(n_954),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1014),
.Y(n_1091)
);

NAND2x1_ASAP7_75t_L g1092 ( 
.A(n_967),
.B(n_991),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1075),
.B(n_1084),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1027),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_975),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1078),
.B(n_996),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_985),
.B(n_982),
.Y(n_1097)
);

AO21x1_ASAP7_75t_L g1098 ( 
.A1(n_978),
.A2(n_948),
.B(n_968),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_955),
.A2(n_1073),
.B(n_1015),
.C(n_959),
.Y(n_1099)
);

NOR4xp25_ASAP7_75t_L g1100 ( 
.A(n_1004),
.B(n_1001),
.C(n_959),
.D(n_1028),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_1081),
.A2(n_973),
.B1(n_972),
.B2(n_964),
.Y(n_1101)
);

OR2x6_ASAP7_75t_L g1102 ( 
.A(n_1060),
.B(n_1079),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_947),
.B(n_1000),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_968),
.B(n_1056),
.Y(n_1104)
);

AO31x2_ASAP7_75t_L g1105 ( 
.A1(n_974),
.A2(n_1006),
.A3(n_1057),
.B(n_1043),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1074),
.A2(n_1080),
.B(n_1076),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_983),
.B(n_1000),
.Y(n_1107)
);

AOI221x1_ASAP7_75t_L g1108 ( 
.A1(n_1076),
.A2(n_1037),
.B1(n_997),
.B2(n_1009),
.C(n_1036),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_945),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_1016),
.A2(n_995),
.B(n_1067),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_949),
.Y(n_1111)
);

O2A1O1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_957),
.A2(n_947),
.B(n_964),
.C(n_965),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_993),
.B(n_1085),
.Y(n_1113)
);

AO31x2_ASAP7_75t_L g1114 ( 
.A1(n_963),
.A2(n_1038),
.A3(n_981),
.B(n_1041),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1013),
.A2(n_1008),
.B(n_1037),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1053),
.B(n_1039),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_976),
.A2(n_990),
.B(n_962),
.C(n_1045),
.Y(n_1117)
);

AO21x2_ASAP7_75t_L g1118 ( 
.A1(n_1036),
.A2(n_979),
.B(n_1030),
.Y(n_1118)
);

INVx1_ASAP7_75t_SL g1119 ( 
.A(n_970),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1055),
.A2(n_1061),
.B(n_1035),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_994),
.B(n_1086),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1055),
.A2(n_1063),
.B(n_1052),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_965),
.A2(n_1029),
.B1(n_1003),
.B2(n_1019),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1068),
.A2(n_1059),
.B(n_1066),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_969),
.A2(n_1017),
.B(n_1065),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_956),
.Y(n_1126)
);

AOI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1051),
.A2(n_1005),
.B(n_1012),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_975),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_1062),
.Y(n_1129)
);

INVx3_ASAP7_75t_SL g1130 ( 
.A(n_966),
.Y(n_1130)
);

BUFx4f_ASAP7_75t_L g1131 ( 
.A(n_1070),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1058),
.A2(n_1051),
.B(n_1031),
.Y(n_1132)
);

O2A1O1Ixp5_ASAP7_75t_L g1133 ( 
.A1(n_1048),
.A2(n_951),
.B(n_992),
.C(n_1049),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1047),
.A2(n_1022),
.B(n_1021),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_998),
.Y(n_1135)
);

OR2x6_ASAP7_75t_SL g1136 ( 
.A(n_1050),
.B(n_1034),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_1070),
.B(n_1071),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_1022),
.A2(n_1021),
.B(n_958),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1025),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_1011),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1017),
.A2(n_1069),
.B(n_1026),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1033),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_977),
.B(n_988),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_958),
.A2(n_1046),
.B(n_1044),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_SL g1145 ( 
.A1(n_1007),
.A2(n_1010),
.B(n_1023),
.C(n_1077),
.Y(n_1145)
);

AO31x2_ASAP7_75t_L g1146 ( 
.A1(n_1054),
.A2(n_1020),
.A3(n_991),
.B(n_967),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_988),
.B(n_1032),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_952),
.B(n_1071),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_999),
.A2(n_1018),
.B(n_1032),
.C(n_1062),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_946),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_946),
.Y(n_1151)
);

AOI221x1_ASAP7_75t_L g1152 ( 
.A1(n_1069),
.A2(n_1062),
.B1(n_1054),
.B2(n_1020),
.C(n_961),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1069),
.B(n_946),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_986),
.B(n_984),
.Y(n_1154)
);

AO31x2_ASAP7_75t_L g1155 ( 
.A1(n_1054),
.A2(n_1064),
.A3(n_1026),
.B(n_984),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_953),
.B(n_961),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_953),
.A2(n_961),
.B(n_980),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_953),
.A2(n_980),
.B(n_987),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_980),
.A2(n_987),
.B(n_1024),
.Y(n_1159)
);

INVx5_ASAP7_75t_L g1160 ( 
.A(n_987),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1024),
.A2(n_1042),
.B(n_950),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_1024),
.Y(n_1162)
);

INVx4_ASAP7_75t_L g1163 ( 
.A(n_1042),
.Y(n_1163)
);

AO31x2_ASAP7_75t_L g1164 ( 
.A1(n_960),
.A2(n_644),
.A3(n_974),
.B(n_1002),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_948),
.A2(n_605),
.B(n_767),
.C(n_884),
.Y(n_1165)
);

INVxp67_ASAP7_75t_L g1166 ( 
.A(n_973),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1074),
.A2(n_1080),
.B(n_1076),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1016),
.A2(n_820),
.B(n_995),
.Y(n_1168)
);

INVx2_ASAP7_75t_SL g1169 ( 
.A(n_954),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1016),
.A2(n_820),
.B(n_995),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1074),
.A2(n_1080),
.B(n_1076),
.Y(n_1171)
);

OAI21xp33_ASAP7_75t_L g1172 ( 
.A1(n_1084),
.A2(n_786),
.B(n_767),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1016),
.A2(n_820),
.B(n_995),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1074),
.A2(n_1080),
.B(n_1076),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_1075),
.B(n_542),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_954),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_945),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1016),
.A2(n_820),
.B(n_995),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1075),
.B(n_1078),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_948),
.A2(n_605),
.B(n_767),
.C(n_884),
.Y(n_1180)
);

AO31x2_ASAP7_75t_L g1181 ( 
.A1(n_960),
.A2(n_644),
.A3(n_974),
.B(n_1002),
.Y(n_1181)
);

OAI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1073),
.A2(n_1001),
.B(n_767),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1074),
.A2(n_1080),
.B(n_1076),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1014),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_975),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1014),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1084),
.A2(n_767),
.B1(n_605),
.B2(n_1075),
.Y(n_1187)
);

AO31x2_ASAP7_75t_L g1188 ( 
.A1(n_960),
.A2(n_644),
.A3(n_974),
.B(n_1002),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_972),
.B(n_310),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_985),
.B(n_600),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1075),
.B(n_767),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1016),
.A2(n_820),
.B(n_995),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1014),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_960),
.A2(n_644),
.A3(n_974),
.B(n_1002),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1062),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1075),
.B(n_767),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_985),
.B(n_600),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1016),
.A2(n_820),
.B(n_995),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1073),
.A2(n_1001),
.B(n_767),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1014),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1075),
.B(n_1078),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_945),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_985),
.B(n_600),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1014),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_985),
.B(n_600),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1014),
.Y(n_1206)
);

OAI21xp5_ASAP7_75t_SL g1207 ( 
.A1(n_1004),
.A2(n_786),
.B(n_605),
.Y(n_1207)
);

O2A1O1Ixp5_ASAP7_75t_L g1208 ( 
.A1(n_1076),
.A2(n_551),
.B(n_1073),
.C(n_963),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1014),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_945),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1074),
.A2(n_1080),
.B(n_1076),
.Y(n_1211)
);

BUFx2_ASAP7_75t_L g1212 ( 
.A(n_1085),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1075),
.B(n_1078),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1075),
.B(n_767),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1014),
.Y(n_1215)
);

BUFx2_ASAP7_75t_R g1216 ( 
.A(n_1086),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1014),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_SL g1218 ( 
.A(n_971),
.B(n_571),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1016),
.A2(n_820),
.B(n_995),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1084),
.A2(n_767),
.B1(n_605),
.B2(n_1075),
.Y(n_1220)
);

INVxp67_ASAP7_75t_L g1221 ( 
.A(n_973),
.Y(n_1221)
);

NOR2x1_ASAP7_75t_L g1222 ( 
.A(n_1011),
.B(n_811),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1074),
.A2(n_1080),
.B(n_1076),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_954),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1014),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1014),
.Y(n_1226)
);

BUFx8_ASAP7_75t_L g1227 ( 
.A(n_1095),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1218),
.A2(n_1172),
.B1(n_1187),
.B2(n_1220),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1094),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1179),
.A2(n_1201),
.B1(n_1213),
.B2(n_1175),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1104),
.A2(n_1226),
.B1(n_1088),
.B2(n_1225),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1126),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1216),
.Y(n_1233)
);

BUFx12f_ASAP7_75t_L g1234 ( 
.A(n_1095),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1146),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_1095),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_SL g1237 ( 
.A1(n_1121),
.A2(n_1113),
.B1(n_1221),
.B2(n_1166),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_SL g1238 ( 
.A1(n_1093),
.A2(n_1196),
.B1(n_1214),
.B2(n_1191),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1135),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_SL g1240 ( 
.A1(n_1093),
.A2(n_1196),
.B1(n_1214),
.B2(n_1191),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1123),
.A2(n_1203),
.B1(n_1205),
.B2(n_1197),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1123),
.A2(n_1190),
.B1(n_1189),
.B2(n_1098),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1101),
.A2(n_1097),
.B1(n_1116),
.B2(n_1096),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_SL g1244 ( 
.A1(n_1207),
.A2(n_1186),
.B1(n_1200),
.B2(n_1217),
.Y(n_1244)
);

INVx4_ASAP7_75t_L g1245 ( 
.A(n_1128),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1101),
.A2(n_1107),
.B1(n_1103),
.B2(n_1212),
.Y(n_1246)
);

CKINVDCx10_ASAP7_75t_R g1247 ( 
.A(n_1102),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_SL g1248 ( 
.A1(n_1165),
.A2(n_1180),
.B(n_1087),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_SL g1249 ( 
.A1(n_1207),
.A2(n_1193),
.B1(n_1215),
.B2(n_1091),
.Y(n_1249)
);

INVx6_ASAP7_75t_L g1250 ( 
.A(n_1128),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1128),
.Y(n_1251)
);

BUFx10_ASAP7_75t_L g1252 ( 
.A(n_1185),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1137),
.B(n_1147),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1185),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1104),
.B(n_1184),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1106),
.A2(n_1183),
.B(n_1223),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1131),
.Y(n_1257)
);

CKINVDCx11_ASAP7_75t_R g1258 ( 
.A(n_1130),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1204),
.A2(n_1206),
.B1(n_1209),
.B2(n_1136),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1119),
.A2(n_1143),
.B1(n_1137),
.B2(n_1102),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1119),
.A2(n_1102),
.B1(n_1122),
.B2(n_1147),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1182),
.A2(n_1199),
.B1(n_1148),
.B2(n_1142),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_1176),
.Y(n_1263)
);

INVx5_ASAP7_75t_L g1264 ( 
.A(n_1160),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1109),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1182),
.A2(n_1199),
.B1(n_1139),
.B2(n_1120),
.Y(n_1266)
);

OAI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1089),
.A2(n_1108),
.B1(n_1177),
.B2(n_1202),
.Y(n_1267)
);

CKINVDCx11_ASAP7_75t_R g1268 ( 
.A(n_1090),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_L g1269 ( 
.A(n_1154),
.Y(n_1269)
);

INVx2_ASAP7_75t_SL g1270 ( 
.A(n_1224),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_SL g1271 ( 
.A1(n_1115),
.A2(n_1125),
.B1(n_1118),
.B2(n_1100),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1210),
.A2(n_1115),
.B1(n_1169),
.B2(n_1118),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1222),
.A2(n_1154),
.B1(n_1144),
.B2(n_1124),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1132),
.A2(n_1150),
.B1(n_1151),
.B2(n_1195),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1129),
.A2(n_1195),
.B1(n_1211),
.B2(n_1171),
.Y(n_1275)
);

BUFx2_ASAP7_75t_SL g1276 ( 
.A(n_1140),
.Y(n_1276)
);

AOI22x1_ASAP7_75t_SL g1277 ( 
.A1(n_1129),
.A2(n_1163),
.B1(n_1090),
.B2(n_1112),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1133),
.Y(n_1278)
);

BUFx12f_ASAP7_75t_L g1279 ( 
.A(n_1163),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1167),
.A2(n_1174),
.B1(n_1138),
.B2(n_1162),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1134),
.Y(n_1281)
);

BUFx2_ASAP7_75t_R g1282 ( 
.A(n_1153),
.Y(n_1282)
);

CKINVDCx11_ASAP7_75t_R g1283 ( 
.A(n_1161),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1100),
.B(n_1099),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1153),
.A2(n_1159),
.B1(n_1156),
.B2(n_1141),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_SL g1286 ( 
.A1(n_1117),
.A2(n_1152),
.B(n_1127),
.Y(n_1286)
);

INVx8_ASAP7_75t_L g1287 ( 
.A(n_1092),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1110),
.A2(n_1158),
.B1(n_1157),
.B2(n_1219),
.Y(n_1288)
);

BUFx8_ASAP7_75t_L g1289 ( 
.A(n_1155),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1155),
.Y(n_1290)
);

INVx8_ASAP7_75t_L g1291 ( 
.A(n_1149),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1155),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1145),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1208),
.A2(n_1194),
.B1(n_1188),
.B2(n_1164),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1168),
.A2(n_1198),
.B1(n_1192),
.B2(n_1170),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1173),
.A2(n_1178),
.B1(n_1181),
.B2(n_1188),
.Y(n_1296)
);

BUFx4f_ASAP7_75t_L g1297 ( 
.A(n_1181),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1188),
.A2(n_1194),
.B1(n_1105),
.B2(n_1114),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1194),
.A2(n_1172),
.B1(n_1218),
.B2(n_767),
.Y(n_1299)
);

CKINVDCx20_ASAP7_75t_R g1300 ( 
.A(n_1105),
.Y(n_1300)
);

INVx1_ASAP7_75t_SL g1301 ( 
.A(n_1114),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1114),
.A2(n_1218),
.B1(n_1172),
.B2(n_884),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1218),
.A2(n_1172),
.B1(n_884),
.B2(n_971),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1218),
.A2(n_1172),
.B1(n_884),
.B2(n_971),
.Y(n_1304)
);

INVx6_ASAP7_75t_L g1305 ( 
.A(n_1095),
.Y(n_1305)
);

BUFx10_ASAP7_75t_L g1306 ( 
.A(n_1121),
.Y(n_1306)
);

OAI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1218),
.A2(n_1207),
.B1(n_1201),
.B2(n_1179),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1095),
.Y(n_1308)
);

OAI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1218),
.A2(n_1207),
.B1(n_1201),
.B2(n_1179),
.Y(n_1309)
);

BUFx10_ASAP7_75t_L g1310 ( 
.A(n_1121),
.Y(n_1310)
);

BUFx10_ASAP7_75t_L g1311 ( 
.A(n_1121),
.Y(n_1311)
);

BUFx8_ASAP7_75t_L g1312 ( 
.A(n_1095),
.Y(n_1312)
);

INVx1_ASAP7_75t_SL g1313 ( 
.A(n_1107),
.Y(n_1313)
);

INVx1_ASAP7_75t_SL g1314 ( 
.A(n_1107),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_SL g1315 ( 
.A1(n_1218),
.A2(n_1004),
.B1(n_542),
.B2(n_971),
.Y(n_1315)
);

CKINVDCx6p67_ASAP7_75t_R g1316 ( 
.A(n_1130),
.Y(n_1316)
);

INVx1_ASAP7_75t_SL g1317 ( 
.A(n_1107),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1094),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1094),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1107),
.Y(n_1320)
);

INVx2_ASAP7_75t_SL g1321 ( 
.A(n_1176),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1218),
.A2(n_1172),
.B1(n_884),
.B2(n_971),
.Y(n_1322)
);

INVx6_ASAP7_75t_L g1323 ( 
.A(n_1095),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_1216),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1094),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_SL g1326 ( 
.A1(n_1218),
.A2(n_1004),
.B1(n_542),
.B2(n_971),
.Y(n_1326)
);

OAI21xp33_ASAP7_75t_L g1327 ( 
.A1(n_1172),
.A2(n_605),
.B(n_884),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1111),
.Y(n_1328)
);

OAI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1218),
.A2(n_1207),
.B1(n_1201),
.B2(n_1179),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1097),
.B(n_1190),
.Y(n_1330)
);

INVx1_ASAP7_75t_SL g1331 ( 
.A(n_1107),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1094),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_SL g1333 ( 
.A1(n_1218),
.A2(n_1004),
.B1(n_542),
.B2(n_971),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1218),
.A2(n_1004),
.B1(n_542),
.B2(n_971),
.Y(n_1334)
);

INVx6_ASAP7_75t_L g1335 ( 
.A(n_1095),
.Y(n_1335)
);

INVx6_ASAP7_75t_L g1336 ( 
.A(n_1095),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1104),
.A2(n_767),
.B1(n_605),
.B2(n_1084),
.Y(n_1337)
);

INVx6_ASAP7_75t_L g1338 ( 
.A(n_1095),
.Y(n_1338)
);

BUFx12f_ASAP7_75t_L g1339 ( 
.A(n_1095),
.Y(n_1339)
);

AOI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1256),
.A2(n_1278),
.B(n_1284),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1290),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1238),
.B(n_1240),
.Y(n_1342)
);

INVx1_ASAP7_75t_SL g1343 ( 
.A(n_1313),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1281),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1315),
.A2(n_1333),
.B1(n_1326),
.B2(n_1334),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1292),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1298),
.B(n_1235),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1235),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1301),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1297),
.Y(n_1350)
);

INVx1_ASAP7_75t_SL g1351 ( 
.A(n_1314),
.Y(n_1351)
);

OR2x6_ASAP7_75t_L g1352 ( 
.A(n_1248),
.B(n_1256),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1238),
.B(n_1240),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1299),
.B(n_1228),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1231),
.B(n_1255),
.Y(n_1355)
);

INVx4_ASAP7_75t_L g1356 ( 
.A(n_1264),
.Y(n_1356)
);

INVx2_ASAP7_75t_SL g1357 ( 
.A(n_1289),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1300),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1289),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_1229),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_1264),
.Y(n_1361)
);

INVx1_ASAP7_75t_SL g1362 ( 
.A(n_1317),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1232),
.Y(n_1363)
);

AO21x2_ASAP7_75t_L g1364 ( 
.A1(n_1286),
.A2(n_1267),
.B(n_1307),
.Y(n_1364)
);

AOI221x1_ASAP7_75t_L g1365 ( 
.A1(n_1327),
.A2(n_1337),
.B1(n_1259),
.B2(n_1231),
.C(n_1239),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1299),
.B(n_1315),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1326),
.B(n_1333),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1318),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1319),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1325),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1295),
.A2(n_1296),
.B(n_1280),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1332),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1267),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1271),
.Y(n_1374)
);

AO21x2_ASAP7_75t_L g1375 ( 
.A1(n_1307),
.A2(n_1309),
.B(n_1329),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1271),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1288),
.A2(n_1275),
.B(n_1266),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1302),
.B(n_1243),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1294),
.Y(n_1379)
);

AO21x2_ASAP7_75t_L g1380 ( 
.A1(n_1309),
.A2(n_1329),
.B(n_1337),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1334),
.B(n_1244),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1294),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1328),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1265),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1272),
.Y(n_1385)
);

AOI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1259),
.A2(n_1253),
.B(n_1330),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1291),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1320),
.Y(n_1388)
);

OA21x2_ASAP7_75t_L g1389 ( 
.A1(n_1262),
.A2(n_1304),
.B(n_1303),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1322),
.A2(n_1230),
.B(n_1249),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1293),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1244),
.B(n_1249),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1331),
.Y(n_1393)
);

BUFx3_ASAP7_75t_L g1394 ( 
.A(n_1264),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1283),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1274),
.Y(n_1396)
);

BUFx4f_ASAP7_75t_SL g1397 ( 
.A(n_1234),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_1257),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1273),
.A2(n_1261),
.B(n_1285),
.Y(n_1399)
);

NOR3xp33_ASAP7_75t_L g1400 ( 
.A(n_1245),
.B(n_1268),
.C(n_1308),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1277),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1242),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1287),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1287),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1237),
.B(n_1311),
.Y(n_1405)
);

OR2x6_ASAP7_75t_L g1406 ( 
.A(n_1269),
.B(n_1276),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1241),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1246),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1260),
.B(n_1282),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1282),
.B(n_1308),
.Y(n_1410)
);

AO21x1_ASAP7_75t_SL g1411 ( 
.A1(n_1247),
.A2(n_1227),
.B(n_1312),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1358),
.B(n_1311),
.Y(n_1412)
);

INVxp67_ASAP7_75t_L g1413 ( 
.A(n_1393),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1358),
.B(n_1310),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1365),
.A2(n_1270),
.B(n_1321),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1358),
.B(n_1306),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1352),
.A2(n_1245),
.B(n_1254),
.Y(n_1417)
);

OAI211xp5_ASAP7_75t_L g1418 ( 
.A1(n_1390),
.A2(n_1258),
.B(n_1233),
.C(n_1324),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1350),
.B(n_1263),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1345),
.A2(n_1335),
.B1(n_1336),
.B2(n_1250),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1405),
.B(n_1306),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1367),
.A2(n_1310),
.B1(n_1316),
.B2(n_1339),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_SL g1423 ( 
.A(n_1395),
.B(n_1227),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_SL g1424 ( 
.A1(n_1390),
.A2(n_1312),
.B(n_1279),
.Y(n_1424)
);

A2O1A1Ixp33_ASAP7_75t_L g1425 ( 
.A1(n_1367),
.A2(n_1236),
.B(n_1254),
.C(n_1251),
.Y(n_1425)
);

O2A1O1Ixp33_ASAP7_75t_L g1426 ( 
.A1(n_1402),
.A2(n_1252),
.B(n_1250),
.C(n_1305),
.Y(n_1426)
);

NOR2x1_ASAP7_75t_SL g1427 ( 
.A(n_1352),
.B(n_1252),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_SL g1428 ( 
.A1(n_1395),
.A2(n_1323),
.B(n_1335),
.Y(n_1428)
);

A2O1A1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1381),
.A2(n_1323),
.B(n_1335),
.C(n_1336),
.Y(n_1429)
);

AO21x1_ASAP7_75t_L g1430 ( 
.A1(n_1391),
.A2(n_1336),
.B(n_1338),
.Y(n_1430)
);

NOR2x1_ASAP7_75t_SL g1431 ( 
.A(n_1352),
.B(n_1338),
.Y(n_1431)
);

NAND2x1p5_ASAP7_75t_L g1432 ( 
.A(n_1395),
.B(n_1403),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1359),
.B(n_1357),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1365),
.A2(n_1399),
.B(n_1352),
.Y(n_1434)
);

NAND4xp25_ASAP7_75t_L g1435 ( 
.A(n_1402),
.B(n_1408),
.C(n_1343),
.D(n_1362),
.Y(n_1435)
);

A2O1A1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1381),
.A2(n_1392),
.B(n_1342),
.C(n_1353),
.Y(n_1436)
);

NAND3xp33_ASAP7_75t_L g1437 ( 
.A(n_1408),
.B(n_1352),
.C(n_1353),
.Y(n_1437)
);

INVx5_ASAP7_75t_SL g1438 ( 
.A(n_1395),
.Y(n_1438)
);

INVx1_ASAP7_75t_SL g1439 ( 
.A(n_1343),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1360),
.B(n_1393),
.Y(n_1440)
);

A2O1A1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1392),
.A2(n_1342),
.B(n_1366),
.C(n_1378),
.Y(n_1441)
);

AO32x2_ASAP7_75t_L g1442 ( 
.A1(n_1357),
.A2(n_1361),
.A3(n_1356),
.B1(n_1360),
.B2(n_1382),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1351),
.B(n_1362),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1398),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1388),
.B(n_1410),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1410),
.B(n_1359),
.Y(n_1446)
);

AOI221xp5_ASAP7_75t_L g1447 ( 
.A1(n_1374),
.A2(n_1376),
.B1(n_1373),
.B2(n_1354),
.C(n_1385),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_SL g1448 ( 
.A1(n_1357),
.A2(n_1355),
.B(n_1359),
.Y(n_1448)
);

A2O1A1Ixp33_ASAP7_75t_L g1449 ( 
.A1(n_1378),
.A2(n_1399),
.B(n_1391),
.C(n_1409),
.Y(n_1449)
);

AOI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1389),
.A2(n_1375),
.B1(n_1407),
.B2(n_1380),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1363),
.B(n_1370),
.Y(n_1451)
);

NAND4xp25_ASAP7_75t_L g1452 ( 
.A(n_1373),
.B(n_1374),
.C(n_1376),
.D(n_1407),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1397),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1368),
.B(n_1369),
.Y(n_1454)
);

INVx5_ASAP7_75t_L g1455 ( 
.A(n_1395),
.Y(n_1455)
);

AO32x2_ASAP7_75t_L g1456 ( 
.A1(n_1361),
.A2(n_1356),
.A3(n_1379),
.B1(n_1382),
.B2(n_1372),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1384),
.B(n_1383),
.Y(n_1457)
);

NOR2x1_ASAP7_75t_SL g1458 ( 
.A(n_1386),
.B(n_1406),
.Y(n_1458)
);

NOR2xp67_ASAP7_75t_SL g1459 ( 
.A(n_1395),
.B(n_1403),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1341),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1341),
.Y(n_1461)
);

O2A1O1Ixp33_ASAP7_75t_SL g1462 ( 
.A1(n_1401),
.A2(n_1391),
.B(n_1404),
.C(n_1387),
.Y(n_1462)
);

AOI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1389),
.A2(n_1375),
.B1(n_1380),
.B2(n_1364),
.Y(n_1463)
);

OAI21xp33_ASAP7_75t_L g1464 ( 
.A1(n_1396),
.A2(n_1385),
.B(n_1386),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1454),
.B(n_1379),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1456),
.B(n_1340),
.Y(n_1466)
);

NAND2x1p5_ASAP7_75t_L g1467 ( 
.A(n_1463),
.B(n_1377),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1456),
.B(n_1364),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1456),
.B(n_1364),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1460),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1431),
.B(n_1344),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1461),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1442),
.B(n_1364),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1442),
.B(n_1451),
.Y(n_1474)
);

AOI21xp5_ASAP7_75t_SL g1475 ( 
.A1(n_1426),
.A2(n_1406),
.B(n_1389),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1442),
.B(n_1346),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_SL g1477 ( 
.A1(n_1437),
.A2(n_1375),
.B1(n_1380),
.B2(n_1389),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1457),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1448),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1458),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1440),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1413),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1434),
.B(n_1346),
.Y(n_1483)
);

NOR2x1_ASAP7_75t_L g1484 ( 
.A(n_1435),
.B(n_1415),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_1444),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1464),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1450),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1450),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1463),
.B(n_1347),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1415),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1470),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1470),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1474),
.B(n_1449),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1487),
.B(n_1348),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1474),
.B(n_1371),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1476),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1474),
.B(n_1371),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1472),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_1480),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1476),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1472),
.Y(n_1501)
);

INVx4_ASAP7_75t_L g1502 ( 
.A(n_1485),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1487),
.B(n_1348),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1473),
.B(n_1468),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1488),
.B(n_1439),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1476),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1471),
.B(n_1427),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1480),
.Y(n_1508)
);

INVxp67_ASAP7_75t_SL g1509 ( 
.A(n_1490),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1478),
.B(n_1443),
.Y(n_1510)
);

NAND3xp33_ASAP7_75t_L g1511 ( 
.A(n_1477),
.B(n_1441),
.C(n_1447),
.Y(n_1511)
);

NOR2x1_ASAP7_75t_SL g1512 ( 
.A(n_1468),
.B(n_1455),
.Y(n_1512)
);

NAND2x1_ASAP7_75t_L g1513 ( 
.A(n_1475),
.B(n_1459),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1486),
.B(n_1349),
.Y(n_1514)
);

AOI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1477),
.A2(n_1375),
.B1(n_1436),
.B2(n_1418),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1490),
.Y(n_1516)
);

NOR2x1_ASAP7_75t_SL g1517 ( 
.A(n_1493),
.B(n_1479),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1511),
.A2(n_1486),
.B1(n_1489),
.B2(n_1484),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1496),
.B(n_1489),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1496),
.B(n_1489),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1492),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1492),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1500),
.B(n_1469),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1500),
.B(n_1469),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1502),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1506),
.B(n_1467),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1491),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1493),
.B(n_1482),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1493),
.B(n_1482),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1502),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1512),
.B(n_1480),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1498),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_SL g1533 ( 
.A(n_1511),
.B(n_1455),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1506),
.B(n_1504),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1509),
.B(n_1481),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1498),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1505),
.B(n_1465),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1509),
.B(n_1465),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1514),
.B(n_1481),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1514),
.B(n_1484),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1504),
.B(n_1467),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1501),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1491),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1516),
.B(n_1483),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1501),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1516),
.B(n_1483),
.Y(n_1546)
);

INVx5_ASAP7_75t_L g1547 ( 
.A(n_1502),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1491),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1494),
.B(n_1483),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1491),
.Y(n_1550)
);

INVx3_ASAP7_75t_L g1551 ( 
.A(n_1502),
.Y(n_1551)
);

AND2x4_ASAP7_75t_SL g1552 ( 
.A(n_1502),
.B(n_1406),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1504),
.B(n_1467),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1494),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1554),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1517),
.B(n_1495),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1517),
.B(n_1512),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1534),
.B(n_1495),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1518),
.B(n_1495),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1554),
.Y(n_1560)
);

INVxp33_ASAP7_75t_L g1561 ( 
.A(n_1533),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1527),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1521),
.Y(n_1563)
);

AOI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1528),
.A2(n_1515),
.B1(n_1513),
.B2(n_1423),
.Y(n_1564)
);

NOR2xp67_ASAP7_75t_L g1565 ( 
.A(n_1547),
.B(n_1480),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1521),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1528),
.B(n_1497),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1540),
.B(n_1494),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1547),
.B(n_1507),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1540),
.B(n_1503),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1534),
.B(n_1497),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1534),
.B(n_1497),
.Y(n_1572)
);

INVx3_ASAP7_75t_L g1573 ( 
.A(n_1547),
.Y(n_1573)
);

INVxp67_ASAP7_75t_SL g1574 ( 
.A(n_1527),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1541),
.B(n_1507),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1541),
.B(n_1507),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1522),
.Y(n_1577)
);

INVx3_ASAP7_75t_R g1578 ( 
.A(n_1525),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1527),
.Y(n_1579)
);

INVxp67_ASAP7_75t_SL g1580 ( 
.A(n_1529),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1522),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1543),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1543),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1541),
.B(n_1507),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1529),
.B(n_1549),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1532),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1553),
.B(n_1526),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1543),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1548),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1553),
.B(n_1507),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_SL g1591 ( 
.A1(n_1519),
.A2(n_1467),
.B1(n_1466),
.B2(n_1515),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1549),
.B(n_1510),
.Y(n_1592)
);

NAND2x1_ASAP7_75t_L g1593 ( 
.A(n_1531),
.B(n_1499),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1532),
.Y(n_1594)
);

CKINVDCx16_ASAP7_75t_R g1595 ( 
.A(n_1525),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1547),
.B(n_1499),
.Y(n_1596)
);

AOI21xp33_ASAP7_75t_L g1597 ( 
.A1(n_1561),
.A2(n_1513),
.B(n_1547),
.Y(n_1597)
);

AOI221xp5_ASAP7_75t_L g1598 ( 
.A1(n_1591),
.A2(n_1526),
.B1(n_1546),
.B2(n_1544),
.C(n_1539),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1595),
.Y(n_1599)
);

O2A1O1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1559),
.A2(n_1513),
.B(n_1519),
.C(n_1520),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1563),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1556),
.B(n_1553),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1580),
.B(n_1539),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1563),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1562),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1559),
.B(n_1421),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1585),
.B(n_1537),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1591),
.B(n_1537),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1556),
.B(n_1531),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1562),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1566),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1566),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1585),
.B(n_1520),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1577),
.Y(n_1614)
);

NAND4xp25_ASAP7_75t_L g1615 ( 
.A(n_1564),
.B(n_1422),
.C(n_1429),
.D(n_1452),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1592),
.B(n_1567),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1564),
.B(n_1544),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1592),
.B(n_1519),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1595),
.B(n_1453),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1567),
.B(n_1546),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1568),
.B(n_1505),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1557),
.B(n_1531),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1578),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1568),
.B(n_1505),
.Y(n_1624)
);

INVxp67_ASAP7_75t_L g1625 ( 
.A(n_1555),
.Y(n_1625)
);

AOI211x1_ASAP7_75t_L g1626 ( 
.A1(n_1558),
.A2(n_1524),
.B(n_1523),
.C(n_1526),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1557),
.B(n_1531),
.Y(n_1627)
);

INVx2_ASAP7_75t_SL g1628 ( 
.A(n_1557),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1570),
.B(n_1535),
.Y(n_1629)
);

NAND4xp25_ASAP7_75t_L g1630 ( 
.A(n_1555),
.B(n_1400),
.C(n_1401),
.D(n_1416),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1570),
.B(n_1560),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1601),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1599),
.A2(n_1623),
.B1(n_1606),
.B2(n_1598),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1623),
.A2(n_1557),
.B1(n_1547),
.B2(n_1593),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1619),
.B(n_1609),
.Y(n_1635)
);

AOI221xp5_ASAP7_75t_SL g1636 ( 
.A1(n_1600),
.A2(n_1578),
.B1(n_1560),
.B2(n_1523),
.C(n_1524),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1604),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1606),
.B(n_1558),
.Y(n_1638)
);

NAND2xp33_ASAP7_75t_L g1639 ( 
.A(n_1617),
.B(n_1400),
.Y(n_1639)
);

OAI21xp33_ASAP7_75t_L g1640 ( 
.A1(n_1608),
.A2(n_1569),
.B(n_1587),
.Y(n_1640)
);

INVx2_ASAP7_75t_SL g1641 ( 
.A(n_1628),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1611),
.Y(n_1642)
);

OAI32xp33_ASAP7_75t_L g1643 ( 
.A1(n_1615),
.A2(n_1573),
.A3(n_1530),
.B1(n_1551),
.B2(n_1538),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1628),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1613),
.B(n_1571),
.Y(n_1645)
);

OAI221xp5_ASAP7_75t_L g1646 ( 
.A1(n_1597),
.A2(n_1630),
.B1(n_1619),
.B2(n_1625),
.C(n_1631),
.Y(n_1646)
);

AOI21xp33_ASAP7_75t_L g1647 ( 
.A1(n_1603),
.A2(n_1573),
.B(n_1593),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1622),
.B(n_1575),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1612),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1614),
.Y(n_1650)
);

INVxp67_ASAP7_75t_L g1651 ( 
.A(n_1622),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1629),
.B(n_1573),
.Y(n_1652)
);

AOI31xp33_ASAP7_75t_L g1653 ( 
.A1(n_1627),
.A2(n_1411),
.A3(n_1432),
.B(n_1569),
.Y(n_1653)
);

OAI32xp33_ASAP7_75t_L g1654 ( 
.A1(n_1618),
.A2(n_1573),
.A3(n_1551),
.B1(n_1530),
.B2(n_1538),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1626),
.B(n_1571),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1607),
.B(n_1569),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1633),
.A2(n_1547),
.B1(n_1616),
.B2(n_1621),
.Y(n_1657)
);

AOI31xp33_ASAP7_75t_L g1658 ( 
.A1(n_1636),
.A2(n_1627),
.A3(n_1411),
.B(n_1624),
.Y(n_1658)
);

OAI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1655),
.A2(n_1653),
.B1(n_1646),
.B2(n_1638),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1644),
.Y(n_1660)
);

OA21x2_ASAP7_75t_L g1661 ( 
.A1(n_1644),
.A2(n_1610),
.B(n_1605),
.Y(n_1661)
);

OAI21xp5_ASAP7_75t_SL g1662 ( 
.A1(n_1635),
.A2(n_1569),
.B(n_1609),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1639),
.A2(n_1531),
.B1(n_1596),
.B2(n_1602),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1632),
.Y(n_1664)
);

AOI22x1_ASAP7_75t_L g1665 ( 
.A1(n_1641),
.A2(n_1596),
.B1(n_1530),
.B2(n_1551),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1651),
.B(n_1602),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1639),
.B(n_1620),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1641),
.B(n_1572),
.Y(n_1668)
);

AOI222xp33_ASAP7_75t_L g1669 ( 
.A1(n_1640),
.A2(n_1643),
.B1(n_1652),
.B2(n_1650),
.C1(n_1649),
.C2(n_1642),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1652),
.B(n_1572),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1656),
.B(n_1587),
.Y(n_1671)
);

OAI31xp33_ASAP7_75t_SL g1672 ( 
.A1(n_1634),
.A2(n_1596),
.A3(n_1574),
.B(n_1584),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1656),
.B(n_1605),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1645),
.A2(n_1565),
.B1(n_1596),
.B2(n_1576),
.Y(n_1674)
);

OAI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1647),
.A2(n_1565),
.B1(n_1530),
.B2(n_1551),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1667),
.B(n_1659),
.Y(n_1676)
);

AO21x1_ASAP7_75t_L g1677 ( 
.A1(n_1658),
.A2(n_1637),
.B(n_1610),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1660),
.B(n_1648),
.Y(n_1678)
);

O2A1O1Ixp33_ASAP7_75t_L g1679 ( 
.A1(n_1657),
.A2(n_1654),
.B(n_1648),
.C(n_1574),
.Y(n_1679)
);

XNOR2xp5_ASAP7_75t_L g1680 ( 
.A(n_1671),
.B(n_1412),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1663),
.A2(n_1670),
.B1(n_1666),
.B2(n_1668),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1661),
.Y(n_1682)
);

O2A1O1Ixp33_ASAP7_75t_L g1683 ( 
.A1(n_1669),
.A2(n_1538),
.B(n_1535),
.C(n_1594),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1673),
.B(n_1577),
.Y(n_1684)
);

AOI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1662),
.A2(n_1674),
.B1(n_1675),
.B2(n_1664),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1682),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1678),
.B(n_1672),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1684),
.Y(n_1688)
);

NAND3xp33_ASAP7_75t_SL g1689 ( 
.A(n_1683),
.B(n_1665),
.C(n_1430),
.Y(n_1689)
);

NOR3xp33_ASAP7_75t_SL g1690 ( 
.A(n_1676),
.B(n_1661),
.C(n_1420),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1681),
.B(n_1445),
.Y(n_1691)
);

NOR3x1_ASAP7_75t_L g1692 ( 
.A(n_1677),
.B(n_1508),
.C(n_1499),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_SL g1693 ( 
.A(n_1679),
.B(n_1685),
.Y(n_1693)
);

OAI211xp5_ASAP7_75t_SL g1694 ( 
.A1(n_1680),
.A2(n_1562),
.B(n_1589),
.C(n_1588),
.Y(n_1694)
);

AOI221xp5_ASAP7_75t_L g1695 ( 
.A1(n_1693),
.A2(n_1582),
.B1(n_1579),
.B2(n_1589),
.C(n_1588),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1691),
.B(n_1575),
.Y(n_1696)
);

AOI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1689),
.A2(n_1583),
.B1(n_1579),
.B2(n_1589),
.C(n_1588),
.Y(n_1697)
);

NAND3xp33_ASAP7_75t_SL g1698 ( 
.A(n_1687),
.B(n_1414),
.C(n_1409),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1690),
.B(n_1576),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1698),
.A2(n_1694),
.B1(n_1688),
.B2(n_1686),
.Y(n_1700)
);

AOI211xp5_ASAP7_75t_L g1701 ( 
.A1(n_1699),
.A2(n_1692),
.B(n_1428),
.C(n_1446),
.Y(n_1701)
);

AOI221xp5_ASAP7_75t_SL g1702 ( 
.A1(n_1696),
.A2(n_1579),
.B1(n_1582),
.B2(n_1583),
.C(n_1594),
.Y(n_1702)
);

OAI322xp33_ASAP7_75t_L g1703 ( 
.A1(n_1695),
.A2(n_1583),
.A3(n_1582),
.B1(n_1581),
.B2(n_1586),
.C1(n_1524),
.C2(n_1523),
.Y(n_1703)
);

OAI221xp5_ASAP7_75t_L g1704 ( 
.A1(n_1697),
.A2(n_1586),
.B1(n_1581),
.B2(n_1479),
.C(n_1508),
.Y(n_1704)
);

OAI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1698),
.A2(n_1590),
.B(n_1584),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1700),
.B(n_1590),
.Y(n_1706)
);

NOR2x1_ASAP7_75t_L g1707 ( 
.A(n_1703),
.B(n_1479),
.Y(n_1707)
);

INVxp33_ASAP7_75t_SL g1708 ( 
.A(n_1705),
.Y(n_1708)
);

NOR3xp33_ASAP7_75t_SL g1709 ( 
.A(n_1704),
.B(n_1425),
.C(n_1417),
.Y(n_1709)
);

AO22x1_ASAP7_75t_L g1710 ( 
.A1(n_1701),
.A2(n_1479),
.B1(n_1508),
.B2(n_1419),
.Y(n_1710)
);

AOI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1708),
.A2(n_1702),
.B1(n_1433),
.B2(n_1552),
.Y(n_1711)
);

AOI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1706),
.A2(n_1552),
.B1(n_1419),
.B2(n_1438),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1707),
.Y(n_1713)
);

AOI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1713),
.A2(n_1711),
.B1(n_1712),
.B2(n_1710),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1714),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1715),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1716),
.A2(n_1709),
.B1(n_1548),
.B2(n_1550),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1717),
.A2(n_1424),
.B(n_1550),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1718),
.Y(n_1719)
);

NAND3xp33_ASAP7_75t_L g1720 ( 
.A(n_1719),
.B(n_1398),
.C(n_1550),
.Y(n_1720)
);

INVxp33_ASAP7_75t_SL g1721 ( 
.A(n_1719),
.Y(n_1721)
);

OAI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1720),
.A2(n_1548),
.B1(n_1536),
.B2(n_1545),
.Y(n_1722)
);

XNOR2xp5_ASAP7_75t_L g1723 ( 
.A(n_1721),
.B(n_1406),
.Y(n_1723)
);

AOI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1723),
.A2(n_1545),
.B1(n_1542),
.B2(n_1536),
.C(n_1462),
.Y(n_1724)
);

AOI211xp5_ASAP7_75t_L g1725 ( 
.A1(n_1724),
.A2(n_1722),
.B(n_1398),
.C(n_1394),
.Y(n_1725)
);


endmodule