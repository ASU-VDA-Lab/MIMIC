module fake_jpeg_25467_n_35 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_35);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_35;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_18;
wire n_20;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_32;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

AOI21xp33_ASAP7_75t_SL g17 ( 
.A1(n_12),
.A2(n_9),
.B(n_2),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_4),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_1),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_18),
.B(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_21),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_23),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_26),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_7),
.B1(n_14),
.B2(n_10),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_25),
.A2(n_8),
.B1(n_15),
.B2(n_16),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_17),
.B(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_30),
.B(n_24),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_30),
.B(n_2),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_1),
.Y(n_34)
);

AOI322xp5_ASAP7_75t_L g35 ( 
.A1(n_34),
.A2(n_3),
.A3(n_19),
.B1(n_27),
.B2(n_28),
.C1(n_22),
.C2(n_26),
.Y(n_35)
);


endmodule