module fake_jpeg_8254_n_321 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_8),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_18),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_35),
.Y(n_49)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_41),
.Y(n_53)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_25),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_51),
.B(n_59),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_21),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_56),
.Y(n_77)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_54),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_58),
.Y(n_82)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_40),
.B(n_25),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_61),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_21),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_62),
.B(n_73),
.C(n_28),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_64),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_49),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_65),
.B(n_63),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_35),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_83),
.Y(n_97)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_69),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_24),
.B1(n_27),
.B2(n_22),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_68),
.A2(n_72),
.B1(n_79),
.B2(n_87),
.Y(n_105)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_24),
.B1(n_27),
.B2(n_22),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_SL g73 ( 
.A1(n_56),
.A2(n_38),
.B(n_39),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_74),
.Y(n_90)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_76),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx4f_ASAP7_75t_SL g80 ( 
.A(n_53),
.Y(n_80)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

CKINVDCx12_ASAP7_75t_R g81 ( 
.A(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_43),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_24),
.B1(n_35),
.B2(n_22),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_84),
.A2(n_36),
.B1(n_28),
.B2(n_25),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_50),
.A2(n_24),
.B1(n_22),
.B2(n_32),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_73),
.B(n_78),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_89),
.A2(n_92),
.B1(n_95),
.B2(n_36),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_45),
.B(n_18),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_102),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_36),
.B1(n_42),
.B2(n_40),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_34),
.Y(n_100)
);

FAx1_ASAP7_75t_SL g118 ( 
.A(n_100),
.B(n_112),
.CI(n_114),
.CON(n_118),
.SN(n_118)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_106),
.Y(n_132)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_63),
.A2(n_34),
.B1(n_42),
.B2(n_45),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_107),
.A2(n_109),
.B1(n_36),
.B2(n_71),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_108),
.B(n_31),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_57),
.B1(n_64),
.B2(n_42),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_111),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_31),
.B1(n_23),
.B2(n_32),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_62),
.B(n_39),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_53),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_39),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_41),
.Y(n_121)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_117),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_125),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_121),
.B(n_105),
.Y(n_147)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_122),
.A2(n_133),
.B1(n_138),
.B2(n_140),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_123),
.A2(n_130),
.B(n_131),
.Y(n_163)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_128),
.Y(n_161)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_127),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_107),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_71),
.Y(n_129)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_97),
.Y(n_130)
);

NAND2xp33_ASAP7_75t_SL g131 ( 
.A(n_89),
.B(n_41),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_135),
.A2(n_137),
.B1(n_67),
.B2(n_69),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_136),
.A2(n_113),
.B1(n_106),
.B2(n_101),
.Y(n_153)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_141),
.A2(n_144),
.B(n_129),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_71),
.Y(n_142)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_81),
.C(n_70),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_115),
.C(n_92),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_99),
.B(n_16),
.Y(n_144)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_148),
.C(n_151),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_SL g207 ( 
.A(n_147),
.B(n_155),
.C(n_174),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_143),
.B(n_110),
.C(n_91),
.Y(n_148)
);

NAND3xp33_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_10),
.C(n_15),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_150),
.B(n_23),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_74),
.C(n_53),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_176),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_162),
.B1(n_173),
.B2(n_133),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_76),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_160),
.C(n_164),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_120),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_157),
.B(n_168),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_127),
.A2(n_119),
.B1(n_136),
.B2(n_123),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_158),
.A2(n_170),
.B1(n_142),
.B2(n_138),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_41),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_126),
.A2(n_86),
.B1(n_79),
.B2(n_54),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_118),
.B(n_41),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_41),
.C(n_47),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_121),
.C(n_39),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_132),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_169),
.B(n_177),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_131),
.A2(n_46),
.B1(n_86),
.B2(n_88),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_125),
.A2(n_46),
.B1(n_75),
.B2(n_16),
.Y(n_173)
);

BUFx12_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_180),
.A2(n_181),
.B1(n_26),
.B2(n_33),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_117),
.B1(n_116),
.B2(n_135),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_189),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_183),
.A2(n_197),
.B1(n_33),
.B2(n_26),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_121),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_192),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_195),
.Y(n_223)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_191),
.Y(n_210)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_146),
.B(n_138),
.C(n_124),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_163),
.A2(n_32),
.B(n_31),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_193),
.A2(n_200),
.B(n_171),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_140),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_148),
.B(n_39),
.C(n_38),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_39),
.C(n_38),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_198),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_170),
.A2(n_104),
.B1(n_23),
.B2(n_28),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_163),
.A2(n_18),
.B(n_104),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_203),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_38),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_167),
.Y(n_212)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

AND2x6_ASAP7_75t_L g204 ( 
.A(n_147),
.B(n_166),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_204),
.Y(n_231)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_176),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_145),
.A2(n_16),
.B1(n_30),
.B2(n_20),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_206),
.A2(n_33),
.B1(n_26),
.B2(n_20),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_218),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_212),
.B(n_19),
.C(n_17),
.Y(n_253)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

OA21x2_ASAP7_75t_L g215 ( 
.A1(n_207),
.A2(n_149),
.B(n_172),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_179),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_168),
.Y(n_221)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_221),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_224),
.A2(n_232),
.B1(n_187),
.B2(n_26),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_199),
.B(n_30),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_228),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_183),
.A2(n_176),
.B1(n_30),
.B2(n_20),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_226),
.A2(n_33),
.B1(n_20),
.B2(n_29),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_227),
.Y(n_235)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_186),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_29),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_206),
.B1(n_204),
.B2(n_196),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_212),
.B(n_185),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_234),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_186),
.Y(n_234)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_214),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_240),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_231),
.A2(n_192),
.B1(n_178),
.B2(n_195),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_238),
.A2(n_247),
.B1(n_221),
.B2(n_229),
.Y(n_255)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_223),
.B(n_202),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_249),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_245),
.A2(n_251),
.B1(n_228),
.B2(n_213),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_178),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_250),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_38),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_208),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_218),
.C(n_213),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_238),
.A2(n_231),
.B(n_210),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_254),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_255),
.A2(n_266),
.B1(n_19),
.B2(n_17),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_223),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_260),
.C(n_261),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_222),
.Y(n_258)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_258),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_259),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_209),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_219),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_265),
.C(n_270),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_215),
.C(n_211),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_243),
.A2(n_215),
.B1(n_222),
.B2(n_227),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_235),
.A2(n_252),
.B1(n_242),
.B2(n_240),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_267),
.B(n_269),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_242),
.A2(n_225),
.B1(n_19),
.B2(n_9),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_19),
.C(n_18),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_244),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_277),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_248),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_276),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_262),
.Y(n_275)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_275),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_239),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_261),
.A2(n_237),
.B(n_236),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_253),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_264),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_251),
.B(n_9),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_283),
.A2(n_6),
.B(n_11),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_284),
.A2(n_18),
.B1(n_17),
.B2(n_2),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_257),
.C(n_268),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_287),
.C(n_291),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_293),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_264),
.C(n_260),
.Y(n_287)
);

OAI321xp33_ASAP7_75t_L g289 ( 
.A1(n_282),
.A2(n_9),
.A3(n_15),
.B1(n_12),
.B2(n_11),
.C(n_4),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_289),
.A2(n_290),
.B1(n_284),
.B2(n_279),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_278),
.A2(n_7),
.B1(n_15),
.B2(n_11),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_19),
.C(n_1),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_0),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_274),
.A2(n_5),
.B(n_10),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_283),
.Y(n_297)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_297),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g299 ( 
.A(n_296),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_300),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_302),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_274),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_272),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_305),
.C(n_5),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_281),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_287),
.C(n_285),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_306),
.A2(n_308),
.B1(n_311),
.B2(n_6),
.Y(n_313)
);

OAI22xp33_ASAP7_75t_L g308 ( 
.A1(n_297),
.A2(n_292),
.B1(n_291),
.B2(n_2),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_307),
.A2(n_298),
.B1(n_303),
.B2(n_7),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_312),
.A2(n_313),
.B(n_314),
.Y(n_315)
);

AO21x1_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_4),
.B(n_7),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_309),
.A3(n_314),
.B1(n_310),
.B2(n_10),
.C1(n_17),
.C2(n_3),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_0),
.C(n_1),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_1),
.B(n_3),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_1),
.B(n_3),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_17),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_17),
.Y(n_321)
);


endmodule