module fake_jpeg_2509_n_227 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_227);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_9),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_0),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_6),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_13),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_13),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_2),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_86),
.Y(n_93)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_25),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_88),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_0),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_61),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_89),
.A2(n_62),
.B1(n_70),
.B2(n_74),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_87),
.B(n_74),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_90),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_89),
.A2(n_67),
.B1(n_73),
.B2(n_76),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_92),
.A2(n_62),
.B1(n_59),
.B2(n_60),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_57),
.B1(n_73),
.B2(n_78),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_100),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_57),
.B1(n_75),
.B2(n_78),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_65),
.B1(n_71),
.B2(n_58),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_58),
.B1(n_70),
.B2(n_79),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

CKINVDCx12_ASAP7_75t_R g105 ( 
.A(n_93),
.Y(n_105)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_86),
.B1(n_75),
.B2(n_77),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_111),
.B1(n_113),
.B2(n_120),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_88),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_115),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_102),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_55),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_77),
.B1(n_76),
.B2(n_68),
.Y(n_113)
);

BUFx16f_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_114),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_72),
.Y(n_115)
);

BUFx8_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_116),
.Y(n_127)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_97),
.A2(n_69),
.B1(n_79),
.B2(n_64),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_90),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_121),
.B(n_116),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_123),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_114),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_133),
.Y(n_156)
);

OAI32xp33_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_90),
.A3(n_95),
.B1(n_98),
.B2(n_64),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_132),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_90),
.B(n_81),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_11),
.B(n_12),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_80),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_107),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_138),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_1),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_135),
.B(n_139),
.Y(n_168)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_113),
.B(n_1),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_106),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_140),
.Y(n_147)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_110),
.B(n_3),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_151),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_131),
.A2(n_63),
.B(n_4),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_149),
.A2(n_157),
.B(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_138),
.A2(n_63),
.A3(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_152),
.A2(n_15),
.B(n_16),
.Y(n_187)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_154),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_54),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_137),
.A2(n_27),
.B1(n_51),
.B2(n_48),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_159),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_3),
.B1(n_5),
.B2(n_8),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_28),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_165),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_26),
.C(n_46),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_166),
.C(n_29),
.Y(n_174)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_23),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_142),
.B1(n_122),
.B2(n_144),
.Y(n_169)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_150),
.A2(n_164),
.B1(n_162),
.B2(n_147),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_170),
.A2(n_145),
.B1(n_152),
.B2(n_148),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_122),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_174),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_156),
.A2(n_11),
.B(n_12),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_185),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_154),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_184),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_30),
.C(n_45),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_182),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_52),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_14),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_161),
.A2(n_44),
.B(n_22),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_186),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_17),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_160),
.A2(n_15),
.B(n_16),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_188),
.B(n_157),
.Y(n_194)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_194),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_170),
.B(n_148),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_199),
.Y(n_207)
);

AO22x1_ASAP7_75t_L g196 ( 
.A1(n_183),
.A2(n_161),
.B1(n_18),
.B2(n_19),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_196),
.A2(n_176),
.B1(n_188),
.B2(n_181),
.Y(n_202)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_202),
.A2(n_204),
.B1(n_208),
.B2(n_203),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_195),
.A2(n_172),
.B1(n_179),
.B2(n_175),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_190),
.B(n_173),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_208),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_198),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_209),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_207),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_212),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_205),
.A2(n_198),
.B1(n_194),
.B2(n_185),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_213),
.A2(n_175),
.B1(n_201),
.B2(n_187),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_192),
.C(n_200),
.Y(n_215)
);

OAI21xp33_ASAP7_75t_L g217 ( 
.A1(n_215),
.A2(n_178),
.B(n_174),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_212),
.C(n_211),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_217),
.A2(n_215),
.B(n_182),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_220),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_218),
.C(n_214),
.Y(n_222)
);

AOI322xp5_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_35),
.A3(n_41),
.B1(n_39),
.B2(n_21),
.C1(n_34),
.C2(n_38),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_223),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_163),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_36),
.B1(n_18),
.B2(n_20),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_17),
.Y(n_227)
);


endmodule