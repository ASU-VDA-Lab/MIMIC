module fake_jpeg_20417_n_157 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_157);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_157;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_149;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_8),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_26),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_43),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_46),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_32),
.Y(n_75)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_79),
.Y(n_93)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_2),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_80),
.B(n_82),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_22),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_76),
.A2(n_50),
.B1(n_69),
.B2(n_65),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_66),
.B1(n_63),
.B2(n_64),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_62),
.B1(n_74),
.B2(n_72),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_53),
.B1(n_73),
.B2(n_75),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_55),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_67),
.B1(n_59),
.B2(n_71),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_94),
.A2(n_97),
.B1(n_101),
.B2(n_103),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_57),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_96),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_90),
.A2(n_85),
.B1(n_52),
.B2(n_67),
.Y(n_97)
);

NAND2x1_ASAP7_75t_SL g98 ( 
.A(n_91),
.B(n_52),
.Y(n_98)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_66),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_104),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_88),
.B1(n_70),
.B2(n_68),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_70),
.B1(n_68),
.B2(n_60),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_88),
.A2(n_60),
.B1(n_61),
.B2(n_51),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_105),
.A2(n_61),
.B1(n_3),
.B2(n_4),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_2),
.Y(n_122)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_109),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

AND2x6_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_25),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_110),
.B(n_120),
.Y(n_133)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_114),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_116),
.A2(n_9),
.B1(n_15),
.B2(n_17),
.Y(n_134)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_119),
.Y(n_129)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

AO21x2_ASAP7_75t_L g128 ( 
.A1(n_121),
.A2(n_30),
.B(n_45),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_112),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_124),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_5),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_125),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_29),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_131),
.B(n_134),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_128),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_33),
.C(n_12),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_132),
.A2(n_18),
.B(n_20),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_127),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_135),
.Y(n_144)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_136),
.A2(n_139),
.B1(n_142),
.B2(n_128),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_128),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_140),
.A2(n_138),
.B1(n_129),
.B2(n_133),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_145),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_145),
.B(n_137),
.C(n_141),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_147),
.A2(n_138),
.B1(n_144),
.B2(n_133),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_146),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_149),
.B(n_21),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_27),
.B1(n_34),
.B2(n_35),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_36),
.B(n_37),
.Y(n_152)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_38),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_154),
.A2(n_40),
.B(n_42),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_47),
.Y(n_157)
);


endmodule