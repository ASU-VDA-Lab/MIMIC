module fake_ariane_1524_n_242 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_38, n_2, n_18, n_32, n_28, n_37, n_9, n_11, n_34, n_26, n_3, n_14, n_0, n_36, n_33, n_19, n_30, n_39, n_40, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_242);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_38;
input n_2;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_11;
input n_34;
input n_26;
input n_3;
input n_14;
input n_0;
input n_36;
input n_33;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_242;

wire n_83;
wire n_233;
wire n_56;
wire n_60;
wire n_170;
wire n_190;
wire n_160;
wire n_64;
wire n_179;
wire n_180;
wire n_119;
wire n_124;
wire n_240;
wire n_167;
wire n_90;
wire n_195;
wire n_213;
wire n_47;
wire n_110;
wire n_153;
wire n_197;
wire n_221;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_158;
wire n_237;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_203;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_236;
wire n_205;
wire n_71;
wire n_109;
wire n_208;
wire n_96;
wire n_156;
wire n_209;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_187;
wire n_132;
wire n_62;
wire n_225;
wire n_147;
wire n_204;
wire n_235;
wire n_210;
wire n_200;
wire n_51;
wire n_166;
wire n_76;
wire n_218;
wire n_103;
wire n_79;
wire n_226;
wire n_46;
wire n_220;
wire n_84;
wire n_199;
wire n_91;
wire n_159;
wire n_107;
wire n_189;
wire n_72;
wire n_105;
wire n_128;
wire n_217;
wire n_44;
wire n_224;
wire n_82;
wire n_178;
wire n_42;
wire n_57;
wire n_131;
wire n_201;
wire n_229;
wire n_70;
wire n_222;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_214;
wire n_227;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_188;
wire n_185;
wire n_58;
wire n_65;
wire n_123;
wire n_212;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_198;
wire n_148;
wire n_232;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_228;
wire n_121;
wire n_93;
wire n_118;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_196;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_206;
wire n_207;
wire n_241;
wire n_238;
wire n_41;
wire n_219;
wire n_140;
wire n_55;
wire n_191;
wire n_151;
wire n_136;
wire n_231;
wire n_192;
wire n_80;
wire n_146;
wire n_234;
wire n_230;
wire n_211;
wire n_194;
wire n_97;
wire n_154;
wire n_215;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_202;
wire n_145;
wire n_78;
wire n_193;
wire n_59;
wire n_63;
wire n_99;
wire n_216;
wire n_155;
wire n_127;
wire n_239;
wire n_223;
wire n_54;

INVxp67_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_27),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVxp33_ASAP7_75t_SL g57 ( 
.A(n_3),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVxp33_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_4),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_13),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_11),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

INVxp33_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_28),
.Y(n_73)
);

INVxp33_ASAP7_75t_SL g74 ( 
.A(n_36),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_44),
.Y(n_76)
);

AND2x4_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_75),
.Y(n_77)
);

OAI21x1_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_19),
.B(n_32),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_0),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g83 ( 
.A(n_57),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_60),
.A2(n_0),
.B1(n_2),
.B2(n_6),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

BUFx8_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_56),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_61),
.Y(n_94)
);

NAND2x1p5_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_7),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_49),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_54),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_2),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_59),
.B(n_71),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_41),
.B(n_12),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_76),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_105),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

INVxp33_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

AND2x6_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_104),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_80),
.A2(n_61),
.B1(n_73),
.B2(n_71),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_97),
.B(n_74),
.Y(n_118)
);

AND2x4_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_46),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_94),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_94),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_98),
.B(n_67),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_73),
.Y(n_129)
);

AO22x2_ASAP7_75t_L g130 ( 
.A1(n_80),
.A2(n_24),
.B1(n_30),
.B2(n_34),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

NAND2x1p5_ASAP7_75t_L g132 ( 
.A(n_87),
.B(n_93),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_77),
.B(n_106),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_83),
.Y(n_135)
);

AO22x2_ASAP7_75t_L g136 ( 
.A1(n_92),
.A2(n_104),
.B1(n_84),
.B2(n_96),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_82),
.B(n_89),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_122),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_135),
.Y(n_140)
);

NAND2x2_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_99),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_109),
.B(n_82),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_87),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_91),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_102),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_103),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_103),
.Y(n_154)
);

NOR2xp67_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_107),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_101),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

NOR2x1p5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_86),
.Y(n_158)
);

BUFx8_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

NOR3xp33_ASAP7_75t_SL g160 ( 
.A(n_118),
.B(n_126),
.C(n_113),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_108),
.Y(n_162)
);

INVxp67_ASAP7_75t_SL g163 ( 
.A(n_121),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

AND2x4_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_110),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

CKINVDCx11_ASAP7_75t_R g169 ( 
.A(n_141),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_136),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

AND2x4_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_117),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_140),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

NAND2xp33_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_130),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_145),
.A2(n_151),
.B(n_152),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_155),
.B(n_95),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_164),
.A2(n_130),
.B1(n_136),
.B2(n_116),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_164),
.A2(n_95),
.B1(n_132),
.B2(n_131),
.Y(n_189)
);

AO21x2_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_78),
.B(n_116),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_159),
.A2(n_120),
.B1(n_124),
.B2(n_116),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_171),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_170),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_184),
.A2(n_149),
.B(n_150),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_178),
.A2(n_158),
.B1(n_139),
.B2(n_120),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_170),
.B(n_150),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_178),
.A2(n_124),
.B1(n_141),
.B2(n_147),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_173),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_116),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_167),
.A2(n_163),
.B(n_150),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_187),
.A2(n_149),
.B1(n_146),
.B2(n_101),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_101),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_175),
.A2(n_157),
.B1(n_144),
.B2(n_121),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_172),
.A2(n_144),
.B1(n_188),
.B2(n_182),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_192),
.A2(n_183),
.B1(n_189),
.B2(n_172),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_191),
.A2(n_144),
.B1(n_174),
.B2(n_166),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_165),
.A2(n_186),
.B1(n_177),
.B2(n_168),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_173),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_180),
.Y(n_211)
);

OAI21x1_ASAP7_75t_L g212 ( 
.A1(n_195),
.A2(n_174),
.B(n_166),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

OAI21x1_ASAP7_75t_L g214 ( 
.A1(n_202),
.A2(n_181),
.B(n_168),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_194),
.A2(n_176),
.B1(n_165),
.B2(n_186),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_196),
.A2(n_165),
.B1(n_181),
.B2(n_173),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_204),
.A2(n_173),
.B1(n_168),
.B2(n_185),
.Y(n_217)
);

OA21x2_ASAP7_75t_L g218 ( 
.A1(n_209),
.A2(n_190),
.B(n_185),
.Y(n_218)
);

AOI221x1_ASAP7_75t_SL g219 ( 
.A1(n_194),
.A2(n_169),
.B1(n_185),
.B2(n_190),
.C(n_198),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_201),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_207),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_217),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_215),
.A2(n_206),
.B1(n_197),
.B2(n_203),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_212),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_220),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_218),
.Y(n_227)
);

OAI221xp5_ASAP7_75t_L g228 ( 
.A1(n_224),
.A2(n_219),
.B1(n_216),
.B2(n_217),
.C(n_197),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_227),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_227),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_230),
.A2(n_228),
.B(n_222),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_229),
.Y(n_232)
);

NOR3x1_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_169),
.C(n_200),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_233),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_234),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_235),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_236),
.A2(n_231),
.B1(n_222),
.B2(n_225),
.Y(n_237)
);

NOR3xp33_ASAP7_75t_SL g238 ( 
.A(n_237),
.B(n_216),
.C(n_210),
.Y(n_238)
);

NOR3xp33_ASAP7_75t_L g239 ( 
.A(n_238),
.B(n_210),
.C(n_200),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_205),
.Y(n_240)
);

AOI222xp33_ASAP7_75t_L g241 ( 
.A1(n_240),
.A2(n_208),
.B1(n_210),
.B2(n_218),
.C1(n_223),
.C2(n_237),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_241),
.A2(n_223),
.B(n_218),
.Y(n_242)
);


endmodule