module real_aes_2206_n_3 (n_0, n_2, n_1, n_3);
input n_0;
input n_2;
input n_1;
output n_3;
wire n_4;
wire n_5;
wire n_7;
wire n_8;
wire n_6;
wire n_9;
wire n_10;
wire n_11;
CKINVDCx20_ASAP7_75t_R g5 ( .A(n_0), .Y(n_5) );
NAND2xp5_ASAP7_75t_L g7 ( .A(n_0), .B(n_8), .Y(n_7) );
AOI21xp5_ASAP7_75t_L g4 ( .A1(n_1), .A2(n_5), .B(n_6), .Y(n_4) );
CKINVDCx16_ASAP7_75t_R g8 ( .A(n_1), .Y(n_8) );
CKINVDCx16_ASAP7_75t_R g10 ( .A(n_2), .Y(n_10) );
AOI22xp33_ASAP7_75t_SL g3 ( .A1(n_4), .A2(n_6), .B1(n_9), .B2(n_11), .Y(n_3) );
INVx2_ASAP7_75t_L g6 ( .A(n_7), .Y(n_6) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_9), .Y(n_11) );
CKINVDCx16_ASAP7_75t_R g9 ( .A(n_10), .Y(n_9) );
endmodule