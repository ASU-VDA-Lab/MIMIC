module real_jpeg_4219_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_1),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_2),
.A2(n_21),
.B1(n_27),
.B2(n_28),
.Y(n_20)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_4),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_5),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_5),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_5),
.A2(n_44),
.B1(n_88),
.B2(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_5),
.A2(n_88),
.B1(n_215),
.B2(n_218),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_6),
.A2(n_94),
.B1(n_97),
.B2(n_98),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_6),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_6),
.A2(n_98),
.B1(n_182),
.B2(n_184),
.Y(n_181)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_8),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_9),
.A2(n_35),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_9),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_10),
.B(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_10),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_10),
.A2(n_119),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_10),
.B(n_176),
.C(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_10),
.B(n_111),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_10),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_10),
.B(n_92),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_11),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_11),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_12),
.A2(n_22),
.B1(n_39),
.B2(n_42),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_12),
.A2(n_42),
.B1(n_123),
.B2(n_125),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_12),
.A2(n_42),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_161),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_159),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_127),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_16),
.B(n_127),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_65),
.C(n_99),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_17),
.B(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_43),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_18),
.B(n_43),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_30),
.B(n_32),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_20),
.A2(n_33),
.B1(n_154),
.B2(n_157),
.Y(n_153)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx4_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_26),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_30),
.Y(n_221)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_31),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_31),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_32),
.A2(n_214),
.B(n_220),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_38),
.Y(n_32)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_33),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_33),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_36),
.Y(n_155)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_37),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_37),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_38),
.B(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_41),
.Y(n_178)
);

AOI32xp33_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_49),
.A3(n_51),
.B1(n_55),
.B2(n_59),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_47),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_47),
.Y(n_151)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_48),
.Y(n_124)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_48),
.Y(n_150)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_49),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_50),
.Y(n_174)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_57),
.A2(n_104),
.B1(n_107),
.B2(n_108),
.Y(n_103)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_62),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AO22x2_ASAP7_75t_L g111 ( 
.A1(n_63),
.A2(n_79),
.B1(n_112),
.B2(n_114),
.Y(n_111)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_65),
.A2(n_99),
.B1(n_100),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_65),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_86),
.B1(n_91),
.B2(n_93),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_66),
.A2(n_93),
.B(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_66),
.A2(n_131),
.B(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_67),
.B(n_132),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_80),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_73),
.B1(n_76),
.B2(n_79),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_72),
.Y(n_168)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_80),
.A2(n_86),
.B(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_84),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g219 ( 
.A(n_84),
.Y(n_219)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_92),
.B(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_115),
.B(n_121),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_111),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_119),
.B(n_120),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_146),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_119),
.A2(n_188),
.B(n_189),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_126),
.A2(n_139),
.B(n_142),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_137),
.B2(n_158),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_136),
.Y(n_129)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_144),
.Y(n_137)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_153),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_233),
.B(n_238),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_198),
.B(n_232),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_179),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_164),
.B(n_179),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_171),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_165),
.A2(n_171),
.B1(n_172),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_165),
.Y(n_230)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_192),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_180),
.B(n_193),
.C(n_197),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_188),
.B(n_189),
.Y(n_180)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_196),
.B2(n_197),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_224),
.B(n_231),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_212),
.B(n_223),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_211),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_208),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_222),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_222),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_229),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_229),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_235),
.Y(n_238)
);


endmodule