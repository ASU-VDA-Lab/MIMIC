module fake_jpeg_13992_n_346 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_346);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_346;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_12),
.Y(n_37)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_10),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_23),
.B(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_52),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_23),
.B(n_0),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_25),
.B(n_14),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_21),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx6_ASAP7_75t_SL g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx2_ASAP7_75t_R g70 ( 
.A(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_83),
.Y(n_113)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_71),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_63),
.A2(n_40),
.B1(n_37),
.B2(n_36),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_79),
.A2(n_27),
.B1(n_22),
.B2(n_49),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_81),
.B(n_82),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_25),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_40),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_62),
.A2(n_40),
.B1(n_37),
.B2(n_24),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_99),
.B1(n_104),
.B2(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_41),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_93),
.Y(n_128)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_41),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_35),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_97),
.B(n_98),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_35),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_44),
.A2(n_19),
.B1(n_26),
.B2(n_21),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_37),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_101),
.Y(n_146)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_45),
.A2(n_42),
.B1(n_29),
.B2(n_22),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_47),
.B(n_18),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_51),
.A2(n_24),
.B1(n_27),
.B2(n_39),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_110),
.A2(n_38),
.B1(n_34),
.B2(n_30),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_56),
.B(n_20),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_87),
.A2(n_24),
.B1(n_42),
.B2(n_29),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_116),
.A2(n_124),
.B1(n_151),
.B2(n_148),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_26),
.C(n_19),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_119),
.B(n_85),
.C(n_8),
.Y(n_172)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_100),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_122),
.B(n_137),
.Y(n_186)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_110),
.A2(n_34),
.B1(n_66),
.B2(n_18),
.Y(n_124)
);

AOI22x1_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_70),
.B1(n_111),
.B2(n_76),
.Y(n_153)
);

INVx3_ASAP7_75t_SL g127 ( 
.A(n_109),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g181 ( 
.A(n_127),
.Y(n_181)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_95),
.A2(n_34),
.B1(n_30),
.B2(n_3),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g161 ( 
.A1(n_129),
.A2(n_133),
.B1(n_111),
.B2(n_103),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_83),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_130)
);

OAI32xp33_ASAP7_75t_L g188 ( 
.A1(n_130),
.A2(n_14),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_188)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_131),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_132),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_91),
.A2(n_30),
.B1(n_2),
.B2(n_3),
.Y(n_133)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_138),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_84),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_84),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_105),
.A2(n_30),
.B1(n_4),
.B2(n_5),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_142),
.A2(n_71),
.B1(n_89),
.B2(n_80),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_102),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_147),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_102),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_76),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_153),
.A2(n_127),
.B1(n_129),
.B2(n_136),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_149),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_167),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_159),
.B(n_161),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_145),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_162),
.B(n_146),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_77),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_176),
.C(n_187),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_164),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_109),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_129),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_121),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_120),
.A2(n_102),
.B(n_69),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_170),
.A2(n_152),
.B(n_132),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_180),
.Y(n_190)
);

AND2x2_ASAP7_75t_SL g175 ( 
.A(n_120),
.B(n_69),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_150),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_113),
.B(n_88),
.C(n_86),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_124),
.A2(n_74),
.B1(n_68),
.B2(n_10),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_118),
.Y(n_178)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_131),
.Y(n_179)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_119),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_185),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_115),
.B(n_68),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_129),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_158),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_191),
.B(n_193),
.Y(n_238)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_194),
.B(n_205),
.Y(n_224)
);

NAND3xp33_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_204),
.C(n_175),
.Y(n_225)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_197),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_163),
.B(n_117),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_200),
.B(n_207),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_166),
.B(n_135),
.Y(n_204)
);

NOR2x1_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_130),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_157),
.A2(n_135),
.B(n_146),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_215),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_173),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_219),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_210),
.A2(n_132),
.B1(n_12),
.B2(n_13),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_138),
.C(n_125),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_171),
.C(n_160),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_165),
.Y(n_213)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_156),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_221),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_157),
.A2(n_125),
.B(n_150),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_217),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_170),
.A2(n_134),
.B(n_132),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_174),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_176),
.B(n_152),
.Y(n_219)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_208),
.A2(n_161),
.B1(n_159),
.B2(n_175),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_223),
.A2(n_227),
.B1(n_218),
.B2(n_211),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_L g262 ( 
.A1(n_225),
.A2(n_198),
.B(n_216),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_208),
.A2(n_161),
.B1(n_153),
.B2(n_181),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_155),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_228),
.B(n_237),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_233),
.A2(n_241),
.B(n_215),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_161),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_234),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_246),
.C(n_212),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_206),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_188),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_243),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_210),
.A2(n_153),
.B1(n_184),
.B2(n_171),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_240),
.A2(n_245),
.B1(n_201),
.B2(n_199),
.Y(n_254)
);

OA21x2_ASAP7_75t_L g241 ( 
.A1(n_208),
.A2(n_165),
.B(n_174),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_181),
.Y(n_243)
);

AND2x6_ASAP7_75t_L g244 ( 
.A(n_190),
.B(n_6),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_205),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_196),
.B(n_11),
.C(n_13),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_202),
.Y(n_247)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_202),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_248),
.Y(n_250)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_251),
.A2(n_229),
.B1(n_268),
.B2(n_234),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_252),
.A2(n_233),
.B(n_234),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_232),
.B(n_196),
.Y(n_253)
);

XNOR2x1_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_235),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_264),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_238),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_257),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_226),
.A2(n_199),
.B1(n_201),
.B2(n_217),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_258),
.A2(n_229),
.B(n_233),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_243),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_261),
.Y(n_284)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

NOR3xp33_ASAP7_75t_SL g287 ( 
.A(n_262),
.B(n_224),
.C(n_244),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_223),
.B(n_198),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_193),
.Y(n_289)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_246),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_203),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_226),
.Y(n_275)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_236),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_269),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_222),
.B(n_197),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_270),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_273),
.B(n_275),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_278),
.C(n_273),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_277),
.A2(n_285),
.B(n_258),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_226),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_271),
.B(n_231),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_288),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_282),
.A2(n_283),
.B1(n_286),
.B2(n_263),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_251),
.A2(n_240),
.B1(n_241),
.B2(n_229),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_241),
.B1(n_239),
.B2(n_227),
.Y(n_286)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_270),
.Y(n_288)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_303),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_291),
.A2(n_283),
.B1(n_286),
.B2(n_285),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_256),
.Y(n_292)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_292),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_284),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_293),
.B(n_297),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_294),
.Y(n_309)
);

AOI21xp33_ASAP7_75t_R g297 ( 
.A1(n_275),
.A2(n_256),
.B(n_267),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_289),
.Y(n_298)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_266),
.C(n_252),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_282),
.C(n_277),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_272),
.Y(n_302)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_302),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_257),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_272),
.B(n_269),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_304),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_290),
.C(n_301),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_310),
.A2(n_296),
.B1(n_291),
.B2(n_294),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_274),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_313),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_264),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_314),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_325),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_292),
.Y(n_319)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_319),
.Y(n_331)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_306),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_320),
.B(n_321),
.Y(n_326)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_307),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_322),
.B(n_324),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_310),
.A2(n_304),
.B1(n_254),
.B2(n_295),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_316),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_323),
.A2(n_315),
.B(n_308),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_327),
.A2(n_332),
.B(n_317),
.Y(n_333)
);

AOI21x1_ASAP7_75t_L g328 ( 
.A1(n_319),
.A2(n_309),
.B(n_287),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_328),
.B(n_265),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_318),
.A2(n_309),
.B(n_305),
.Y(n_332)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_333),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_330),
.B(n_324),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_334),
.B(n_336),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_331),
.A2(n_301),
.B(n_322),
.Y(n_335)
);

NAND3xp33_ASAP7_75t_SL g339 ( 
.A(n_335),
.B(n_337),
.C(n_326),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_221),
.Y(n_336)
);

OAI31xp33_ASAP7_75t_SL g342 ( 
.A1(n_339),
.A2(n_250),
.A3(n_259),
.B(n_261),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_338),
.A2(n_329),
.B1(n_280),
.B2(n_259),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_341),
.B(n_342),
.C(n_250),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_343),
.Y(n_344)
);

OAI321xp33_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_13),
.A3(n_192),
.B1(n_220),
.B2(n_340),
.C(n_338),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_192),
.Y(n_346)
);


endmodule