module fake_netlist_5_1535_n_191 (n_29, n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_30, n_20, n_5, n_14, n_2, n_31, n_23, n_13, n_3, n_6, n_191);

input n_29;
input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_14;
input n_2;
input n_31;
input n_23;
input n_13;
input n_3;
input n_6;

output n_191;

wire n_137;
wire n_168;
wire n_164;
wire n_91;
wire n_82;
wire n_122;
wire n_142;
wire n_176;
wire n_140;
wire n_124;
wire n_86;
wire n_136;
wire n_146;
wire n_182;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_180;
wire n_184;
wire n_78;
wire n_65;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_189;
wire n_165;
wire n_111;
wire n_108;
wire n_129;
wire n_66;
wire n_98;
wire n_177;
wire n_60;
wire n_155;
wire n_152;
wire n_43;
wire n_107;
wire n_69;
wire n_58;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_123;
wire n_139;
wire n_105;
wire n_80;
wire n_179;
wire n_125;
wire n_35;
wire n_167;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_156;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_157;
wire n_79;
wire n_131;
wire n_151;
wire n_47;
wire n_173;
wire n_53;
wire n_160;
wire n_188;
wire n_190;
wire n_158;
wire n_44;
wire n_40;
wire n_34;
wire n_154;
wire n_62;
wire n_138;
wire n_148;
wire n_71;
wire n_100;
wire n_109;
wire n_112;
wire n_85;
wire n_159;
wire n_163;
wire n_95;
wire n_119;
wire n_183;
wire n_185;
wire n_175;
wire n_169;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_181;
wire n_49;
wire n_39;
wire n_54;
wire n_147;
wire n_178;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_150;
wire n_170;
wire n_162;
wire n_77;
wire n_106;
wire n_102;
wire n_64;
wire n_161;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_174;
wire n_186;
wire n_134;
wire n_187;
wire n_32;
wire n_41;
wire n_104;
wire n_172;
wire n_103;
wire n_141;
wire n_51;
wire n_97;
wire n_63;
wire n_56;
wire n_166;
wire n_171;
wire n_153;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_20),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVxp67_ASAP7_75t_SL g34 ( 
.A(n_15),
.Y(n_34)
);

INVxp33_ASAP7_75t_SL g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

INVxp33_ASAP7_75t_SL g41 ( 
.A(n_24),
.Y(n_41)
);

INVxp67_ASAP7_75t_SL g42 ( 
.A(n_26),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

INVxp33_ASAP7_75t_SL g46 ( 
.A(n_9),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVxp33_ASAP7_75t_SL g53 ( 
.A(n_13),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_SL g58 ( 
.A(n_33),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_0),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_1),
.Y(n_61)
);

AND2x4_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_51),
.B(n_2),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_52),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_51),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_43),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

OAI221xp5_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_47),
.B1(n_49),
.B2(n_38),
.C(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

AO22x2_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_49),
.B1(n_42),
.B2(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

NAND2x1p5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_41),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_53),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_72),
.B(n_43),
.Y(n_86)
);

XNOR2x2_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_46),
.Y(n_87)
);

OAI221xp5_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_32),
.B1(n_40),
.B2(n_35),
.C(n_8),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_61),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_4),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_90),
.B1(n_79),
.B2(n_85),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_74),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_73),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_74),
.Y(n_98)
);

CKINVDCx11_ASAP7_75t_R g99 ( 
.A(n_87),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_73),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_74),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_79),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_86),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_103),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

BUFx4_ASAP7_75t_R g109 ( 
.A(n_99),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_98),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_98),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_97),
.B(n_92),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_79),
.B1(n_102),
.B2(n_97),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_102),
.Y(n_118)
);

NAND3xp33_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_105),
.C(n_108),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_107),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_118),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_112),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

OR2x6_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_112),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_120),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_65),
.B(n_117),
.Y(n_130)
);

NAND4xp25_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_88),
.C(n_64),
.D(n_70),
.Y(n_131)
);

NAND4xp25_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_64),
.C(n_70),
.D(n_69),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_123),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_133),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_126),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_124),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_117),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_134),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_130),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_141),
.A2(n_130),
.B1(n_132),
.B2(n_131),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_136),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

AOI221xp5_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_63),
.B1(n_58),
.B2(n_60),
.C(n_69),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_137),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_146),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_140),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_139),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_60),
.Y(n_155)
);

OAI211xp5_ASAP7_75t_L g156 ( 
.A1(n_145),
.A2(n_148),
.B(n_143),
.C(n_142),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_127),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_68),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_68),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_73),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_149),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_160),
.Y(n_163)
);

NOR3xp33_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_153),
.C(n_159),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_56),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_56),
.Y(n_169)
);

OAI221xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_81),
.B1(n_89),
.B2(n_100),
.C(n_84),
.Y(n_170)
);

NOR3x1_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_89),
.C(n_109),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

OA21x2_ASAP7_75t_L g173 ( 
.A1(n_163),
.A2(n_100),
.B(n_101),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_169),
.A2(n_81),
.B(n_73),
.Y(n_174)
);

INVxp67_ASAP7_75t_SL g175 ( 
.A(n_165),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_6),
.Y(n_176)
);

OA211x2_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_109),
.B(n_8),
.C(n_10),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_170),
.A2(n_162),
.B1(n_167),
.B2(n_164),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_174),
.A2(n_58),
.B1(n_81),
.B2(n_114),
.Y(n_179)
);

AOI31xp33_ASAP7_75t_SL g180 ( 
.A1(n_171),
.A2(n_7),
.A3(n_11),
.B(n_12),
.Y(n_180)
);

NAND4xp75_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_7),
.C(n_12),
.D(n_101),
.Y(n_181)
);

AND2x4_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_113),
.Y(n_182)
);

AND4x1_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_176),
.C(n_172),
.D(n_175),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_178),
.A2(n_173),
.B1(n_176),
.B2(n_114),
.Y(n_184)
);

AOI322xp5_ASAP7_75t_L g185 ( 
.A1(n_180),
.A2(n_181),
.A3(n_182),
.B1(n_173),
.B2(n_58),
.C1(n_113),
.C2(n_115),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_173),
.Y(n_186)
);

OAI322xp33_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_114),
.A3(n_113),
.B1(n_115),
.B2(n_22),
.C1(n_25),
.C2(n_29),
.Y(n_187)
);

OAI322xp33_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_114),
.A3(n_18),
.B1(n_21),
.B2(n_30),
.C1(n_14),
.C2(n_94),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_183),
.A2(n_114),
.B1(n_96),
.B2(n_94),
.Y(n_189)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_185),
.B(n_96),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_188),
.B1(n_187),
.B2(n_94),
.Y(n_191)
);


endmodule