module fake_jpeg_18565_n_187 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_187);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_31),
.B(n_32),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_SL g32 ( 
.A(n_17),
.B(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_14),
.B(n_2),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_43),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_17),
.Y(n_35)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_37),
.B(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_25),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_25),
.Y(n_44)
);

CKINVDCx12_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_27),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_29),
.B1(n_14),
.B2(n_16),
.Y(n_48)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_33),
.Y(n_68)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_35),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_26),
.B1(n_23),
.B2(n_29),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_55),
.B1(n_62),
.B2(n_37),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_23),
.B1(n_26),
.B2(n_16),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_32),
.A2(n_45),
.B1(n_44),
.B2(n_43),
.Y(n_62)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_65),
.Y(n_93)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_67),
.Y(n_97)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_71),
.Y(n_103)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_70),
.A2(n_77),
.B1(n_78),
.B2(n_2),
.Y(n_111)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_39),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_74),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_23),
.B1(n_36),
.B2(n_31),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_73),
.A2(n_76),
.B1(n_79),
.B2(n_24),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_56),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_36),
.B1(n_31),
.B2(n_16),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_36),
.B1(n_35),
.B2(n_40),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_47),
.A2(n_40),
.B1(n_41),
.B2(n_30),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_15),
.B1(n_19),
.B2(n_30),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_81),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_46),
.B(n_19),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_15),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_49),
.A2(n_28),
.B1(n_27),
.B2(n_20),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_86),
.A2(n_92),
.B1(n_52),
.B2(n_57),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_58),
.Y(n_88)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_21),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_66),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_40),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_94),
.A2(n_99),
.B1(n_75),
.B2(n_8),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_52),
.B(n_34),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_96),
.A2(n_75),
.B(n_6),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_21),
.C(n_28),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_107),
.C(n_75),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_41),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_106),
.B(n_111),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_21),
.C(n_20),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_69),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_71),
.B(n_80),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_115),
.A2(n_99),
.B(n_93),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_116),
.B(n_118),
.Y(n_142)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_95),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_90),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_121),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_92),
.C(n_87),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_82),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_123),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_87),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_110),
.B(n_9),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_124),
.B(n_11),
.Y(n_136)
);

AO21x1_ASAP7_75t_L g133 ( 
.A1(n_125),
.A2(n_126),
.B(n_108),
.Y(n_133)
);

AO21x1_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_5),
.B(n_7),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_127),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_100),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

OAI32xp33_ASAP7_75t_L g132 ( 
.A1(n_120),
.A2(n_96),
.A3(n_111),
.B1(n_106),
.B2(n_112),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_132),
.B(n_140),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_144),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_134),
.A2(n_143),
.B(n_129),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_136),
.B(n_11),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_114),
.A2(n_107),
.B1(n_109),
.B2(n_98),
.Y(n_139)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_100),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_108),
.B(n_113),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_122),
.C(n_116),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_147),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_146),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_121),
.C(n_119),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_143),
.A2(n_125),
.B1(n_126),
.B2(n_115),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_149),
.A2(n_134),
.B1(n_135),
.B2(n_8),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_137),
.Y(n_151)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_104),
.Y(n_152)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_152),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_156),
.Y(n_164)
);

INVxp33_ASAP7_75t_SL g155 ( 
.A(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

AOI322xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_8),
.A3(n_12),
.B1(n_104),
.B2(n_129),
.C1(n_132),
.C2(n_142),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_154),
.A2(n_139),
.B1(n_138),
.B2(n_140),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_165),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_147),
.C(n_145),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_171),
.C(n_163),
.Y(n_174)
);

NAND2xp67_ASAP7_75t_SL g167 ( 
.A(n_160),
.B(n_149),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_168),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_158),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_154),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_165),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_176),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_170),
.A2(n_164),
.B1(n_148),
.B2(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_175),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_164),
.C(n_158),
.Y(n_177)
);

OAI21x1_ASAP7_75t_L g180 ( 
.A1(n_177),
.A2(n_167),
.B(n_153),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_180),
.A2(n_173),
.B(n_170),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_169),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_181),
.B(n_173),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_179),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_184),
.C(n_161),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_157),
.B1(n_135),
.B2(n_162),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_12),
.Y(n_187)
);


endmodule