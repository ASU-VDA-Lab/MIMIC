module fake_jpeg_6651_n_46 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

BUFx5_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx6_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx10_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_17),
.A2(n_7),
.B1(n_13),
.B2(n_3),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_18),
.B(n_21),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_1),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_20),
.B(n_9),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_26),
.B1(n_19),
.B2(n_17),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_22),
.B1(n_27),
.B2(n_20),
.Y(n_33)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_30),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_16),
.B(n_15),
.C(n_14),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

AOI221xp5_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_32),
.B1(n_10),
.B2(n_14),
.C(n_6),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_15),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_35),
.A2(n_29),
.B(n_15),
.Y(n_38)
);

XNOR2x1_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_39),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_36),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_43),
.B(n_23),
.Y(n_44)
);

AOI322xp5_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_34),
.A3(n_23),
.B1(n_14),
.B2(n_10),
.C1(n_6),
.C2(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);


endmodule