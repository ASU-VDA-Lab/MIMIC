module fake_aes_8503_n_26 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_26);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_26;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
NOR2xp33_ASAP7_75t_R g13 ( .A(n_1), .B(n_4), .Y(n_13) );
INVxp67_ASAP7_75t_L g14 ( .A(n_11), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_8), .Y(n_15) );
AOI22xp5_ASAP7_75t_L g16 ( .A1(n_0), .A2(n_10), .B1(n_3), .B2(n_5), .Y(n_16) );
NOR2xp33_ASAP7_75t_R g17 ( .A(n_9), .B(n_7), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_14), .Y(n_18) );
AOI21xp5_ASAP7_75t_L g19 ( .A1(n_15), .A2(n_6), .B(n_12), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_18), .B(n_16), .Y(n_20) );
INVx4_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
OAI22xp33_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_20), .B1(n_15), .B2(n_19), .Y(n_22) );
OAI211xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_13), .B(n_17), .C(n_2), .Y(n_23) );
CKINVDCx12_ASAP7_75t_R g24 ( .A(n_23), .Y(n_24) );
XNOR2xp5_ASAP7_75t_L g25 ( .A(n_24), .B(n_0), .Y(n_25) );
AOI22xp33_ASAP7_75t_SL g26 ( .A1(n_25), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_26) );
endmodule