module fake_ibex_69_n_855 (n_151, n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_855);

input n_151;
input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_855;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_418;
wire n_256;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_593;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_187;
wire n_667;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_723;
wire n_270;
wire n_170;
wire n_383;
wire n_346;
wire n_840;
wire n_561;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_791;
wire n_715;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_439;
wire n_433;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_564;
wire n_562;
wire n_506;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_397;
wire n_366;
wire n_803;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_415;
wire n_597;
wire n_288;
wire n_320;
wire n_247;
wire n_285;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_342;
wire n_385;
wire n_414;
wire n_233;
wire n_430;
wire n_807;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_668;
wire n_779;
wire n_266;
wire n_294;
wire n_485;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_693;
wire n_311;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_687;
wire n_202;
wire n_298;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_559;
wire n_425;

INVx2_ASAP7_75t_L g165 ( 
.A(n_118),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_10),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_97),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_164),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_57),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_22),
.Y(n_172)
);

INVxp33_ASAP7_75t_L g173 ( 
.A(n_107),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_56),
.B(n_44),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_76),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_31),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_114),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_146),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_52),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_26),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_21),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_36),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_109),
.Y(n_185)
);

INVxp67_ASAP7_75t_SL g186 ( 
.A(n_100),
.Y(n_186)
);

BUFx2_ASAP7_75t_SL g187 ( 
.A(n_158),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_48),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_92),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_66),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_122),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_135),
.Y(n_192)
);

BUFx10_ASAP7_75t_L g193 ( 
.A(n_11),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_22),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_88),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_106),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_46),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_116),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_115),
.Y(n_199)
);

NOR2xp67_ASAP7_75t_L g200 ( 
.A(n_133),
.B(n_6),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_55),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_23),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_87),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_136),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_111),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_127),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_18),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_159),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_42),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_61),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_123),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_18),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_150),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_125),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_38),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_74),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_120),
.Y(n_218)
);

INVxp33_ASAP7_75t_SL g219 ( 
.A(n_80),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_5),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_30),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_91),
.Y(n_222)
);

INVxp67_ASAP7_75t_SL g223 ( 
.A(n_34),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_144),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_1),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_145),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_17),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_16),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_81),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_37),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_143),
.Y(n_231)
);

CKINVDCx11_ASAP7_75t_R g232 ( 
.A(n_43),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_142),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_16),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_79),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_151),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_60),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_82),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_45),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_99),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_128),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_89),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_53),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_62),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_117),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_28),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_24),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_132),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_83),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_84),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_73),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_34),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_29),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_37),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_59),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_39),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_71),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_41),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_35),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_148),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_157),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_10),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_131),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_160),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_119),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_54),
.Y(n_266)
);

INVxp33_ASAP7_75t_SL g267 ( 
.A(n_65),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_140),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_141),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_101),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_205),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_221),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_232),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_219),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_274)
);

OAI21x1_ASAP7_75t_L g275 ( 
.A1(n_165),
.A2(n_85),
.B(n_162),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_202),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_207),
.B(n_246),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_218),
.B(n_3),
.Y(n_278)
);

AND2x4_ASAP7_75t_L g279 ( 
.A(n_202),
.B(n_4),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_221),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_221),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_172),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_240),
.B(n_6),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_232),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_175),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_175),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_229),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_221),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_176),
.Y(n_289)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_239),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_249),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_172),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_194),
.B(n_7),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_234),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_254),
.Y(n_295)
);

CKINVDCx6p67_ASAP7_75t_R g296 ( 
.A(n_239),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_219),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_173),
.B(n_8),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_254),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_197),
.Y(n_300)
);

AND2x2_ASAP7_75t_SL g301 ( 
.A(n_167),
.B(n_168),
.Y(n_301)
);

BUFx12f_ASAP7_75t_L g302 ( 
.A(n_193),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_262),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_197),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_234),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_261),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_267),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_307)
);

AND2x4_ASAP7_75t_L g308 ( 
.A(n_259),
.B(n_12),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_173),
.B(n_13),
.Y(n_309)
);

BUFx12f_ASAP7_75t_L g310 ( 
.A(n_193),
.Y(n_310)
);

INVx6_ASAP7_75t_L g311 ( 
.A(n_193),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_261),
.Y(n_312)
);

AND2x4_ASAP7_75t_L g313 ( 
.A(n_166),
.B(n_14),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_178),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_180),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_262),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_182),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_234),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_177),
.B(n_15),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_184),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_171),
.B(n_195),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_181),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_234),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_213),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_227),
.B(n_19),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_228),
.B(n_20),
.Y(n_326)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_247),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_247),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_188),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_189),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_252),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_253),
.B(n_223),
.Y(n_332)
);

AND2x4_ASAP7_75t_L g333 ( 
.A(n_191),
.B(n_20),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_198),
.Y(n_334)
);

OAI21x1_ASAP7_75t_L g335 ( 
.A1(n_201),
.A2(n_95),
.B(n_161),
.Y(n_335)
);

OAI21x1_ASAP7_75t_L g336 ( 
.A1(n_204),
.A2(n_94),
.B(n_154),
.Y(n_336)
);

BUFx12f_ASAP7_75t_L g337 ( 
.A(n_247),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_270),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_206),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_214),
.B(n_21),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_209),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_267),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_272),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_272),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_279),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_R g346 ( 
.A(n_273),
.B(n_266),
.Y(n_346)
);

INVx5_ASAP7_75t_L g347 ( 
.A(n_279),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_272),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_272),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_279),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_280),
.Y(n_351)
);

NAND2xp33_ASAP7_75t_L g352 ( 
.A(n_340),
.B(n_179),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_301),
.A2(n_269),
.B1(n_169),
.B2(n_192),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_322),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_280),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_327),
.B(n_215),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_327),
.B(n_251),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_321),
.B(n_251),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_328),
.B(n_287),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_280),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_311),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_329),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_329),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_329),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_R g365 ( 
.A(n_284),
.B(n_322),
.Y(n_365)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_311),
.Y(n_366)
);

AO21x2_ASAP7_75t_L g367 ( 
.A1(n_275),
.A2(n_212),
.B(n_211),
.Y(n_367)
);

INVx11_ASAP7_75t_L g368 ( 
.A(n_302),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_308),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_311),
.B(n_255),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_328),
.B(n_291),
.Y(n_371)
);

NAND2xp33_ASAP7_75t_SL g372 ( 
.A(n_340),
.B(n_169),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_301),
.B(n_257),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_276),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_284),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_280),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_281),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_308),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_275),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_339),
.B(n_257),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_281),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_281),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_313),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_288),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_302),
.B(n_258),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_310),
.B(n_258),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_277),
.B(n_303),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_310),
.B(n_260),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_L g389 ( 
.A1(n_313),
.A2(n_220),
.B1(n_225),
.B2(n_230),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_337),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_337),
.B(n_333),
.Y(n_391)
);

NAND2xp33_ASAP7_75t_L g392 ( 
.A(n_338),
.B(n_260),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_290),
.B(n_263),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_313),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_325),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_333),
.B(n_263),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_325),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_338),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_338),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_290),
.B(n_264),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_296),
.Y(n_401)
);

AND3x2_ASAP7_75t_L g402 ( 
.A(n_325),
.B(n_186),
.C(n_256),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_296),
.Y(n_403)
);

NOR2x1p5_ASAP7_75t_L g404 ( 
.A(n_332),
.B(n_183),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_326),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_326),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_333),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_331),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_298),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_314),
.B(n_265),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_331),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_294),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_294),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_332),
.B(n_265),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_335),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_320),
.B(n_187),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_309),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_SL g418 ( 
.A1(n_316),
.A2(n_269),
.B1(n_185),
.B2(n_192),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_278),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_285),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_L g421 ( 
.A1(n_324),
.A2(n_243),
.B1(n_250),
.B2(n_231),
.Y(n_421)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_315),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_285),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_294),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_286),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_283),
.A2(n_185),
.B1(n_222),
.B2(n_224),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_305),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_341),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_305),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_317),
.B(n_190),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_409),
.B(n_317),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_419),
.B(n_293),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_401),
.B(n_319),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_408),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_417),
.B(n_196),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_370),
.B(n_330),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_358),
.B(n_330),
.Y(n_437)
);

INVx2_ASAP7_75t_SL g438 ( 
.A(n_370),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_380),
.B(n_334),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_416),
.B(n_334),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_368),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_398),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_416),
.B(n_199),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_411),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_414),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_410),
.B(n_282),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_391),
.B(n_271),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_387),
.B(n_282),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_387),
.B(n_292),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_403),
.B(n_342),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_359),
.B(n_295),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_404),
.A2(n_274),
.B1(n_297),
.B2(n_307),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_354),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_393),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_379),
.Y(n_455)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_368),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_390),
.B(n_292),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_378),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_373),
.A2(n_352),
.B1(n_389),
.B2(n_426),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_402),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_398),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_374),
.B(n_292),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_407),
.A2(n_394),
.B1(n_395),
.B2(n_383),
.Y(n_463)
);

NAND2xp33_ASAP7_75t_L g464 ( 
.A(n_415),
.B(n_203),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_371),
.B(n_299),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_397),
.B(n_208),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_379),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_396),
.A2(n_335),
.B(n_336),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_403),
.B(n_210),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_405),
.A2(n_174),
.B1(n_304),
.B2(n_289),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_406),
.B(n_216),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_372),
.B(n_289),
.Y(n_472)
);

NAND3xp33_ASAP7_75t_L g473 ( 
.A(n_352),
.B(n_341),
.C(n_244),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_428),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_345),
.A2(n_336),
.B(n_300),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_385),
.B(n_300),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_430),
.B(n_235),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_365),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_422),
.Y(n_479)
);

NOR2x1p5_ASAP7_75t_L g480 ( 
.A(n_375),
.B(n_236),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_350),
.B(n_238),
.Y(n_481)
);

NAND2xp33_ASAP7_75t_L g482 ( 
.A(n_415),
.B(n_248),
.Y(n_482)
);

OR2x2_ASAP7_75t_SL g483 ( 
.A(n_418),
.B(n_217),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_372),
.B(n_304),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_369),
.A2(n_306),
.B1(n_312),
.B2(n_341),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_400),
.B(n_306),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_347),
.B(n_361),
.Y(n_487)
);

O2A1O1Ixp33_ASAP7_75t_L g488 ( 
.A1(n_386),
.A2(n_237),
.B(n_226),
.C(n_233),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_347),
.B(n_170),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_420),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_361),
.B(n_241),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_366),
.B(n_268),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_366),
.B(n_341),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_423),
.A2(n_341),
.B1(n_245),
.B2(n_242),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_425),
.Y(n_495)
);

OAI22xp33_ASAP7_75t_L g496 ( 
.A1(n_353),
.A2(n_200),
.B1(n_323),
.B2(n_305),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_421),
.B(n_323),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_356),
.B(n_323),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_357),
.B(n_318),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_388),
.B(n_318),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_392),
.B(n_25),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_392),
.B(n_26),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_379),
.B(n_40),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_367),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_367),
.B(n_27),
.Y(n_505)
);

AOI21x1_ASAP7_75t_L g506 ( 
.A1(n_475),
.A2(n_468),
.B(n_504),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_431),
.B(n_346),
.Y(n_507)
);

AND2x2_ASAP7_75t_SL g508 ( 
.A(n_456),
.B(n_415),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_456),
.B(n_367),
.Y(n_509)
);

CKINVDCx10_ASAP7_75t_R g510 ( 
.A(n_441),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_453),
.B(n_362),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_447),
.A2(n_362),
.B1(n_363),
.B2(n_364),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_445),
.B(n_363),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_457),
.Y(n_514)
);

NOR2xp67_ASAP7_75t_L g515 ( 
.A(n_460),
.B(n_27),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_469),
.B(n_364),
.Y(n_516)
);

INVxp67_ASAP7_75t_SL g517 ( 
.A(n_470),
.Y(n_517)
);

BUFx8_ASAP7_75t_SL g518 ( 
.A(n_447),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_454),
.A2(n_486),
.B(n_439),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_455),
.Y(n_520)
);

INVx3_ASAP7_75t_SL g521 ( 
.A(n_476),
.Y(n_521)
);

AND2x6_ASAP7_75t_L g522 ( 
.A(n_458),
.B(n_399),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_448),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_440),
.B(n_30),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_449),
.B(n_31),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_432),
.Y(n_526)
);

NOR2xp67_ASAP7_75t_L g527 ( 
.A(n_452),
.B(n_32),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_437),
.B(n_438),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_459),
.A2(n_429),
.B1(n_427),
.B2(n_424),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_478),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_437),
.A2(n_413),
.B(n_412),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_463),
.A2(n_436),
.B(n_455),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_503),
.A2(n_413),
.B(n_412),
.Y(n_533)
);

O2A1O1Ixp33_ASAP7_75t_L g534 ( 
.A1(n_496),
.A2(n_384),
.B(n_382),
.C(n_381),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_478),
.B(n_480),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_479),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_490),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_450),
.A2(n_351),
.B1(n_377),
.B2(n_376),
.Y(n_538)
);

AO21x1_ASAP7_75t_L g539 ( 
.A1(n_505),
.A2(n_502),
.B(n_501),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_483),
.A2(n_360),
.B1(n_355),
.B2(n_351),
.Y(n_540)
);

AO21x1_ASAP7_75t_L g541 ( 
.A1(n_491),
.A2(n_493),
.B(n_499),
.Y(n_541)
);

AO21x1_ASAP7_75t_L g542 ( 
.A1(n_491),
.A2(n_355),
.B(n_349),
.Y(n_542)
);

O2A1O1Ixp33_ASAP7_75t_L g543 ( 
.A1(n_472),
.A2(n_348),
.B(n_344),
.C(n_343),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_495),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_462),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_435),
.B(n_33),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_434),
.A2(n_105),
.B(n_152),
.Y(n_547)
);

O2A1O1Ixp33_ASAP7_75t_L g548 ( 
.A1(n_484),
.A2(n_33),
.B(n_35),
.C(n_36),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_476),
.B(n_163),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_467),
.A2(n_47),
.B(n_49),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_443),
.A2(n_50),
.B(n_51),
.Y(n_551)
);

NAND3xp33_ASAP7_75t_L g552 ( 
.A(n_473),
.B(n_58),
.C(n_63),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_465),
.B(n_451),
.Y(n_553)
);

A2O1A1Ixp33_ASAP7_75t_L g554 ( 
.A1(n_444),
.A2(n_64),
.B(n_67),
.C(n_68),
.Y(n_554)
);

O2A1O1Ixp33_ASAP7_75t_L g555 ( 
.A1(n_446),
.A2(n_69),
.B(n_70),
.C(n_72),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_497),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_485),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_465),
.B(n_433),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_489),
.Y(n_559)
);

O2A1O1Ixp33_ASAP7_75t_L g560 ( 
.A1(n_488),
.A2(n_147),
.B(n_90),
.C(n_93),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_500),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_466),
.A2(n_86),
.B1(n_96),
.B2(n_98),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_485),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_563)
);

OR2x6_ASAP7_75t_L g564 ( 
.A(n_471),
.B(n_108),
.Y(n_564)
);

O2A1O1Ixp33_ASAP7_75t_L g565 ( 
.A1(n_481),
.A2(n_110),
.B(n_112),
.C(n_113),
.Y(n_565)
);

BUFx12f_ASAP7_75t_L g566 ( 
.A(n_494),
.Y(n_566)
);

O2A1O1Ixp33_ASAP7_75t_L g567 ( 
.A1(n_477),
.A2(n_121),
.B(n_124),
.C(n_126),
.Y(n_567)
);

NOR3xp33_ASAP7_75t_L g568 ( 
.A(n_492),
.B(n_130),
.C(n_134),
.Y(n_568)
);

AO21x2_ASAP7_75t_L g569 ( 
.A1(n_464),
.A2(n_137),
.B(n_138),
.Y(n_569)
);

CKINVDCx10_ASAP7_75t_R g570 ( 
.A(n_498),
.Y(n_570)
);

CKINVDCx8_ASAP7_75t_R g571 ( 
.A(n_498),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_487),
.B(n_139),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_523),
.B(n_442),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_517),
.B(n_482),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_537),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_528),
.B(n_461),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_566),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_SL g578 ( 
.A(n_516),
.B(n_474),
.Y(n_578)
);

OAI21x1_ASAP7_75t_SL g579 ( 
.A1(n_547),
.A2(n_541),
.B(n_563),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_544),
.Y(n_580)
);

AO32x2_ASAP7_75t_L g581 ( 
.A1(n_540),
.A2(n_529),
.A3(n_557),
.B1(n_563),
.B2(n_542),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_521),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_553),
.B(n_558),
.Y(n_583)
);

NAND2xp33_ASAP7_75t_R g584 ( 
.A(n_509),
.B(n_564),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_518),
.Y(n_585)
);

BUFx2_ASAP7_75t_L g586 ( 
.A(n_559),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_525),
.B(n_526),
.Y(n_587)
);

AOI21xp33_ASAP7_75t_L g588 ( 
.A1(n_509),
.A2(n_535),
.B(n_508),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_530),
.B(n_545),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_524),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_514),
.B(n_546),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_510),
.Y(n_592)
);

BUFx12f_ASAP7_75t_L g593 ( 
.A(n_564),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_570),
.Y(n_594)
);

AO31x2_ASAP7_75t_L g595 ( 
.A1(n_529),
.A2(n_554),
.A3(n_557),
.B(n_556),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_571),
.B(n_512),
.Y(n_596)
);

A2O1A1Ixp33_ASAP7_75t_L g597 ( 
.A1(n_560),
.A2(n_534),
.B(n_543),
.C(n_551),
.Y(n_597)
);

INVx5_ASAP7_75t_L g598 ( 
.A(n_522),
.Y(n_598)
);

AO31x2_ASAP7_75t_L g599 ( 
.A1(n_550),
.A2(n_549),
.A3(n_531),
.B(n_572),
.Y(n_599)
);

CKINVDCx8_ASAP7_75t_R g600 ( 
.A(n_522),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_513),
.B(n_511),
.Y(n_601)
);

AO21x1_ASAP7_75t_L g602 ( 
.A1(n_567),
.A2(n_555),
.B(n_568),
.Y(n_602)
);

CKINVDCx11_ASAP7_75t_R g603 ( 
.A(n_515),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_565),
.A2(n_569),
.B(n_552),
.Y(n_604)
);

AO31x2_ASAP7_75t_L g605 ( 
.A1(n_522),
.A2(n_539),
.A3(n_541),
.B(n_542),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_522),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_538),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_562),
.B(n_387),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_514),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_518),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_536),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_537),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_537),
.Y(n_613)
);

AOI221x1_ASAP7_75t_L g614 ( 
.A1(n_540),
.A2(n_532),
.B1(n_505),
.B2(n_568),
.C(n_547),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_519),
.A2(n_533),
.B(n_532),
.Y(n_615)
);

NOR3xp33_ASAP7_75t_L g616 ( 
.A(n_507),
.B(n_527),
.C(n_517),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_566),
.Y(n_617)
);

AOI21x1_ASAP7_75t_L g618 ( 
.A1(n_506),
.A2(n_539),
.B(n_541),
.Y(n_618)
);

NOR2xp67_ASAP7_75t_L g619 ( 
.A(n_527),
.B(n_456),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_518),
.B(n_453),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_517),
.B(n_431),
.Y(n_621)
);

AO31x2_ASAP7_75t_L g622 ( 
.A1(n_539),
.A2(n_541),
.A3(n_542),
.B(n_504),
.Y(n_622)
);

NOR4xp25_ASAP7_75t_L g623 ( 
.A(n_548),
.B(n_496),
.C(n_540),
.D(n_342),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_519),
.A2(n_533),
.B(n_532),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_519),
.A2(n_533),
.B(n_532),
.Y(n_625)
);

A2O1A1Ixp33_ASAP7_75t_L g626 ( 
.A1(n_519),
.A2(n_437),
.B(n_532),
.C(n_561),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_520),
.Y(n_627)
);

AOI21x1_ASAP7_75t_L g628 ( 
.A1(n_506),
.A2(n_539),
.B(n_541),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_537),
.Y(n_629)
);

AO22x2_ASAP7_75t_L g630 ( 
.A1(n_540),
.A2(n_470),
.B1(n_517),
.B2(n_453),
.Y(n_630)
);

AO32x2_ASAP7_75t_L g631 ( 
.A1(n_540),
.A2(n_529),
.A3(n_563),
.B1(n_557),
.B2(n_539),
.Y(n_631)
);

BUFx2_ASAP7_75t_SL g632 ( 
.A(n_527),
.Y(n_632)
);

OR2x6_ASAP7_75t_L g633 ( 
.A(n_527),
.B(n_456),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_517),
.B(n_431),
.Y(n_634)
);

A2O1A1Ixp33_ASAP7_75t_L g635 ( 
.A1(n_519),
.A2(n_437),
.B(n_532),
.C(n_561),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_523),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_523),
.Y(n_637)
);

BUFx10_ASAP7_75t_L g638 ( 
.A(n_546),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_523),
.B(n_387),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_523),
.Y(n_640)
);

NOR3xp33_ASAP7_75t_L g641 ( 
.A(n_507),
.B(n_527),
.C(n_517),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_517),
.B(n_431),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_517),
.B(n_431),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_517),
.B(n_431),
.Y(n_644)
);

AOI21xp33_ASAP7_75t_SL g645 ( 
.A1(n_592),
.A2(n_594),
.B(n_620),
.Y(n_645)
);

AO31x2_ASAP7_75t_L g646 ( 
.A1(n_614),
.A2(n_624),
.A3(n_615),
.B(n_625),
.Y(n_646)
);

CKINVDCx11_ASAP7_75t_R g647 ( 
.A(n_610),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_SL g648 ( 
.A(n_600),
.B(n_593),
.Y(n_648)
);

AOI21xp33_ASAP7_75t_SL g649 ( 
.A1(n_633),
.A2(n_584),
.B(n_616),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_583),
.B(n_639),
.Y(n_650)
);

BUFx10_ASAP7_75t_L g651 ( 
.A(n_633),
.Y(n_651)
);

AO21x2_ASAP7_75t_L g652 ( 
.A1(n_579),
.A2(n_604),
.B(n_628),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_609),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_580),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_585),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_612),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_586),
.B(n_617),
.Y(n_657)
);

AO31x2_ASAP7_75t_L g658 ( 
.A1(n_626),
.A2(n_635),
.A3(n_602),
.B(n_597),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_640),
.B(n_589),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_577),
.B(n_636),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_596),
.B(n_577),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_613),
.Y(n_662)
);

BUFx2_ASAP7_75t_R g663 ( 
.A(n_632),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_621),
.B(n_644),
.Y(n_664)
);

CKINVDCx11_ASAP7_75t_R g665 ( 
.A(n_582),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_629),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_603),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_606),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_634),
.B(n_643),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_642),
.B(n_608),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_578),
.A2(n_590),
.B(n_574),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_641),
.A2(n_630),
.B1(n_619),
.B2(n_607),
.Y(n_672)
);

OA21x2_ASAP7_75t_L g673 ( 
.A1(n_588),
.A2(n_581),
.B(n_622),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_598),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_598),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g676 ( 
.A1(n_623),
.A2(n_587),
.B(n_576),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_598),
.B(n_611),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_637),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_591),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_573),
.B(n_601),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_573),
.Y(n_681)
);

OA21x2_ASAP7_75t_L g682 ( 
.A1(n_581),
.A2(n_622),
.B(n_631),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_630),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_627),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_638),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_638),
.B(n_601),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_622),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_605),
.B(n_595),
.Y(n_688)
);

AO31x2_ASAP7_75t_L g689 ( 
.A1(n_631),
.A2(n_605),
.A3(n_595),
.B(n_599),
.Y(n_689)
);

OA21x2_ASAP7_75t_L g690 ( 
.A1(n_605),
.A2(n_595),
.B(n_599),
.Y(n_690)
);

AO31x2_ASAP7_75t_L g691 ( 
.A1(n_599),
.A2(n_539),
.A3(n_614),
.B(n_615),
.Y(n_691)
);

OA21x2_ASAP7_75t_L g692 ( 
.A1(n_614),
.A2(n_604),
.B(n_618),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_575),
.Y(n_693)
);

NAND2x1p5_ASAP7_75t_L g694 ( 
.A(n_598),
.B(n_606),
.Y(n_694)
);

BUFx2_ASAP7_75t_L g695 ( 
.A(n_586),
.Y(n_695)
);

INVx4_ASAP7_75t_L g696 ( 
.A(n_598),
.Y(n_696)
);

NAND2x1p5_ASAP7_75t_L g697 ( 
.A(n_598),
.B(n_606),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_575),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_575),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_575),
.Y(n_700)
);

AOI211xp5_ASAP7_75t_L g701 ( 
.A1(n_616),
.A2(n_527),
.B(n_641),
.C(n_496),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_575),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_586),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_575),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_650),
.B(n_664),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_650),
.B(n_664),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_687),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_654),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_656),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_662),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_666),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_659),
.B(n_679),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_693),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_646),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_698),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_676),
.B(n_670),
.Y(n_716)
);

BUFx2_ASAP7_75t_L g717 ( 
.A(n_684),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_699),
.B(n_704),
.Y(n_718)
);

BUFx2_ASAP7_75t_SL g719 ( 
.A(n_668),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_700),
.B(n_702),
.Y(n_720)
);

INVxp67_ASAP7_75t_L g721 ( 
.A(n_695),
.Y(n_721)
);

OAI21xp5_ASAP7_75t_SL g722 ( 
.A1(n_649),
.A2(n_672),
.B(n_645),
.Y(n_722)
);

OAI21xp5_ASAP7_75t_L g723 ( 
.A1(n_671),
.A2(n_669),
.B(n_701),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_673),
.B(n_680),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_651),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_683),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_647),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_691),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_703),
.Y(n_729)
);

AO21x1_ASAP7_75t_L g730 ( 
.A1(n_688),
.A2(n_696),
.B(n_677),
.Y(n_730)
);

OR2x6_ASAP7_75t_L g731 ( 
.A(n_694),
.B(n_697),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_658),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_661),
.B(n_657),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_673),
.B(n_689),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_673),
.B(n_680),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_661),
.B(n_681),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_694),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_658),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_680),
.B(n_653),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_724),
.B(n_690),
.Y(n_740)
);

NOR2x1_ASAP7_75t_L g741 ( 
.A(n_722),
.B(n_696),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_716),
.B(n_682),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_719),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_724),
.B(n_735),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_707),
.Y(n_745)
);

AOI222xp33_ASAP7_75t_L g746 ( 
.A1(n_705),
.A2(n_648),
.B1(n_651),
.B2(n_647),
.C1(n_665),
.C2(n_686),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_706),
.B(n_665),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_719),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_735),
.B(n_690),
.Y(n_749)
);

NOR2x1p5_ASAP7_75t_L g750 ( 
.A(n_737),
.B(n_674),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_712),
.B(n_685),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_718),
.B(n_720),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_716),
.B(n_690),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_733),
.A2(n_677),
.B1(n_678),
.B2(n_682),
.Y(n_754)
);

OR2x6_ASAP7_75t_L g755 ( 
.A(n_730),
.B(n_697),
.Y(n_755)
);

AND2x4_ASAP7_75t_SL g756 ( 
.A(n_731),
.B(n_677),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_726),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_720),
.B(n_689),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_732),
.B(n_658),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_736),
.A2(n_668),
.B1(n_674),
.B2(n_675),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_723),
.A2(n_653),
.B1(n_660),
.B2(n_675),
.Y(n_761)
);

BUFx2_ASAP7_75t_L g762 ( 
.A(n_730),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_717),
.B(n_652),
.Y(n_763)
);

INVx4_ASAP7_75t_L g764 ( 
.A(n_731),
.Y(n_764)
);

NAND2xp33_ASAP7_75t_R g765 ( 
.A(n_731),
.B(n_663),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_717),
.B(n_692),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_737),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_745),
.Y(n_768)
);

INVxp67_ASAP7_75t_SL g769 ( 
.A(n_766),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_744),
.B(n_738),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_745),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_767),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_744),
.B(n_738),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_747),
.B(n_727),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_752),
.B(n_711),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_740),
.B(n_714),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_753),
.B(n_734),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_758),
.B(n_753),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_758),
.B(n_742),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_740),
.B(n_728),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_749),
.B(n_728),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_778),
.B(n_749),
.Y(n_782)
);

INVxp67_ASAP7_75t_L g783 ( 
.A(n_772),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_775),
.B(n_757),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_778),
.B(n_759),
.Y(n_785)
);

INVxp67_ASAP7_75t_L g786 ( 
.A(n_769),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_776),
.B(n_762),
.Y(n_787)
);

OR2x2_ASAP7_75t_L g788 ( 
.A(n_777),
.B(n_742),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_770),
.B(n_773),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_768),
.Y(n_790)
);

OR2x2_ASAP7_75t_L g791 ( 
.A(n_777),
.B(n_763),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_780),
.B(n_781),
.Y(n_792)
);

AND2x4_ASAP7_75t_L g793 ( 
.A(n_776),
.B(n_762),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_771),
.Y(n_794)
);

INVxp33_ASAP7_75t_L g795 ( 
.A(n_791),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_782),
.B(n_780),
.Y(n_796)
);

OAI211xp5_ASAP7_75t_L g797 ( 
.A1(n_786),
.A2(n_746),
.B(n_748),
.C(n_743),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_782),
.B(n_789),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_789),
.B(n_781),
.Y(n_799)
);

AND2x2_ASAP7_75t_SL g800 ( 
.A(n_787),
.B(n_764),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_794),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_794),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_785),
.B(n_776),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_790),
.Y(n_804)
);

OR2x2_ASAP7_75t_L g805 ( 
.A(n_792),
.B(n_779),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_791),
.B(n_779),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_800),
.A2(n_764),
.B1(n_788),
.B2(n_783),
.Y(n_807)
);

NAND2x1_ASAP7_75t_L g808 ( 
.A(n_798),
.B(n_787),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_798),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_804),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_799),
.B(n_796),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_803),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_806),
.B(n_788),
.Y(n_813)
);

AOI221xp5_ASAP7_75t_L g814 ( 
.A1(n_795),
.A2(n_784),
.B1(n_721),
.B2(n_785),
.C(n_751),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_797),
.A2(n_793),
.B1(n_787),
.B2(n_746),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_804),
.Y(n_816)
);

A2O1A1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_808),
.A2(n_800),
.B(n_796),
.C(n_799),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_812),
.B(n_803),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_811),
.B(n_806),
.Y(n_819)
);

OAI22xp33_ASAP7_75t_SL g820 ( 
.A1(n_815),
.A2(n_805),
.B1(n_764),
.B2(n_760),
.Y(n_820)
);

AOI21xp33_ASAP7_75t_L g821 ( 
.A1(n_820),
.A2(n_774),
.B(n_765),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_817),
.A2(n_807),
.B(n_814),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_818),
.B(n_807),
.Y(n_823)
);

NAND3xp33_ASAP7_75t_L g824 ( 
.A(n_822),
.B(n_729),
.C(n_816),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_823),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_825),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_824),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_826),
.A2(n_821),
.B(n_667),
.C(n_655),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_827),
.B(n_819),
.Y(n_829)
);

XNOR2xp5_ASAP7_75t_L g830 ( 
.A(n_829),
.B(n_667),
.Y(n_830)
);

NAND3xp33_ASAP7_75t_SL g831 ( 
.A(n_828),
.B(n_826),
.C(n_655),
.Y(n_831)
);

OAI21x1_ASAP7_75t_SL g832 ( 
.A1(n_830),
.A2(n_725),
.B(n_741),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_831),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_830),
.B(n_810),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_833),
.A2(n_725),
.B(n_741),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_834),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_832),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_833),
.A2(n_809),
.B1(n_760),
.B2(n_761),
.Y(n_838)
);

AOI22x1_ASAP7_75t_L g839 ( 
.A1(n_833),
.A2(n_750),
.B1(n_813),
.B2(n_764),
.Y(n_839)
);

AOI221xp5_ASAP7_75t_L g840 ( 
.A1(n_837),
.A2(n_711),
.B1(n_710),
.B2(n_708),
.C(n_709),
.Y(n_840)
);

AOI21x1_ASAP7_75t_L g841 ( 
.A1(n_836),
.A2(n_739),
.B(n_731),
.Y(n_841)
);

AOI21xp33_ASAP7_75t_SL g842 ( 
.A1(n_839),
.A2(n_805),
.B(n_767),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_838),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_835),
.A2(n_713),
.B(n_708),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_836),
.B(n_801),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_838),
.A2(n_750),
.B1(n_754),
.B2(n_755),
.Y(n_846)
);

XNOR2xp5_ASAP7_75t_L g847 ( 
.A(n_843),
.B(n_709),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_844),
.B(n_710),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_846),
.A2(n_801),
.B1(n_793),
.B2(n_737),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_845),
.A2(n_793),
.B1(n_802),
.B2(n_713),
.Y(n_850)
);

OA21x2_ASAP7_75t_L g851 ( 
.A1(n_847),
.A2(n_841),
.B(n_848),
.Y(n_851)
);

OA21x2_ASAP7_75t_L g852 ( 
.A1(n_849),
.A2(n_840),
.B(n_842),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_852),
.B(n_850),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_851),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_854),
.A2(n_853),
.B1(n_756),
.B2(n_715),
.Y(n_855)
);


endmodule