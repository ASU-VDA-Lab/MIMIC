module real_aes_7376_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_119;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_148;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g550 ( .A1(n_0), .A2(n_175), .B(n_551), .C(n_554), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_1), .B(n_501), .Y(n_555) );
INVx1_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
INVx1_ASAP7_75t_L g187 ( .A(n_3), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_4), .B(n_147), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_5), .A2(n_474), .B(n_495), .Y(n_494) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_6), .A2(n_167), .B(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_7), .A2(n_38), .B1(n_141), .B2(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_8), .B(n_167), .Y(n_176) );
AND2x6_ASAP7_75t_L g159 ( .A(n_9), .B(n_160), .Y(n_159) );
A2O1A1Ixp33_ASAP7_75t_L g563 ( .A1(n_10), .A2(n_159), .B(n_479), .C(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g110 ( .A(n_11), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_11), .B(n_39), .Y(n_435) );
INVx1_ASAP7_75t_L g137 ( .A(n_12), .Y(n_137) );
INVx1_ASAP7_75t_L g180 ( .A(n_13), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_14), .B(n_145), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_15), .B(n_147), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_16), .B(n_133), .Y(n_251) );
AO32x2_ASAP7_75t_L g193 ( .A1(n_17), .A2(n_132), .A3(n_158), .B1(n_167), .B2(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_18), .B(n_141), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_19), .B(n_133), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_20), .A2(n_54), .B1(n_141), .B2(n_196), .Y(n_197) );
AOI22xp33_ASAP7_75t_SL g235 ( .A1(n_21), .A2(n_81), .B1(n_141), .B2(n_145), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_22), .B(n_141), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_23), .A2(n_158), .B(n_479), .C(n_528), .Y(n_527) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_24), .A2(n_60), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_24), .Y(n_123) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_25), .A2(n_158), .B(n_479), .C(n_507), .Y(n_506) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_26), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_27), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_28), .B(n_440), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_29), .A2(n_474), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_30), .B(n_162), .Y(n_210) );
INVx2_ASAP7_75t_L g143 ( .A(n_31), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_32), .A2(n_477), .B(n_487), .C(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_33), .B(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_34), .B(n_162), .Y(n_221) );
XNOR2x2_ASAP7_75t_SL g120 ( .A(n_35), .B(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_36), .B(n_217), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_37), .A2(n_85), .B1(n_456), .B2(n_457), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_37), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_39), .B(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_40), .B(n_526), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_41), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_42), .B(n_147), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_43), .B(n_474), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_44), .A2(n_477), .B(n_481), .C(n_487), .Y(n_476) );
OAI321xp33_ASAP7_75t_L g119 ( .A1(n_45), .A2(n_120), .A3(n_429), .B1(n_436), .B2(n_437), .C(n_439), .Y(n_119) );
INVx1_ASAP7_75t_L g436 ( .A(n_45), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_46), .B(n_141), .Y(n_170) );
INVx1_ASAP7_75t_L g552 ( .A(n_47), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_48), .A2(n_91), .B1(n_196), .B2(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g482 ( .A(n_49), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_50), .B(n_141), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_51), .B(n_141), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_52), .B(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_53), .B(n_153), .Y(n_174) );
AOI22xp33_ASAP7_75t_SL g249 ( .A1(n_55), .A2(n_61), .B1(n_141), .B2(n_145), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_56), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_57), .B(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_58), .B(n_141), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_59), .B(n_141), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_60), .Y(n_124) );
OAI22xp5_ASAP7_75t_SL g462 ( .A1(n_60), .A2(n_124), .B1(n_125), .B2(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g160 ( .A(n_62), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_63), .B(n_474), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_64), .B(n_501), .Y(n_500) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_65), .A2(n_153), .B(n_183), .C(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_66), .B(n_141), .Y(n_188) );
INVx1_ASAP7_75t_L g136 ( .A(n_67), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_68), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_69), .B(n_147), .Y(n_519) );
AO32x2_ASAP7_75t_L g231 ( .A1(n_70), .A2(n_158), .A3(n_167), .B1(n_232), .B2(n_236), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_71), .B(n_148), .Y(n_565) );
INVx1_ASAP7_75t_L g151 ( .A(n_72), .Y(n_151) );
INVx1_ASAP7_75t_L g205 ( .A(n_73), .Y(n_205) );
CKINVDCx16_ASAP7_75t_R g549 ( .A(n_74), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_75), .B(n_484), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_76), .A2(n_479), .B(n_487), .C(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_77), .B(n_145), .Y(n_206) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_78), .Y(n_496) );
INVx1_ASAP7_75t_L g115 ( .A(n_79), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_80), .B(n_483), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_82), .B(n_196), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_83), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_84), .B(n_145), .Y(n_209) );
INVx1_ASAP7_75t_L g457 ( .A(n_85), .Y(n_457) );
INVx2_ASAP7_75t_L g134 ( .A(n_86), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_87), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_88), .B(n_157), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_89), .B(n_145), .Y(n_171) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_90), .B(n_112), .C(n_113), .Y(n_111) );
OR2x2_ASAP7_75t_L g432 ( .A(n_90), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g449 ( .A(n_90), .Y(n_449) );
OR2x2_ASAP7_75t_L g461 ( .A(n_90), .B(n_434), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_92), .A2(n_103), .B1(n_145), .B2(n_146), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_93), .B(n_474), .Y(n_515) );
INVx1_ASAP7_75t_L g518 ( .A(n_94), .Y(n_518) );
INVxp67_ASAP7_75t_L g499 ( .A(n_95), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_96), .B(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_97), .B(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g540 ( .A(n_98), .Y(n_540) );
INVx1_ASAP7_75t_L g561 ( .A(n_99), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_100), .A2(n_105), .B1(n_116), .B2(n_770), .Y(n_104) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_101), .A2(n_453), .B1(n_454), .B2(n_455), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_101), .Y(n_453) );
AND2x2_ASAP7_75t_L g489 ( .A(n_102), .B(n_162), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx5_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
CKINVDCx9p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
BUFx2_ASAP7_75t_L g770 ( .A(n_108), .Y(n_770) );
OR2x4_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
AND2x2_ASAP7_75t_L g434 ( .A(n_112), .B(n_435), .Y(n_434) );
OA211x2_ASAP7_75t_L g116 ( .A1(n_113), .A2(n_117), .B(n_119), .C(n_443), .Y(n_116) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g444 ( .A(n_118), .Y(n_444) );
NAND2x1p5_ASAP7_75t_L g437 ( .A(n_120), .B(n_438), .Y(n_437) );
XNOR2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_125), .Y(n_121) );
INVx1_ASAP7_75t_SL g463 ( .A(n_125), .Y(n_463) );
OR3x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_357), .C(n_406), .Y(n_125) );
NAND5xp2_ASAP7_75t_L g126 ( .A(n_127), .B(n_272), .C(n_300), .D(n_330), .E(n_344), .Y(n_126) );
AOI221xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_190), .B1(n_222), .B2(n_227), .C(n_238), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_129), .B(n_163), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_129), .B(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g252 ( .A(n_130), .Y(n_252) );
AND2x2_ASAP7_75t_L g260 ( .A(n_130), .B(n_166), .Y(n_260) );
AND2x2_ASAP7_75t_L g283 ( .A(n_130), .B(n_165), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_130), .B(n_177), .Y(n_298) );
OR2x2_ASAP7_75t_L g307 ( .A(n_130), .B(n_245), .Y(n_307) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_130), .Y(n_310) );
AND2x2_ASAP7_75t_L g418 ( .A(n_130), .B(n_245), .Y(n_418) );
OA21x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_138), .B(n_161), .Y(n_130) );
OA21x2_ASAP7_75t_L g177 ( .A1(n_131), .A2(n_178), .B(n_189), .Y(n_177) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_132), .B(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_133), .Y(n_167) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x2_ASAP7_75t_SL g162 ( .A(n_134), .B(n_135), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
OAI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_150), .B(n_158), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_144), .B(n_147), .Y(n_139) );
INVx3_ASAP7_75t_L g204 ( .A(n_141), .Y(n_204) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_141), .Y(n_542) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g196 ( .A(n_142), .Y(n_196) );
BUFx3_ASAP7_75t_L g234 ( .A(n_142), .Y(n_234) );
AND2x6_ASAP7_75t_L g479 ( .A(n_142), .B(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g146 ( .A(n_143), .Y(n_146) );
INVx1_ASAP7_75t_L g154 ( .A(n_143), .Y(n_154) );
INVx2_ASAP7_75t_L g181 ( .A(n_145), .Y(n_181) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_147), .A2(n_170), .B(n_171), .Y(n_169) );
INVx2_ASAP7_75t_L g175 ( .A(n_147), .Y(n_175) );
O2A1O1Ixp5_ASAP7_75t_SL g203 ( .A1(n_147), .A2(n_204), .B(n_205), .C(n_206), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_147), .B(n_499), .Y(n_498) );
INVx5_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
OAI22xp5_ASAP7_75t_SL g232 ( .A1(n_148), .A2(n_157), .B1(n_233), .B2(n_235), .Y(n_232) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_149), .Y(n_157) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_149), .Y(n_185) );
INVx1_ASAP7_75t_L g217 ( .A(n_149), .Y(n_217) );
AND2x2_ASAP7_75t_L g475 ( .A(n_149), .B(n_154), .Y(n_475) );
INVx1_ASAP7_75t_L g480 ( .A(n_149), .Y(n_480) );
O2A1O1Ixp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_155), .C(n_156), .Y(n_150) );
O2A1O1Ixp33_ASAP7_75t_L g186 ( .A1(n_152), .A2(n_175), .B(n_187), .C(n_188), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_152), .A2(n_529), .B(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_156), .A2(n_219), .B(n_220), .Y(n_218) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
OAI22xp5_ASAP7_75t_L g194 ( .A1(n_157), .A2(n_175), .B1(n_195), .B2(n_197), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_157), .A2(n_175), .B1(n_248), .B2(n_249), .Y(n_247) );
INVx4_ASAP7_75t_L g553 ( .A(n_157), .Y(n_553) );
NAND3xp33_ASAP7_75t_L g271 ( .A(n_158), .B(n_246), .C(n_247), .Y(n_271) );
BUFx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
OAI21xp5_ASAP7_75t_L g168 ( .A1(n_159), .A2(n_169), .B(n_172), .Y(n_168) );
OAI21xp5_ASAP7_75t_L g178 ( .A1(n_159), .A2(n_179), .B(n_186), .Y(n_178) );
OAI21xp5_ASAP7_75t_L g202 ( .A1(n_159), .A2(n_203), .B(n_207), .Y(n_202) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_159), .A2(n_213), .B(n_218), .Y(n_212) );
AND2x4_ASAP7_75t_L g474 ( .A(n_159), .B(n_475), .Y(n_474) );
INVx4_ASAP7_75t_SL g488 ( .A(n_159), .Y(n_488) );
NAND2x1p5_ASAP7_75t_L g562 ( .A(n_159), .B(n_475), .Y(n_562) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_162), .A2(n_202), .B(n_210), .Y(n_201) );
OA21x2_ASAP7_75t_L g211 ( .A1(n_162), .A2(n_212), .B(n_221), .Y(n_211) );
INVx2_ASAP7_75t_L g236 ( .A(n_162), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_162), .A2(n_473), .B(n_476), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_162), .A2(n_515), .B(n_516), .Y(n_514) );
INVx1_ASAP7_75t_L g534 ( .A(n_162), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_163), .B(n_310), .Y(n_366) );
INVx2_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
OAI311xp33_ASAP7_75t_L g308 ( .A1(n_164), .A2(n_309), .A3(n_310), .B1(n_311), .C1(n_326), .Y(n_308) );
AND2x2_ASAP7_75t_L g164 ( .A(n_165), .B(n_177), .Y(n_164) );
AND2x2_ASAP7_75t_L g269 ( .A(n_165), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g276 ( .A(n_165), .Y(n_276) );
AND2x2_ASAP7_75t_L g397 ( .A(n_165), .B(n_226), .Y(n_397) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_166), .B(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g253 ( .A(n_166), .B(n_177), .Y(n_253) );
AND2x2_ASAP7_75t_L g305 ( .A(n_166), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g319 ( .A(n_166), .B(n_252), .Y(n_319) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_176), .Y(n_166) );
INVx4_ASAP7_75t_L g246 ( .A(n_167), .Y(n_246) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_167), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_167), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_175), .Y(n_172) );
INVx2_ASAP7_75t_L g226 ( .A(n_177), .Y(n_226) );
AND2x2_ASAP7_75t_L g268 ( .A(n_177), .B(n_252), .Y(n_268) );
O2A1O1Ixp33_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_182), .C(n_183), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_181), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_181), .A2(n_565), .B(n_566), .Y(n_564) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_183), .A2(n_540), .B(n_541), .C(n_542), .Y(n_539) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_184), .A2(n_208), .B(n_209), .Y(n_207) );
INVx4_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g484 ( .A(n_185), .Y(n_484) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_198), .Y(n_190) );
OR2x2_ASAP7_75t_L g363 ( .A(n_191), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_191), .B(n_369), .Y(n_380) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_192), .B(n_376), .Y(n_375) );
BUFx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g237 ( .A(n_193), .Y(n_237) );
AND2x2_ASAP7_75t_L g304 ( .A(n_193), .B(n_231), .Y(n_304) );
AND2x2_ASAP7_75t_L g315 ( .A(n_193), .B(n_211), .Y(n_315) );
AND2x2_ASAP7_75t_L g324 ( .A(n_193), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_198), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_198), .B(n_265), .Y(n_309) );
INVx2_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
OR2x2_ASAP7_75t_L g296 ( .A(n_199), .B(n_255), .Y(n_296) );
OR2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_211), .Y(n_199) );
INVx2_ASAP7_75t_L g229 ( .A(n_200), .Y(n_229) );
AND2x2_ASAP7_75t_L g323 ( .A(n_200), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g241 ( .A(n_201), .Y(n_241) );
OR2x2_ASAP7_75t_L g340 ( .A(n_201), .B(n_341), .Y(n_340) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_201), .Y(n_403) );
AND2x2_ASAP7_75t_L g242 ( .A(n_211), .B(n_237), .Y(n_242) );
INVx1_ASAP7_75t_L g263 ( .A(n_211), .Y(n_263) );
AND2x2_ASAP7_75t_L g284 ( .A(n_211), .B(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g325 ( .A(n_211), .Y(n_325) );
INVx1_ASAP7_75t_L g341 ( .A(n_211), .Y(n_341) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_211), .Y(n_416) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_216), .Y(n_213) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVxp67_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_224), .B(n_329), .Y(n_370) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_224), .A2(n_314), .B1(n_363), .B2(n_373), .Y(n_372) );
INVx1_ASAP7_75t_SL g224 ( .A(n_225), .Y(n_224) );
OAI211xp5_ASAP7_75t_SL g406 ( .A1(n_225), .A2(n_407), .B(n_409), .C(n_427), .Y(n_406) );
INVx2_ASAP7_75t_L g259 ( .A(n_226), .Y(n_259) );
AND2x2_ASAP7_75t_L g317 ( .A(n_226), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g328 ( .A(n_226), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_227), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_230), .Y(n_227) );
AND2x2_ASAP7_75t_L g301 ( .A(n_228), .B(n_265), .Y(n_301) );
BUFx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g333 ( .A(n_229), .B(n_324), .Y(n_333) );
AND2x2_ASAP7_75t_L g352 ( .A(n_229), .B(n_266), .Y(n_352) );
AND2x4_ASAP7_75t_L g288 ( .A(n_230), .B(n_262), .Y(n_288) );
AND2x2_ASAP7_75t_L g426 ( .A(n_230), .B(n_402), .Y(n_426) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_237), .Y(n_230) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_231), .Y(n_255) );
INVx1_ASAP7_75t_L g266 ( .A(n_231), .Y(n_266) );
INVx1_ASAP7_75t_L g365 ( .A(n_231), .Y(n_365) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_234), .Y(n_486) );
INVx2_ASAP7_75t_L g554 ( .A(n_234), .Y(n_554) );
INVx1_ASAP7_75t_L g531 ( .A(n_236), .Y(n_531) );
OR2x2_ASAP7_75t_L g256 ( .A(n_237), .B(n_241), .Y(n_256) );
AND2x2_ASAP7_75t_L g265 ( .A(n_237), .B(n_266), .Y(n_265) );
NOR2xp67_ASAP7_75t_L g285 ( .A(n_237), .B(n_286), .Y(n_285) );
OAI221xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_243), .B1(n_254), .B2(n_257), .C(n_261), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_240), .A2(n_262), .B(n_264), .C(n_267), .Y(n_261) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
INVx1_ASAP7_75t_L g286 ( .A(n_241), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_241), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_SL g369 ( .A(n_241), .B(n_263), .Y(n_369) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_241), .Y(n_376) );
AND2x2_ASAP7_75t_L g294 ( .A(n_242), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g331 ( .A(n_242), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_253), .Y(n_243) );
INVx2_ASAP7_75t_L g322 ( .A(n_244), .Y(n_322) );
AOI222xp33_ASAP7_75t_L g371 ( .A1(n_244), .A2(n_255), .B1(n_372), .B2(n_374), .C1(n_375), .C2(n_377), .Y(n_371) );
AND2x2_ASAP7_75t_L g428 ( .A(n_244), .B(n_397), .Y(n_428) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_252), .Y(n_244) );
INVx1_ASAP7_75t_L g318 ( .A(n_245), .Y(n_318) );
AO21x1_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_247), .B(n_250), .Y(n_245) );
INVx3_ASAP7_75t_L g501 ( .A(n_246), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_246), .B(n_521), .Y(n_520) );
AO21x2_ASAP7_75t_L g536 ( .A1(n_246), .A2(n_537), .B(n_544), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_246), .B(n_545), .Y(n_544) );
AO21x2_ASAP7_75t_L g559 ( .A1(n_246), .A2(n_560), .B(n_567), .Y(n_559) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x4_ASAP7_75t_L g270 ( .A(n_251), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g356 ( .A(n_253), .B(n_290), .Y(n_356) );
AOI21xp33_ASAP7_75t_L g367 ( .A1(n_254), .A2(n_368), .B(n_370), .Y(n_367) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx2_ASAP7_75t_L g295 ( .A(n_255), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_255), .B(n_262), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_255), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
INVx3_ASAP7_75t_L g321 ( .A(n_259), .Y(n_321) );
OR2x2_ASAP7_75t_L g373 ( .A(n_259), .B(n_295), .Y(n_373) );
AND2x2_ASAP7_75t_L g289 ( .A(n_260), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g327 ( .A(n_260), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_260), .B(n_321), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_260), .B(n_317), .Y(n_343) );
AND2x2_ASAP7_75t_L g347 ( .A(n_260), .B(n_329), .Y(n_347) );
INVxp67_ASAP7_75t_L g279 ( .A(n_262), .Y(n_279) );
BUFx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OAI22xp5_ASAP7_75t_L g336 ( .A1(n_264), .A2(n_337), .B1(n_342), .B2(n_343), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_264), .B(n_369), .Y(n_399) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g385 ( .A(n_265), .B(n_376), .Y(n_385) );
AND2x2_ASAP7_75t_L g414 ( .A(n_265), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g419 ( .A(n_265), .B(n_369), .Y(n_419) );
INVx1_ASAP7_75t_L g332 ( .A(n_266), .Y(n_332) );
BUFx2_ASAP7_75t_L g338 ( .A(n_266), .Y(n_338) );
INVx1_ASAP7_75t_L g423 ( .A(n_267), .Y(n_423) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
NAND2x1p5_ASAP7_75t_L g274 ( .A(n_268), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g299 ( .A(n_269), .Y(n_299) );
NOR2x1_ASAP7_75t_L g275 ( .A(n_270), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g282 ( .A(n_270), .B(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g291 ( .A(n_270), .Y(n_291) );
INVx3_ASAP7_75t_L g329 ( .A(n_270), .Y(n_329) );
OR2x2_ASAP7_75t_L g395 ( .A(n_270), .B(n_396), .Y(n_395) );
AOI211xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_277), .B(n_280), .C(n_292), .Y(n_272) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_273), .A2(n_410), .B1(n_417), .B2(n_419), .C(n_420), .Y(n_409) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_281), .B(n_287), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_283), .B(n_321), .Y(n_335) );
AND2x2_ASAP7_75t_L g377 ( .A(n_283), .B(n_317), .Y(n_377) );
INVx1_ASAP7_75t_SL g390 ( .A(n_284), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_284), .B(n_338), .Y(n_393) );
INVx1_ASAP7_75t_L g411 ( .A(n_285), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g378 ( .A1(n_289), .A2(n_379), .B1(n_381), .B2(n_385), .C(n_386), .Y(n_378) );
AND2x2_ASAP7_75t_L g405 ( .A(n_290), .B(n_397), .Y(n_405) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g389 ( .A(n_291), .Y(n_389) );
AOI21xp33_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_296), .B(n_297), .Y(n_292) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g360 ( .A(n_295), .B(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g346 ( .A(n_296), .Y(n_346) );
INVx1_ASAP7_75t_L g374 ( .A(n_297), .Y(n_374) );
OR2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
O2A1O1Ixp33_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_302), .B(n_305), .C(n_308), .Y(n_300) );
OAI31xp33_ASAP7_75t_L g427 ( .A1(n_301), .A2(n_339), .A3(n_426), .B(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g401 ( .A(n_304), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g422 ( .A(n_304), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_306), .B(n_321), .Y(n_349) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g424 ( .A(n_307), .B(n_321), .Y(n_424) );
AOI22xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_316), .B1(n_320), .B2(n_323), .Y(n_311) );
NAND2xp33_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_315), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g351 ( .A(n_315), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g354 ( .A(n_315), .B(n_338), .Y(n_354) );
AND2x2_ASAP7_75t_L g408 ( .A(n_315), .B(n_403), .Y(n_408) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
INVx1_ASAP7_75t_L g383 ( .A(n_319), .Y(n_383) );
NOR2xp67_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
OAI32xp33_ASAP7_75t_L g386 ( .A1(n_321), .A2(n_355), .A3(n_387), .B1(n_389), .B2(n_390), .Y(n_386) );
INVx1_ASAP7_75t_L g361 ( .A(n_324), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_324), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g384 ( .A(n_328), .Y(n_384) );
O2A1O1Ixp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_333), .B(n_334), .C(n_336), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_332), .B(n_369), .Y(n_368) );
AOI221xp5_ASAP7_75t_L g344 ( .A1(n_333), .A2(n_345), .B1(n_346), .B2(n_347), .C(n_348), .Y(n_344) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g345 ( .A(n_343), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_350), .B1(n_353), .B2(n_355), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NAND4xp25_ASAP7_75t_SL g410 ( .A(n_353), .B(n_411), .C(n_412), .D(n_413), .Y(n_410) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
NAND4xp25_ASAP7_75t_SL g357 ( .A(n_358), .B(n_371), .C(n_378), .D(n_391), .Y(n_357) );
O2A1O1Ixp33_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_362), .B(n_366), .C(n_367), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_SL g388 ( .A(n_364), .Y(n_388) );
INVx2_ASAP7_75t_L g412 ( .A(n_369), .Y(n_412) );
OR2x2_ASAP7_75t_L g421 ( .A(n_376), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_394), .B(n_398), .Y(n_391) );
INVxp67_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g417 ( .A(n_397), .B(n_418), .Y(n_417) );
AOI21xp33_ASAP7_75t_SL g398 ( .A1(n_399), .A2(n_400), .B(n_404), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
CKINVDCx16_ASAP7_75t_R g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_423), .B1(n_424), .B2(n_425), .Y(n_420) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g438 ( .A(n_431), .Y(n_438) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_SL g442 ( .A(n_432), .Y(n_442) );
NOR2x2_ASAP7_75t_L g448 ( .A(n_433), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g466 ( .A(n_434), .B(n_449), .Y(n_466) );
NAND4xp25_ASAP7_75t_SL g443 ( .A(n_439), .B(n_444), .C(n_445), .D(n_450), .Y(n_443) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx3_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B1(n_458), .B2(n_765), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_462), .B1(n_464), .B2(n_467), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g766 ( .A(n_460), .Y(n_766) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g767 ( .A(n_462), .Y(n_767) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g768 ( .A(n_465), .Y(n_768) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx4_ASAP7_75t_L g769 ( .A(n_467), .Y(n_769) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
OR5x1_ASAP7_75t_L g468 ( .A(n_469), .B(n_638), .C(n_716), .D(n_740), .E(n_757), .Y(n_468) );
OAI211xp5_ASAP7_75t_SL g469 ( .A1(n_470), .A2(n_510), .B(n_556), .C(n_615), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_490), .Y(n_470) );
AND2x2_ASAP7_75t_L g569 ( .A(n_471), .B(n_492), .Y(n_569) );
INVx5_ASAP7_75t_SL g597 ( .A(n_471), .Y(n_597) );
AND2x2_ASAP7_75t_L g633 ( .A(n_471), .B(n_618), .Y(n_633) );
OR2x2_ASAP7_75t_L g672 ( .A(n_471), .B(n_491), .Y(n_672) );
OR2x2_ASAP7_75t_L g703 ( .A(n_471), .B(n_594), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_471), .B(n_607), .Y(n_739) );
AND2x2_ASAP7_75t_L g751 ( .A(n_471), .B(n_594), .Y(n_751) );
OR2x6_ASAP7_75t_L g471 ( .A(n_472), .B(n_489), .Y(n_471) );
BUFx2_ASAP7_75t_L g526 ( .A(n_474), .Y(n_526) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_478), .A2(n_488), .B(n_496), .C(n_497), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_SL g548 ( .A1(n_478), .A2(n_488), .B(n_549), .C(n_550), .Y(n_548) );
INVx5_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B(n_485), .C(n_486), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g517 ( .A1(n_483), .A2(n_486), .B(n_518), .C(n_519), .Y(n_517) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g750 ( .A(n_490), .B(n_751), .Y(n_750) );
INVx1_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
OR2x2_ASAP7_75t_L g613 ( .A(n_491), .B(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_502), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_492), .B(n_594), .Y(n_593) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_492), .Y(n_606) );
INVx3_ASAP7_75t_L g621 ( .A(n_492), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_492), .B(n_502), .Y(n_645) );
OR2x2_ASAP7_75t_L g654 ( .A(n_492), .B(n_597), .Y(n_654) );
AND2x2_ASAP7_75t_L g658 ( .A(n_492), .B(n_618), .Y(n_658) );
AND2x2_ASAP7_75t_L g664 ( .A(n_492), .B(n_665), .Y(n_664) );
INVxp67_ASAP7_75t_L g701 ( .A(n_492), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_492), .B(n_559), .Y(n_715) );
OA21x2_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_494), .B(n_500), .Y(n_492) );
OA21x2_ASAP7_75t_L g546 ( .A1(n_501), .A2(n_547), .B(n_555), .Y(n_546) );
OR2x2_ASAP7_75t_L g607 ( .A(n_502), .B(n_559), .Y(n_607) );
AND2x2_ASAP7_75t_L g618 ( .A(n_502), .B(n_594), .Y(n_618) );
AND2x2_ASAP7_75t_L g630 ( .A(n_502), .B(n_621), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_502), .B(n_559), .Y(n_653) );
INVx1_ASAP7_75t_SL g665 ( .A(n_502), .Y(n_665) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g558 ( .A(n_503), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_503), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_522), .Y(n_511) );
AND2x2_ASAP7_75t_L g578 ( .A(n_512), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_512), .B(n_535), .Y(n_582) );
AND2x2_ASAP7_75t_L g585 ( .A(n_512), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_512), .B(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g610 ( .A(n_512), .B(n_601), .Y(n_610) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_512), .Y(n_629) );
AND2x2_ASAP7_75t_L g650 ( .A(n_512), .B(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g660 ( .A(n_512), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g706 ( .A(n_512), .B(n_589), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_512), .B(n_612), .Y(n_733) );
INVx5_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
BUFx2_ASAP7_75t_L g603 ( .A(n_513), .Y(n_603) );
AND2x2_ASAP7_75t_L g669 ( .A(n_513), .B(n_601), .Y(n_669) );
AND2x2_ASAP7_75t_L g753 ( .A(n_513), .B(n_621), .Y(n_753) );
OR2x6_ASAP7_75t_L g513 ( .A(n_514), .B(n_520), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_522), .B(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g742 ( .A(n_522), .Y(n_742) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_535), .Y(n_522) );
AND2x2_ASAP7_75t_L g572 ( .A(n_523), .B(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g581 ( .A(n_523), .B(n_579), .Y(n_581) );
INVx5_ASAP7_75t_L g589 ( .A(n_523), .Y(n_589) );
AND2x2_ASAP7_75t_L g612 ( .A(n_523), .B(n_546), .Y(n_612) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_523), .Y(n_649) );
OR2x6_ASAP7_75t_L g523 ( .A(n_524), .B(n_532), .Y(n_523) );
AOI21xp5_ASAP7_75t_SL g524 ( .A1(n_525), .A2(n_527), .B(n_531), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
INVx1_ASAP7_75t_L g690 ( .A(n_535), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_535), .B(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g723 ( .A(n_535), .B(n_589), .Y(n_723) );
A2O1A1Ixp33_ASAP7_75t_L g752 ( .A1(n_535), .A2(n_646), .B(n_753), .C(n_754), .Y(n_752) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_546), .Y(n_535) );
BUFx2_ASAP7_75t_L g573 ( .A(n_536), .Y(n_573) );
INVx2_ASAP7_75t_L g577 ( .A(n_536), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_543), .Y(n_537) );
INVx2_ASAP7_75t_L g579 ( .A(n_546), .Y(n_579) );
AND2x2_ASAP7_75t_L g586 ( .A(n_546), .B(n_577), .Y(n_586) );
AND2x2_ASAP7_75t_L g677 ( .A(n_546), .B(n_589), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
AOI211x1_ASAP7_75t_SL g556 ( .A1(n_557), .A2(n_570), .B(n_583), .C(n_608), .Y(n_556) );
INVx1_ASAP7_75t_L g674 ( .A(n_557), .Y(n_674) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_569), .Y(n_557) );
INVx5_ASAP7_75t_SL g594 ( .A(n_559), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_559), .B(n_664), .Y(n_663) );
AOI311xp33_ASAP7_75t_L g682 ( .A1(n_559), .A2(n_683), .A3(n_685), .B(n_686), .C(n_692), .Y(n_682) );
A2O1A1Ixp33_ASAP7_75t_L g717 ( .A1(n_559), .A2(n_630), .B(n_718), .C(n_721), .Y(n_717) );
OAI21xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_562), .B(n_563), .Y(n_560) );
INVxp67_ASAP7_75t_L g637 ( .A(n_569), .Y(n_637) );
NAND4xp25_ASAP7_75t_SL g570 ( .A(n_571), .B(n_574), .C(n_580), .D(n_582), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_571), .B(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g628 ( .A(n_572), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_578), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_575), .B(n_581), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_575), .B(n_588), .Y(n_708) );
BUFx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_576), .B(n_589), .Y(n_726) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g601 ( .A(n_577), .Y(n_601) );
INVxp67_ASAP7_75t_L g636 ( .A(n_578), .Y(n_636) );
AND2x4_ASAP7_75t_L g588 ( .A(n_579), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g662 ( .A(n_579), .B(n_601), .Y(n_662) );
INVx1_ASAP7_75t_L g689 ( .A(n_579), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_579), .B(n_676), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_580), .B(n_650), .Y(n_670) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_581), .B(n_603), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_581), .B(n_650), .Y(n_749) );
INVx1_ASAP7_75t_L g760 ( .A(n_582), .Y(n_760) );
A2O1A1Ixp33_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_587), .B(n_590), .C(n_598), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g602 ( .A(n_586), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g640 ( .A(n_586), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g622 ( .A(n_587), .Y(n_622) );
AND2x2_ASAP7_75t_L g599 ( .A(n_588), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_588), .B(n_650), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_588), .B(n_669), .Y(n_693) );
OR2x2_ASAP7_75t_L g609 ( .A(n_589), .B(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g641 ( .A(n_589), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_589), .B(n_601), .Y(n_656) );
AND2x2_ASAP7_75t_L g713 ( .A(n_589), .B(n_669), .Y(n_713) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_589), .Y(n_720) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AOI221xp5_ASAP7_75t_L g724 ( .A1(n_591), .A2(n_603), .B1(n_725), .B2(n_727), .C(n_730), .Y(n_724) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_595), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g614 ( .A(n_594), .B(n_597), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_594), .B(n_664), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_594), .B(n_621), .Y(n_729) );
INVx1_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g714 ( .A(n_596), .B(n_715), .Y(n_714) );
OR2x2_ASAP7_75t_L g728 ( .A(n_596), .B(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_597), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g625 ( .A(n_597), .B(n_618), .Y(n_625) );
AND2x2_ASAP7_75t_L g695 ( .A(n_597), .B(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_597), .B(n_644), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_597), .B(n_745), .Y(n_744) );
OAI21xp5_ASAP7_75t_SL g598 ( .A1(n_599), .A2(n_602), .B(n_604), .Y(n_598) );
INVx2_ASAP7_75t_L g631 ( .A(n_599), .Y(n_631) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g651 ( .A(n_601), .Y(n_651) );
OR2x2_ASAP7_75t_L g655 ( .A(n_603), .B(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g758 ( .A(n_603), .B(n_726), .Y(n_758) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
AOI21xp33_ASAP7_75t_SL g608 ( .A1(n_609), .A2(n_611), .B(n_613), .Y(n_608) );
INVx1_ASAP7_75t_L g762 ( .A(n_609), .Y(n_762) );
INVx2_ASAP7_75t_SL g676 ( .A(n_610), .Y(n_676) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
A2O1A1Ixp33_ASAP7_75t_L g757 ( .A1(n_613), .A2(n_694), .B(n_758), .C(n_759), .Y(n_757) );
OAI322xp33_ASAP7_75t_SL g626 ( .A1(n_614), .A2(n_627), .A3(n_630), .B1(n_631), .B2(n_632), .C1(n_634), .C2(n_637), .Y(n_626) );
INVx2_ASAP7_75t_L g646 ( .A(n_614), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_622), .B1(n_623), .B2(n_625), .C(n_626), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OAI22xp33_ASAP7_75t_SL g692 ( .A1(n_617), .A2(n_693), .B1(n_694), .B2(n_697), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_618), .B(n_621), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_618), .B(n_756), .Y(n_755) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g691 ( .A(n_620), .B(n_653), .Y(n_691) );
INVx1_ASAP7_75t_L g681 ( .A(n_621), .Y(n_681) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_625), .A2(n_735), .B(n_737), .Y(n_734) );
AOI21xp33_ASAP7_75t_L g659 ( .A1(n_627), .A2(n_660), .B(n_663), .Y(n_659) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NOR2xp67_ASAP7_75t_SL g688 ( .A(n_629), .B(n_689), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_629), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g745 ( .A(n_630), .Y(n_745) );
INVx1_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND4xp25_ASAP7_75t_L g638 ( .A(n_639), .B(n_666), .C(n_682), .D(n_698), .Y(n_638) );
AOI211xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_642), .B(n_647), .C(n_659), .Y(n_639) );
INVx1_ASAP7_75t_L g731 ( .A(n_640), .Y(n_731) );
AND2x2_ASAP7_75t_L g679 ( .A(n_641), .B(n_662), .Y(n_679) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_646), .B(n_681), .Y(n_680) );
OAI22xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_652), .B1(n_655), .B2(n_657), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_649), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g697 ( .A(n_650), .Y(n_697) );
O2A1O1Ixp33_ASAP7_75t_L g711 ( .A1(n_650), .A2(n_689), .B(n_712), .C(n_714), .Y(n_711) );
OR2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_L g696 ( .A(n_653), .Y(n_696) );
INVx1_ASAP7_75t_L g756 ( .A(n_654), .Y(n_756) );
NAND2xp33_ASAP7_75t_SL g746 ( .A(n_655), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g685 ( .A(n_664), .Y(n_685) );
O2A1O1Ixp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_670), .B(n_671), .C(n_673), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .B1(n_678), .B2(n_680), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_676), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_681), .B(n_702), .Y(n_764) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AOI21xp33_ASAP7_75t_SL g686 ( .A1(n_687), .A2(n_690), .B(n_691), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_704), .B1(n_707), .B2(n_709), .C(n_711), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVxp67_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_714), .A2(n_731), .B1(n_732), .B2(n_733), .Y(n_730) );
NAND3xp33_ASAP7_75t_SL g716 ( .A(n_717), .B(n_724), .C(n_734), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
CKINVDCx16_ASAP7_75t_R g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVxp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OAI211xp5_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_742), .B(n_743), .C(n_752), .Y(n_740) );
INVx1_ASAP7_75t_L g761 ( .A(n_741), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_746), .B1(n_748), .B2(n_750), .Y(n_743) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_761), .B1(n_762), .B2(n_763), .Y(n_759) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
OAI22x1_ASAP7_75t_SL g765 ( .A1(n_766), .A2(n_767), .B1(n_768), .B2(n_769), .Y(n_765) );
endmodule