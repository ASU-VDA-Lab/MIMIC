module fake_jpeg_4575_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_19),
.Y(n_66)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_25),
.B(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_17),
.B1(n_27),
.B2(n_21),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_54),
.B1(n_62),
.B2(n_72),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_33),
.B1(n_23),
.B2(n_25),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_50),
.A2(n_53),
.B1(n_56),
.B2(n_59),
.Y(n_96)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_55),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_33),
.B1(n_23),
.B2(n_25),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_45),
.B1(n_41),
.B2(n_35),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_33),
.B1(n_23),
.B2(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_67),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_33),
.B1(n_32),
.B2(n_16),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_34),
.A2(n_16),
.B1(n_17),
.B2(n_21),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_27),
.Y(n_91)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_38),
.B(n_22),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_29),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_38),
.A2(n_16),
.B1(n_17),
.B2(n_21),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_77),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_32),
.B1(n_18),
.B2(n_19),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

AOI22x1_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_28),
.B1(n_38),
.B2(n_30),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_79),
.A2(n_85),
.B1(n_94),
.B2(n_58),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_81),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_84),
.Y(n_114)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_32),
.B1(n_29),
.B2(n_22),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_22),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_89),
.Y(n_100)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_98),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_19),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_38),
.Y(n_90)
);

OAI32xp33_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_79),
.A3(n_82),
.B1(n_97),
.B2(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_93),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_18),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_63),
.A2(n_27),
.B1(n_18),
.B2(n_20),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_0),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_97),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_57),
.B(n_1),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_63),
.B1(n_71),
.B2(n_52),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_99),
.A2(n_106),
.B1(n_58),
.B2(n_96),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_101),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_104),
.Y(n_136)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_107),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_79),
.A2(n_71),
.B1(n_52),
.B2(n_51),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_108),
.A2(n_73),
.B(n_48),
.Y(n_138)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_110),
.B(n_111),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_80),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_92),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_112),
.Y(n_142)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_113),
.B(n_117),
.Y(n_139)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_92),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_119),
.Y(n_140)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_52),
.B1(n_47),
.B2(n_58),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_120),
.A2(n_121),
.B1(n_78),
.B2(n_90),
.Y(n_130)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_86),
.Y(n_143)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_128),
.A2(n_131),
.B1(n_148),
.B2(n_149),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_103),
.A2(n_90),
.B(n_94),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_100),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_130),
.A2(n_132),
.B1(n_145),
.B2(n_146),
.Y(n_176)
);

AO22x1_ASAP7_75t_SL g131 ( 
.A1(n_121),
.A2(n_102),
.B1(n_108),
.B2(n_99),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_78),
.B1(n_84),
.B2(n_48),
.Y(n_132)
);

BUFx12_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_137),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_116),
.A2(n_67),
.B1(n_84),
.B2(n_98),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_114),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_73),
.C(n_86),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_129),
.C(n_140),
.Y(n_168)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_120),
.A2(n_81),
.B1(n_83),
.B2(n_32),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_108),
.A2(n_83),
.B1(n_32),
.B2(n_69),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_106),
.A2(n_69),
.B(n_65),
.C(n_30),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_147),
.A2(n_153),
.B(n_123),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_113),
.A2(n_32),
.B1(n_69),
.B2(n_65),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_65),
.B1(n_88),
.B2(n_74),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_150),
.B(n_109),
.Y(n_158)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_107),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_SL g153 ( 
.A1(n_112),
.A2(n_30),
.B(n_24),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_151),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_163),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_103),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_157),
.A2(n_172),
.B(n_139),
.Y(n_197)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_146),
.B(n_124),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_166),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_124),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_170),
.Y(n_195)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_151),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_164),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_119),
.B1(n_104),
.B2(n_118),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_165),
.A2(n_132),
.B1(n_130),
.B2(n_134),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_173),
.C(n_175),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_169),
.A2(n_134),
.B1(n_147),
.B2(n_142),
.Y(n_187)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_171),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_114),
.B(n_111),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_131),
.B(n_126),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_110),
.C(n_122),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_184),
.C(n_159),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_136),
.B(n_101),
.Y(n_178)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_135),
.Y(n_183)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_131),
.B(n_123),
.C(n_46),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_185),
.A2(n_186),
.B1(n_191),
.B2(n_205),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_181),
.A2(n_134),
.B1(n_142),
.B2(n_144),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_187),
.A2(n_190),
.B1(n_201),
.B2(n_207),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_128),
.B1(n_147),
.B2(n_144),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_123),
.Y(n_191)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_165),
.A2(n_139),
.B(n_148),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_197),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_198),
.B(n_204),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_184),
.A2(n_145),
.B1(n_153),
.B2(n_155),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_164),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_161),
.A2(n_155),
.B1(n_133),
.B2(n_105),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_209),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_172),
.A2(n_133),
.B1(n_137),
.B2(n_46),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_133),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_208),
.A2(n_157),
.B1(n_182),
.B2(n_180),
.Y(n_216)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_175),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_157),
.C(n_161),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_177),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_211),
.Y(n_227)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_221),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_163),
.Y(n_215)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_215),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_228),
.Y(n_242)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_217),
.B(n_218),
.Y(n_238)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_222),
.C(n_224),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_162),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_166),
.C(n_162),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_171),
.C(n_170),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_231),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_169),
.C(n_183),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_229),
.B(n_233),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_167),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_235),
.Y(n_246)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_199),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_232),
.Y(n_253)
);

NOR4xp25_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_167),
.C(n_133),
.D(n_15),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_185),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_234),
.B(n_236),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_202),
.B(n_26),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_190),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_30),
.Y(n_259)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_240),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_226),
.A2(n_209),
.B1(n_197),
.B2(n_191),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_241),
.A2(n_250),
.B1(n_237),
.B2(n_214),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_227),
.B(n_188),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_244),
.B(n_245),
.Y(n_269)
);

FAx1_ASAP7_75t_SL g245 ( 
.A(n_216),
.B(n_208),
.CI(n_191),
.CON(n_245),
.SN(n_245)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_203),
.B(n_193),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_249),
.A2(n_259),
.B(n_24),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_212),
.A2(n_203),
.B1(n_198),
.B2(n_193),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_214),
.A2(n_188),
.B1(n_194),
.B2(n_115),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_251),
.A2(n_30),
.B1(n_24),
.B2(n_20),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_220),
.B(n_194),
.Y(n_252)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_26),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_258),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_213),
.B(n_15),
.Y(n_255)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_224),
.B(n_222),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_256),
.B(n_14),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_26),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_253),
.B(n_219),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_261),
.B(n_249),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_262),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_263),
.A2(n_277),
.B(n_248),
.Y(n_285)
);

AOI321xp33_ASAP7_75t_L g264 ( 
.A1(n_245),
.A2(n_230),
.A3(n_215),
.B1(n_221),
.B2(n_235),
.C(n_212),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_264),
.A2(n_278),
.B(n_13),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_228),
.C(n_115),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_273),
.C(n_279),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_26),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_274),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_250),
.A2(n_257),
.B1(n_247),
.B2(n_238),
.Y(n_267)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_267),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_268),
.A2(n_76),
.B1(n_24),
.B2(n_20),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_260),
.A2(n_245),
.B1(n_239),
.B2(n_241),
.Y(n_272)
);

A2O1A1Ixp33_ASAP7_75t_SL g286 ( 
.A1(n_272),
.A2(n_257),
.B(n_248),
.C(n_246),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_242),
.B(n_26),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_26),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_76),
.C(n_24),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_275),
.A2(n_260),
.B1(n_258),
.B2(n_254),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_291),
.C(n_295),
.Y(n_304)
);

BUFx24_ASAP7_75t_SL g283 ( 
.A(n_276),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_292),
.Y(n_299)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_284),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_285),
.A2(n_290),
.B(n_293),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_286),
.A2(n_274),
.B(n_271),
.Y(n_305)
);

OAI321xp33_ASAP7_75t_L g309 ( 
.A1(n_287),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_20),
.B1(n_2),
.B2(n_3),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_268),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_26),
.C(n_2),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_263),
.A2(n_13),
.B(n_2),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_294),
.A2(n_1),
.B(n_3),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_270),
.A2(n_13),
.B1(n_2),
.B2(n_3),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_266),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_308),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g297 ( 
.A(n_281),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_297),
.A2(n_305),
.B1(n_286),
.B2(n_282),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_299),
.B(n_303),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_301),
.B(n_306),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_290),
.A2(n_264),
.B1(n_273),
.B2(n_279),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_307),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_291),
.B(n_271),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_286),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_1),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_309),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_319)
);

NOR2x1_ASAP7_75t_L g310 ( 
.A(n_307),
.B(n_300),
.Y(n_310)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_310),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_319),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_286),
.C(n_5),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_7),
.C(n_8),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_4),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_314),
.B(n_320),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_4),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_316),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_297),
.B(n_5),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_321),
.A2(n_324),
.B(n_12),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_323),
.B(n_324),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_9),
.C(n_11),
.Y(n_324)
);

INVx11_ASAP7_75t_L g325 ( 
.A(n_310),
.Y(n_325)
);

AO21x1_ASAP7_75t_L g330 ( 
.A1(n_325),
.A2(n_312),
.B(n_311),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_9),
.C(n_11),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_326),
.A2(n_11),
.B(n_12),
.Y(n_332)
);

AOI21xp33_ASAP7_75t_L g335 ( 
.A1(n_329),
.A2(n_330),
.B(n_331),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_322),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_332),
.Y(n_334)
);

AOI222xp33_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_325),
.B1(n_327),
.B2(n_317),
.C1(n_318),
.C2(n_328),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_321),
.C(n_333),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_337),
.B(n_316),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_334),
.Y(n_339)
);


endmodule