module fake_jpeg_30828_n_139 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_139);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_63),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_0),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_22),
.C(n_41),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_44),
.C(n_59),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_58),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_68),
.Y(n_70)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_67),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_1),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVxp67_ASAP7_75t_SL g77 ( 
.A(n_69),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_72),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_56),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_75),
.B(n_78),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_54),
.B1(n_51),
.B2(n_55),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_49),
.Y(n_78)
);

BUFx16f_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_65),
.B1(n_47),
.B2(n_46),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_83),
.A2(n_91),
.B1(n_15),
.B2(n_16),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_81),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_29),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_79),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_87),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_86),
.B(n_94),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_79),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_43),
.B1(n_2),
.B2(n_3),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_77),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_4),
.B(n_5),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_10),
.B(n_11),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_96),
.A2(n_17),
.B1(n_21),
.B2(n_23),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_70),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_10),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_104),
.B(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_82),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_14),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_108),
.A2(n_109),
.B1(n_100),
.B2(n_114),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_24),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_110),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_98),
.B(n_42),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_114),
.A2(n_88),
.B1(n_32),
.B2(n_33),
.Y(n_117)
);

INVxp33_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_101),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_98),
.B1(n_35),
.B2(n_36),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_121),
.C(n_114),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_31),
.C(n_39),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_122),
.B(n_109),
.Y(n_126)
);

INVxp33_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_102),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_129),
.B1(n_120),
.B2(n_124),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_128),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_130),
.A2(n_131),
.B1(n_123),
.B2(n_108),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_125),
.C(n_111),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_132),
.B1(n_131),
.B2(n_116),
.Y(n_135)
);

INVxp33_ASAP7_75t_SL g136 ( 
.A(n_135),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_116),
.C(n_118),
.Y(n_137)
);

OAI21x1_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_118),
.B(n_113),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_113),
.B(n_99),
.Y(n_139)
);


endmodule