module fake_jpeg_27842_n_43 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx4_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx5_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

AND2x2_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_6),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_15),
.A2(n_18),
.B(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_17),
.Y(n_23)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_0),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_19),
.A2(n_12),
.B1(n_13),
.B2(n_9),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_5),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_12),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_24),
.A2(n_23),
.B1(n_27),
.B2(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_25),
.B(n_28),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_11),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_30),
.Y(n_32)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_11),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_18),
.B(n_22),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_32),
.B(n_36),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_9),
.B1(n_17),
.B2(n_20),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_34),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_20),
.C(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_32),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_31),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_39),
.A2(n_40),
.B1(n_34),
.B2(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_42),
.Y(n_43)
);


endmodule