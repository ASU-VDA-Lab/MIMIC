module fake_jpeg_26071_n_311 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_311);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_145;
wire n_20;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_6),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_15),
.B1(n_23),
.B2(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_36),
.Y(n_64)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_55),
.Y(n_92)
);

CKINVDCx12_ASAP7_75t_R g54 ( 
.A(n_47),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx5_ASAP7_75t_SL g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_15),
.B1(n_29),
.B2(n_28),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_28),
.B1(n_37),
.B2(n_45),
.Y(n_83)
);

CKINVDCx12_ASAP7_75t_R g58 ( 
.A(n_50),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_58),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_29),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_30),
.Y(n_74)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_33),
.C(n_27),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_36),
.Y(n_96)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_33),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_65),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_34),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_69),
.B(n_73),
.Y(n_78)
);

CKINVDCx9p33_ASAP7_75t_R g71 ( 
.A(n_41),
.Y(n_71)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

CKINVDCx12_ASAP7_75t_R g72 ( 
.A(n_50),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_49),
.B1(n_46),
.B2(n_37),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_34),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_74),
.B(n_21),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_32),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_90),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_95),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_55),
.B1(n_48),
.B2(n_45),
.Y(n_103)
);

NAND2xp33_ASAP7_75t_SL g85 ( 
.A(n_71),
.B(n_27),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_88),
.B(n_68),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_86),
.Y(n_120)
);

AOI32xp33_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_49),
.A3(n_46),
.B1(n_37),
.B2(n_28),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_59),
.A2(n_45),
.B1(n_48),
.B2(n_25),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_55),
.B1(n_70),
.B2(n_52),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_31),
.Y(n_90)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_63),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_91),
.C(n_79),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_78),
.B(n_65),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_99),
.B(n_100),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_65),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_62),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_101),
.B(n_104),
.Y(n_146)
);

AO21x1_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_95),
.B(n_91),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_103),
.A2(n_38),
.B1(n_39),
.B2(n_21),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_61),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_53),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_105),
.B(n_109),
.Y(n_134)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_107),
.A2(n_39),
.B1(n_26),
.B2(n_24),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_32),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_114),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_93),
.A2(n_52),
.B1(n_70),
.B2(n_67),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_112),
.A2(n_113),
.B1(n_87),
.B2(n_84),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_67),
.B1(n_30),
.B2(n_31),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_118),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_85),
.A2(n_67),
.B1(n_72),
.B2(n_58),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_36),
.Y(n_117)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_75),
.B(n_54),
.Y(n_122)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

FAx1_ASAP7_75t_SL g123 ( 
.A(n_98),
.B(n_91),
.CI(n_75),
.CON(n_123),
.SN(n_123)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_125),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_128),
.A2(n_133),
.B(n_138),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_108),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_129),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_141),
.C(n_97),
.Y(n_161)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_135),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_84),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_121),
.A2(n_120),
.B1(n_111),
.B2(n_114),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_142),
.B1(n_153),
.B2(n_154),
.Y(n_155)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_148),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_120),
.A2(n_79),
.B1(n_94),
.B2(n_82),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_140),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_77),
.C(n_35),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_100),
.A2(n_87),
.B1(n_94),
.B2(n_38),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_145),
.Y(n_187)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_150),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_99),
.A2(n_22),
.B1(n_16),
.B2(n_23),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_119),
.B(n_109),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_156),
.A2(n_143),
.B(n_147),
.Y(n_190)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_157),
.B(n_160),
.Y(n_212)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_164),
.C(n_180),
.Y(n_203)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_123),
.C(n_141),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_169),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_97),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_175),
.Y(n_206)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_170),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_134),
.B(n_106),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_171),
.Y(n_207)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_181),
.Y(n_198)
);

INVxp33_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_35),
.Y(n_175)
);

OA22x2_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_115),
.B1(n_108),
.B2(n_39),
.Y(n_176)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_124),
.A2(n_6),
.B(n_1),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_179),
.A2(n_185),
.B(n_12),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_123),
.B(n_35),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_135),
.B(n_44),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_148),
.A2(n_20),
.B1(n_17),
.B2(n_19),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_183),
.A2(n_26),
.B1(n_24),
.B2(n_12),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_140),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_184),
.Y(n_195)
);

AND2x6_ASAP7_75t_L g185 ( 
.A(n_124),
.B(n_11),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_127),
.B(n_18),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_186),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_190),
.A2(n_202),
.B(n_204),
.Y(n_216)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_197),
.Y(n_215)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_137),
.Y(n_199)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_166),
.A2(n_132),
.B1(n_126),
.B2(n_138),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_201),
.A2(n_208),
.B1(n_211),
.B2(n_213),
.Y(n_225)
);

NOR2xp67_ASAP7_75t_SL g202 ( 
.A(n_174),
.B(n_142),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_174),
.A2(n_126),
.B(n_152),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_209),
.A2(n_163),
.B(n_177),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_161),
.B(n_56),
.C(n_25),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_164),
.C(n_175),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_187),
.A2(n_26),
.B1(n_24),
.B2(n_21),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_177),
.A2(n_20),
.B1(n_19),
.B2(n_17),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_217),
.A2(n_190),
.B(n_198),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_221),
.C(n_229),
.Y(n_248)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_212),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_233),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_196),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_180),
.C(n_168),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_207),
.A2(n_158),
.B1(n_179),
.B2(n_185),
.Y(n_222)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_156),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_228),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_192),
.A2(n_155),
.B1(n_176),
.B2(n_159),
.Y(n_224)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_192),
.A2(n_176),
.B1(n_160),
.B2(n_173),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_226),
.A2(n_227),
.B1(n_234),
.B2(n_191),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_195),
.A2(n_176),
.B1(n_170),
.B2(n_20),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_206),
.B(n_18),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_206),
.C(n_197),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_198),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_231),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_56),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_189),
.B(n_56),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_232),
.B(n_200),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_25),
.C(n_18),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_195),
.A2(n_19),
.B1(n_17),
.B2(n_12),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_235),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_217),
.A2(n_204),
.B(n_193),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_236),
.B(n_228),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_241),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_238),
.A2(n_244),
.B(n_246),
.Y(n_259)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_214),
.A2(n_199),
.B1(n_188),
.B2(n_191),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_25),
.B1(n_1),
.B2(n_2),
.Y(n_263)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_231),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_188),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_250),
.Y(n_254)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_247),
.B(n_252),
.Y(n_257)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_194),
.Y(n_252)
);

OAI21x1_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_236),
.B(n_216),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_249),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_240),
.A2(n_200),
.B1(n_205),
.B2(n_194),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_261),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_241),
.A2(n_229),
.B1(n_218),
.B2(n_221),
.Y(n_256)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_239),
.A2(n_201),
.B1(n_223),
.B2(n_205),
.Y(n_260)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_260),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_243),
.B(n_213),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_251),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_265),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_0),
.C(n_1),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_267),
.C(n_246),
.Y(n_269)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_0),
.C(n_11),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_262),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_277),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_259),
.A2(n_252),
.B(n_235),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_276),
.B(n_257),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_251),
.C(n_242),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_275),
.A2(n_280),
.B(n_267),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_249),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_244),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_259),
.A2(n_6),
.B(n_2),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_278),
.A2(n_3),
.B(n_4),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_0),
.C(n_11),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_268),
.Y(n_291)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_277),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_280),
.Y(n_297)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_283),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_285),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_274),
.A2(n_258),
.B1(n_264),
.B2(n_263),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_286),
.B(n_288),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_7),
.B1(n_3),
.B2(n_4),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_7),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_289),
.B(n_290),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_281),
.C(n_269),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_279),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_292),
.A2(n_297),
.B(n_287),
.Y(n_300)
);

AOI21x1_ASAP7_75t_L g294 ( 
.A1(n_287),
.A2(n_284),
.B(n_270),
.Y(n_294)
);

NAND2xp33_ASAP7_75t_SL g302 ( 
.A(n_294),
.B(n_298),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_299),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_300),
.A2(n_301),
.B(n_302),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_295),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_301)
);

OA21x2_ASAP7_75t_SL g303 ( 
.A1(n_293),
.A2(n_5),
.B(n_8),
.Y(n_303)
);

OAI21x1_ASAP7_75t_L g306 ( 
.A1(n_304),
.A2(n_298),
.B(n_305),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_296),
.C(n_303),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_10),
.B(n_9),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_9),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_9),
.B1(n_10),
.B2(n_0),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_0),
.B1(n_10),
.B2(n_282),
.Y(n_311)
);


endmodule