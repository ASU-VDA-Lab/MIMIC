module real_jpeg_18331_n_15 (n_108, n_8, n_116, n_0, n_111, n_2, n_10, n_114, n_9, n_12, n_6, n_11, n_14, n_110, n_112, n_7, n_117, n_3, n_119, n_5, n_4, n_109, n_115, n_1, n_118, n_13, n_113, n_15);

input n_108;
input n_8;
input n_116;
input n_0;
input n_111;
input n_2;
input n_10;
input n_114;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_110;
input n_112;
input n_7;
input n_117;
input n_3;
input n_119;
input n_5;
input n_4;
input n_109;
input n_115;
input n_1;
input n_118;
input n_13;
input n_113;

output n_15;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_0),
.B(n_30),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_1),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_1),
.B(n_35),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_2),
.B(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_2),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_3),
.B(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_3),
.Y(n_98)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_SL g73 ( 
.A(n_4),
.B(n_62),
.C(n_69),
.Y(n_73)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_5),
.B(n_42),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_7),
.B(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_8),
.A2(n_60),
.B(n_72),
.Y(n_59)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_8),
.Y(n_74)
);

MAJx2_ASAP7_75t_L g57 ( 
.A(n_9),
.B(n_58),
.C(n_86),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_10),
.Y(n_102)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

AOI322xp5_ASAP7_75t_SL g93 ( 
.A1(n_11),
.A2(n_39),
.A3(n_50),
.B1(n_53),
.B2(n_94),
.C1(n_96),
.C2(n_119),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_12),
.A2(n_17),
.B1(n_18),
.B2(n_23),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_14),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_24),
.Y(n_15)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_20),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_99),
.B(n_104),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI31xp67_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.A3(n_57),
.B(n_90),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_43),
.Y(n_42)
);

NOR3xp33_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_38),
.C(n_44),
.Y(n_33)
);

NOR3xp33_ASAP7_75t_L g94 ( 
.A(n_34),
.B(n_46),
.C(n_95),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

OAI321xp33_ASAP7_75t_L g90 ( 
.A1(n_38),
.A2(n_44),
.A3(n_91),
.B1(n_92),
.B2(n_93),
.C(n_118),
.Y(n_90)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_50),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_56),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_80),
.C(n_81),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_67),
.C(n_68),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B(n_75),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_108),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_109),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_110),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_111),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_112),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_113),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_114),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_115),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_116),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_117),
.Y(n_87)
);


endmodule