module fake_jpeg_10024_n_247 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_14),
.B(n_4),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_29),
.Y(n_49)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx2_ASAP7_75t_SL g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_27),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_38),
.Y(n_65)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

CKINVDCx6p67_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_42),
.Y(n_52)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_55),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_24),
.B1(n_18),
.B2(n_28),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_60),
.B(n_27),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_20),
.Y(n_47)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_30),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_54),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_21),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_19),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_22),
.C(n_23),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_40),
.B(n_28),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_58),
.Y(n_82)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_18),
.B1(n_24),
.B2(n_30),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_26),
.B1(n_42),
.B2(n_21),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_35),
.A2(n_39),
.B1(n_36),
.B2(n_25),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_61),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_36),
.B(n_25),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_29),
.Y(n_85)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_68),
.Y(n_87)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_81),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_39),
.B1(n_42),
.B2(n_31),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_70),
.A2(n_72),
.B1(n_76),
.B2(n_45),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_71),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_39),
.B1(n_31),
.B2(n_35),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_75),
.Y(n_98)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_80),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_84),
.Y(n_102)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_85),
.B(n_48),
.Y(n_89)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_91),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_89),
.B(n_92),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_54),
.C(n_55),
.Y(n_90)
);

XNOR2x1_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_107),
.Y(n_110)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_82),
.B(n_48),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_67),
.B(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_94),
.B(n_99),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_101),
.B1(n_65),
.B2(n_80),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_86),
.B(n_57),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_103),
.Y(n_118)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_71),
.A2(n_43),
.B1(n_42),
.B2(n_52),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_67),
.B(n_15),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_44),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_106),
.Y(n_123)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_58),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_74),
.B(n_52),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_59),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_73),
.B(n_65),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_112),
.B(n_116),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_117),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_105),
.A2(n_76),
.B1(n_73),
.B2(n_68),
.Y(n_114)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_102),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_120),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_104),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_127),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_69),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_132),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_98),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_129),
.Y(n_151)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_94),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_93),
.A2(n_83),
.B1(n_41),
.B2(n_32),
.Y(n_131)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_37),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_95),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_139),
.C(n_143),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_124),
.B(n_97),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_136),
.B(n_145),
.Y(n_167)
);

NOR2xp67_ASAP7_75t_R g137 ( 
.A(n_122),
.B(n_92),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_149),
.B(n_122),
.Y(n_162)
);

XOR2x1_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_89),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_138),
.B(n_142),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_95),
.C(n_107),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_123),
.A2(n_108),
.B(n_96),
.Y(n_142)
);

MAJx2_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_95),
.C(n_107),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_146),
.B(n_147),
.Y(n_173)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_125),
.A2(n_107),
.B(n_88),
.Y(n_149)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_125),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_121),
.C(n_129),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_120),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_144),
.Y(n_156)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_144),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_157),
.A2(n_159),
.B1(n_133),
.B2(n_140),
.Y(n_179)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_160),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_147),
.A2(n_115),
.B1(n_121),
.B2(n_116),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_162),
.B(n_137),
.Y(n_184)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_170),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_139),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_165),
.C(n_169),
.Y(n_177)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_168),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_117),
.C(n_118),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_112),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_135),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_172),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_124),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_127),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_146),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_179),
.A2(n_77),
.B1(n_26),
.B2(n_91),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_155),
.B(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_138),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_189),
.C(n_190),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_174),
.Y(n_183)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_191),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_148),
.B(n_149),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_185),
.A2(n_103),
.B(n_21),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_143),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_169),
.Y(n_194)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_161),
.C(n_165),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_133),
.C(n_145),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_162),
.B(n_118),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_178),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_192),
.A2(n_205),
.B(n_77),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_157),
.B1(n_173),
.B2(n_159),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_193),
.A2(n_196),
.B1(n_180),
.B2(n_187),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_204),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_158),
.B1(n_163),
.B2(n_172),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_197),
.A2(n_191),
.B1(n_183),
.B2(n_84),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_0),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_199),
.A2(n_2),
.B(n_3),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_184),
.A2(n_0),
.B(n_1),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_203),
.A2(n_1),
.B(n_2),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_189),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_206),
.B(n_207),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_209),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_200),
.A2(n_202),
.B1(n_195),
.B2(n_199),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_210),
.A2(n_212),
.B1(n_214),
.B2(n_201),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_211),
.A2(n_3),
.B(n_6),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_203),
.A2(n_177),
.B1(n_182),
.B2(n_5),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_201),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_41),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_198),
.A2(n_62),
.B1(n_50),
.B2(n_29),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_198),
.A2(n_2),
.B(n_3),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_215),
.A2(n_216),
.B(n_19),
.Y(n_221)
);

OA21x2_ASAP7_75t_L g216 ( 
.A1(n_194),
.A2(n_62),
.B(n_50),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_220),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_215),
.A2(n_204),
.B1(n_7),
.B2(n_8),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_9),
.C(n_10),
.Y(n_233)
);

BUFx24_ASAP7_75t_SL g224 ( 
.A(n_217),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_216),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_225),
.A2(n_226),
.B(n_8),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_213),
.A2(n_6),
.B(n_8),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_217),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_227),
.A2(n_9),
.B(n_11),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_230),
.B(n_233),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_221),
.A2(n_216),
.B1(n_211),
.B2(n_208),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_231),
.A2(n_12),
.B1(n_19),
.B2(n_29),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_12),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_229),
.A2(n_228),
.B1(n_230),
.B2(n_218),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_237),
.C(n_12),
.Y(n_239)
);

NAND3xp33_ASAP7_75t_SL g240 ( 
.A(n_236),
.B(n_50),
.C(n_62),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_238),
.B(n_32),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_239),
.A2(n_241),
.B(n_242),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_240),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_41),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_244),
.A2(n_235),
.B1(n_37),
.B2(n_41),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_246),
.Y(n_247)
);

O2A1O1Ixp33_ASAP7_75t_SL g246 ( 
.A1(n_243),
.A2(n_32),
.B(n_37),
.C(n_244),
.Y(n_246)
);


endmodule