module real_aes_7335_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_800;
wire n_778;
wire n_618;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_284;
wire n_656;
wire n_532;
wire n_316;
wire n_746;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_293;
wire n_397;
wire n_358;
wire n_275;
wire n_385;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_720;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_279;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_842;
wire n_475;
wire n_554;
wire n_798;
wire n_797;
wire n_668;
CKINVDCx20_ASAP7_75t_R g390 ( .A(n_0), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_1), .Y(n_797) );
XOR2x2_ASAP7_75t_L g522 ( .A(n_2), .B(n_523), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_3), .A2(n_16), .B1(n_403), .B2(n_406), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_4), .A2(n_225), .B1(n_341), .B2(n_344), .Y(n_652) );
INVx1_ASAP7_75t_L g316 ( .A(n_5), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_6), .A2(n_59), .B1(n_526), .B2(n_568), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_7), .A2(n_177), .B1(n_472), .B2(n_517), .Y(n_814) );
AOI22xp33_ASAP7_75t_SL g839 ( .A1(n_8), .A2(n_104), .B1(n_337), .B2(n_404), .Y(n_839) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_9), .A2(n_111), .B1(n_341), .B2(n_344), .C(n_347), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_10), .A2(n_377), .B1(n_422), .B2(n_423), .Y(n_376) );
INVx1_ASAP7_75t_L g422 ( .A(n_10), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_11), .A2(n_244), .B1(n_326), .B2(n_465), .Y(n_464) );
AOI222xp33_ASAP7_75t_L g542 ( .A1(n_12), .A2(n_30), .B1(n_215), .B2(n_360), .C1(n_543), .C2(n_545), .Y(n_542) );
AOI22xp33_ASAP7_75t_SL g595 ( .A1(n_13), .A2(n_169), .B1(n_289), .B2(n_532), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_14), .A2(n_139), .B1(n_461), .B2(n_597), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_15), .A2(n_71), .B1(n_305), .B2(n_534), .Y(n_533) );
AOI221xp5_ASAP7_75t_L g691 ( .A1(n_17), .A2(n_26), .B1(n_443), .B2(n_461), .C(n_692), .Y(n_691) );
AOI22xp33_ASAP7_75t_SL g626 ( .A1(n_18), .A2(n_217), .B1(n_627), .B2(n_628), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g320 ( .A1(n_19), .A2(n_234), .B1(n_321), .B2(n_326), .C(n_330), .Y(n_320) );
INVx1_ASAP7_75t_L g348 ( .A(n_20), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g287 ( .A1(n_21), .A2(n_69), .B1(n_288), .B2(n_305), .C(n_309), .Y(n_287) );
AOI222xp33_ASAP7_75t_L g359 ( .A1(n_22), .A2(n_34), .B1(n_247), .B2(n_360), .C1(n_362), .C2(n_366), .Y(n_359) );
XOR2x2_ASAP7_75t_L g486 ( .A(n_23), .B(n_487), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_24), .A2(n_73), .B1(n_404), .B2(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g573 ( .A(n_25), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_27), .A2(n_91), .B1(n_545), .B2(n_649), .Y(n_715) );
AO22x2_ASAP7_75t_L g302 ( .A1(n_28), .A2(n_81), .B1(n_294), .B2(n_299), .Y(n_302) );
INVx1_ASAP7_75t_L g789 ( .A(n_28), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_29), .A2(n_43), .B1(n_321), .B2(n_512), .Y(n_840) );
AOI22xp33_ASAP7_75t_SL g619 ( .A1(n_31), .A2(n_33), .B1(n_403), .B2(n_540), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_32), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_35), .A2(n_174), .B1(n_493), .B2(n_545), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_36), .A2(n_178), .B1(n_367), .B2(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_SL g616 ( .A1(n_37), .A2(n_63), .B1(n_478), .B2(n_584), .Y(n_616) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_38), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_39), .A2(n_40), .B1(n_526), .B2(n_527), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_41), .A2(n_52), .B1(n_288), .B2(n_560), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_42), .A2(n_202), .B1(n_329), .B2(n_532), .Y(n_554) );
AO22x2_ASAP7_75t_L g304 ( .A1(n_44), .A2(n_85), .B1(n_294), .B2(n_295), .Y(n_304) );
INVx1_ASAP7_75t_L g790 ( .A(n_44), .Y(n_790) );
AOI22xp33_ASAP7_75t_SL g722 ( .A1(n_45), .A2(n_48), .B1(n_337), .B2(n_510), .Y(n_722) );
AOI22xp33_ASAP7_75t_SL g717 ( .A1(n_46), .A2(n_117), .B1(n_305), .B2(n_718), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_47), .Y(n_803) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_49), .A2(n_268), .B1(n_514), .B2(n_562), .C(n_686), .Y(n_685) );
AOI22xp33_ASAP7_75t_SL g711 ( .A1(n_50), .A2(n_257), .B1(n_392), .B2(n_543), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_51), .A2(n_143), .B1(n_416), .B2(n_420), .Y(n_415) );
AOI22xp33_ASAP7_75t_SL g660 ( .A1(n_53), .A2(n_142), .B1(n_403), .B2(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_54), .B(n_526), .Y(n_586) );
INVx1_ASAP7_75t_L g452 ( .A(n_55), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_56), .A2(n_228), .B1(n_520), .B2(n_521), .Y(n_519) );
AOI22xp5_ASAP7_75t_SL g555 ( .A1(n_57), .A2(n_255), .B1(n_472), .B2(n_556), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_58), .A2(n_118), .B1(n_413), .B2(n_414), .Y(n_412) );
INVx1_ASAP7_75t_L g693 ( .A(n_60), .Y(n_693) );
AOI22xp33_ASAP7_75t_SL g719 ( .A1(n_61), .A2(n_194), .B1(n_420), .B2(n_720), .Y(n_719) );
XOR2x2_ASAP7_75t_L g706 ( .A(n_62), .B(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_64), .B(n_501), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_65), .A2(n_86), .B1(n_321), .B2(n_409), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_66), .A2(n_201), .B1(n_289), .B2(n_445), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_67), .A2(n_249), .B1(n_496), .B2(n_504), .Y(n_569) );
OA22x2_ASAP7_75t_L g639 ( .A1(n_68), .A2(n_640), .B1(n_641), .B2(n_663), .Y(n_639) );
CKINVDCx20_ASAP7_75t_R g640 ( .A(n_68), .Y(n_640) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_70), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_72), .A2(n_179), .B1(n_443), .B2(n_562), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_74), .A2(n_153), .B1(n_321), .B2(n_448), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_75), .A2(n_96), .B1(n_414), .B2(n_468), .Y(n_467) );
AO22x1_ASAP7_75t_L g456 ( .A1(n_76), .A2(n_457), .B1(n_458), .B2(n_484), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_76), .Y(n_484) );
AOI22xp33_ASAP7_75t_SL g583 ( .A1(n_77), .A2(n_146), .B1(n_493), .B2(n_584), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_78), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_79), .A2(n_252), .B1(n_341), .B2(n_476), .Y(n_617) );
AOI22xp33_ASAP7_75t_SL g842 ( .A1(n_80), .A2(n_154), .B1(n_448), .B2(n_471), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_82), .A2(n_172), .B1(n_407), .B2(n_769), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_83), .A2(n_141), .B1(n_421), .B2(n_445), .Y(n_444) );
AOI22xp33_ASAP7_75t_SL g648 ( .A1(n_84), .A2(n_218), .B1(n_649), .B2(n_651), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_87), .A2(n_200), .B1(n_562), .B2(n_565), .Y(n_561) );
AOI22xp33_ASAP7_75t_SL g591 ( .A1(n_88), .A2(n_207), .B1(n_417), .B2(n_538), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_89), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g679 ( .A(n_90), .Y(n_679) );
AND2x2_ASAP7_75t_L g277 ( .A(n_92), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_93), .B(n_499), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_94), .A2(n_131), .B1(n_724), .B2(n_810), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_95), .Y(n_614) );
AOI22xp33_ASAP7_75t_SL g596 ( .A1(n_97), .A2(n_180), .B1(n_540), .B2(n_597), .Y(n_596) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_98), .Y(n_799) );
INVx1_ASAP7_75t_L g274 ( .A(n_99), .Y(n_274) );
INVx1_ASAP7_75t_L g576 ( .A(n_100), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_101), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_102), .A2(n_176), .B1(n_517), .B2(n_765), .Y(n_764) );
AOI22xp33_ASAP7_75t_SL g836 ( .A1(n_103), .A2(n_224), .B1(n_362), .B2(n_504), .Y(n_836) );
AOI22xp33_ASAP7_75t_SL g624 ( .A1(n_105), .A2(n_256), .B1(n_597), .B2(n_625), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_106), .A2(n_229), .B1(n_421), .B2(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_107), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_108), .A2(n_188), .B1(n_508), .B2(n_509), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_109), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_110), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_112), .B(n_395), .Y(n_394) );
AOI222xp33_ASAP7_75t_L g482 ( .A1(n_113), .A2(n_140), .B1(n_258), .B2(n_360), .C1(n_366), .C2(n_483), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g688 ( .A(n_114), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_115), .A2(n_163), .B1(n_362), .B2(n_367), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_116), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_119), .A2(n_123), .B1(n_362), .B2(n_529), .Y(n_528) );
AOI22xp33_ASAP7_75t_SL g654 ( .A1(n_120), .A2(n_213), .B1(n_655), .B2(n_656), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_121), .A2(n_286), .B1(n_370), .B2(n_371), .Y(n_285) );
INVx1_ASAP7_75t_L g370 ( .A(n_121), .Y(n_370) );
INVx1_ASAP7_75t_L g353 ( .A(n_122), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_124), .A2(n_262), .B1(n_538), .B2(n_540), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_125), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_126), .B(n_476), .Y(n_835) );
AOI22xp33_ASAP7_75t_SL g620 ( .A1(n_127), .A2(n_246), .B1(n_472), .B2(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g331 ( .A(n_128), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_129), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_130), .A2(n_166), .B1(n_521), .B2(n_720), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_132), .A2(n_170), .B1(n_627), .B2(n_813), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_133), .A2(n_164), .B1(n_471), .B2(n_472), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_134), .A2(n_245), .B1(n_503), .B2(n_504), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_135), .A2(n_193), .B1(n_512), .B2(n_514), .Y(n_511) );
AOI222xp33_ASAP7_75t_L g738 ( .A1(n_136), .A2(n_171), .B1(n_206), .B2(n_361), .C1(n_366), .C2(n_483), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_137), .Y(n_805) );
INVx1_ASAP7_75t_L g310 ( .A(n_138), .Y(n_310) );
INVx2_ASAP7_75t_L g278 ( .A(n_144), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_145), .A2(n_236), .B1(n_493), .B2(n_494), .Y(n_492) );
AO22x1_ASAP7_75t_L g665 ( .A1(n_147), .A2(n_666), .B1(n_698), .B2(n_699), .Y(n_665) );
INVx1_ASAP7_75t_L g698 ( .A(n_147), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_148), .A2(n_269), .B1(n_483), .B2(n_646), .Y(n_645) );
AOI22xp33_ASAP7_75t_SL g662 ( .A1(n_149), .A2(n_155), .B1(n_406), .B2(n_512), .Y(n_662) );
CKINVDCx20_ASAP7_75t_R g672 ( .A(n_150), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_151), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_152), .A2(n_159), .B1(n_520), .B2(n_521), .Y(n_843) );
INVx1_ASAP7_75t_L g335 ( .A(n_156), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_157), .A2(n_241), .B1(n_584), .B2(n_649), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_158), .A2(n_214), .B1(n_409), .B2(n_517), .Y(n_516) );
AOI22xp33_ASAP7_75t_SL g657 ( .A1(n_160), .A2(n_263), .B1(n_472), .B2(n_658), .Y(n_657) );
AND2x6_ASAP7_75t_L g273 ( .A(n_161), .B(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_161), .Y(n_783) );
AO22x2_ASAP7_75t_L g293 ( .A1(n_162), .A2(n_223), .B1(n_294), .B2(n_295), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_165), .A2(n_220), .B1(n_475), .B2(n_476), .Y(n_474) );
INVx1_ASAP7_75t_L g598 ( .A(n_167), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_168), .A2(n_222), .B1(n_450), .B2(n_451), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_173), .A2(n_261), .B1(n_463), .B2(n_465), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_175), .A2(n_230), .B1(n_538), .B2(n_655), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_181), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_182), .A2(n_211), .B1(n_413), .B2(n_461), .Y(n_460) );
AOI22xp33_ASAP7_75t_SL g592 ( .A1(n_183), .A2(n_216), .B1(n_305), .B2(n_593), .Y(n_592) );
INVxp67_ASAP7_75t_L g825 ( .A(n_184), .Y(n_825) );
XNOR2x1_ASAP7_75t_L g827 ( .A(n_184), .B(n_828), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_185), .B(n_527), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_186), .B(n_366), .Y(n_677) );
AO22x2_ASAP7_75t_L g298 ( .A1(n_187), .A2(n_238), .B1(n_294), .B2(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_189), .B(n_568), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_190), .Y(n_397) );
XOR2x2_ASAP7_75t_L g725 ( .A(n_191), .B(n_726), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g792 ( .A1(n_192), .A2(n_793), .B1(n_815), .B2(n_816), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_192), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_195), .A2(n_740), .B1(n_771), .B2(n_772), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_195), .Y(n_771) );
INVx1_ASAP7_75t_L g695 ( .A(n_196), .Y(n_695) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_197), .Y(n_398) );
INVx1_ASAP7_75t_L g439 ( .A(n_198), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_199), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g674 ( .A(n_203), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_204), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_205), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_208), .B(n_526), .Y(n_834) );
AOI22xp33_ASAP7_75t_SL g588 ( .A1(n_209), .A2(n_264), .B1(n_479), .B2(n_483), .Y(n_588) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_210), .Y(n_757) );
AOI22xp33_ASAP7_75t_SL g723 ( .A1(n_212), .A2(n_260), .B1(n_328), .B2(n_724), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_219), .A2(n_233), .B1(n_478), .B2(n_481), .Y(n_477) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_221), .A2(n_271), .B(n_279), .C(n_791), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_223), .B(n_788), .Y(n_787) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_226), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_227), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_231), .A2(n_242), .B1(n_409), .B2(n_737), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_232), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_235), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g644 ( .A(n_237), .Y(n_644) );
INVx1_ASAP7_75t_L g786 ( .A(n_238), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g687 ( .A(n_239), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_240), .A2(n_265), .B1(n_568), .B2(n_732), .Y(n_731) );
OA22x2_ASAP7_75t_L g603 ( .A1(n_243), .A2(n_604), .B1(n_605), .B2(n_630), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g604 ( .A(n_243), .Y(n_604) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_248), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g612 ( .A(n_250), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_251), .B(n_475), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g380 ( .A(n_253), .Y(n_380) );
INVx1_ASAP7_75t_L g294 ( .A(n_254), .Y(n_294) );
INVx1_ASAP7_75t_L g296 ( .A(n_254), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_259), .B(n_493), .Y(n_801) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_266), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_267), .Y(n_430) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_274), .Y(n_782) );
OAI21xp5_ASAP7_75t_L g823 ( .A1(n_275), .A2(n_781), .B(n_824), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_276), .Y(n_275) );
INVxp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_637), .B1(n_776), .B2(n_777), .C(n_778), .Y(n_279) );
INVx1_ASAP7_75t_L g776 ( .A(n_280), .Y(n_776) );
AOI22xp5_ASAP7_75t_SL g280 ( .A1(n_281), .A2(n_547), .B1(n_548), .B2(n_636), .Y(n_280) );
INVx1_ASAP7_75t_L g636 ( .A(n_281), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B1(n_372), .B2(n_546), .Y(n_281) );
CKINVDCx14_ASAP7_75t_R g282 ( .A(n_283), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g371 ( .A(n_286), .Y(n_371) );
AND4x1_ASAP7_75t_L g286 ( .A(n_287), .B(n_320), .C(n_340), .D(n_359), .Y(n_286) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx3_ASAP7_75t_L g413 ( .A(n_289), .Y(n_413) );
BUFx3_ASAP7_75t_L g627 ( .A(n_289), .Y(n_627) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
BUFx2_ASAP7_75t_SL g443 ( .A(n_290), .Y(n_443) );
INVx2_ASAP7_75t_L g513 ( .A(n_290), .Y(n_513) );
BUFx2_ASAP7_75t_SL g718 ( .A(n_290), .Y(n_718) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_300), .Y(n_290) );
AND2x6_ASAP7_75t_L g323 ( .A(n_291), .B(n_324), .Y(n_323) );
AND2x4_ASAP7_75t_L g329 ( .A(n_291), .B(n_313), .Y(n_329) );
AND2x6_ASAP7_75t_L g361 ( .A(n_291), .B(n_356), .Y(n_361) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_297), .Y(n_291) );
AND2x2_ASAP7_75t_L g308 ( .A(n_292), .B(n_298), .Y(n_308) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g314 ( .A(n_293), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_293), .B(n_298), .Y(n_319) );
AND2x2_ASAP7_75t_L g351 ( .A(n_293), .B(n_302), .Y(n_351) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g299 ( .A(n_296), .Y(n_299) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g315 ( .A(n_298), .Y(n_315) );
INVx1_ASAP7_75t_L g365 ( .A(n_298), .Y(n_365) );
AND2x4_ASAP7_75t_L g307 ( .A(n_300), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_300), .B(n_314), .Y(n_334) );
AND2x4_ASAP7_75t_L g338 ( .A(n_300), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g405 ( .A(n_300), .B(n_314), .Y(n_405) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
AND2x2_ASAP7_75t_L g313 ( .A(n_301), .B(n_304), .Y(n_313) );
OR2x2_ASAP7_75t_L g325 ( .A(n_301), .B(n_304), .Y(n_325) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g356 ( .A(n_302), .B(n_304), .Y(n_356) );
INVx1_ASAP7_75t_L g352 ( .A(n_303), .Y(n_352) );
AND2x2_ASAP7_75t_L g364 ( .A(n_303), .B(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g318 ( .A(n_304), .Y(n_318) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx3_ASAP7_75t_L g414 ( .A(n_307), .Y(n_414) );
BUFx3_ASAP7_75t_L g450 ( .A(n_307), .Y(n_450) );
BUFx3_ASAP7_75t_L g520 ( .A(n_307), .Y(n_520) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_307), .Y(n_564) );
AND2x4_ASAP7_75t_L g343 ( .A(n_308), .B(n_324), .Y(n_343) );
AND2x6_ASAP7_75t_L g346 ( .A(n_308), .B(n_313), .Y(n_346) );
INVx1_ASAP7_75t_L g383 ( .A(n_308), .Y(n_383) );
NAND2x1p5_ASAP7_75t_L g387 ( .A(n_308), .B(n_313), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_311), .B1(n_316), .B2(n_317), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_311), .A2(n_687), .B1(n_688), .B2(n_689), .Y(n_686) );
BUFx2_ASAP7_75t_R g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_313), .B(n_314), .Y(n_312) );
AND2x2_ASAP7_75t_L g419 ( .A(n_313), .B(n_314), .Y(n_419) );
INVx1_ASAP7_75t_L g358 ( .A(n_315), .Y(n_358) );
INVx6_ASAP7_75t_SL g421 ( .A(n_317), .Y(n_421) );
INVx1_ASAP7_75t_SL g765 ( .A(n_317), .Y(n_765) );
OR2x6_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g480 ( .A(n_318), .Y(n_480) );
INVx1_ASAP7_75t_L g339 ( .A(n_319), .Y(n_339) );
INVx4_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_322), .Y(n_469) );
INVx2_ASAP7_75t_SL g508 ( .A(n_322), .Y(n_508) );
INVx2_ASAP7_75t_L g560 ( .A(n_322), .Y(n_560) );
INVx1_ASAP7_75t_L g737 ( .A(n_322), .Y(n_737) );
INVx11_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx11_ASAP7_75t_L g539 ( .A(n_323), .Y(n_539) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g382 ( .A(n_325), .B(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx6_ASAP7_75t_L g410 ( .A(n_329), .Y(n_410) );
BUFx3_ASAP7_75t_L g540 ( .A(n_329), .Y(n_540) );
BUFx3_ASAP7_75t_L g655 ( .A(n_329), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_332), .B1(n_335), .B2(n_336), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
BUFx2_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
BUFx3_ASAP7_75t_L g407 ( .A(n_338), .Y(n_407) );
BUFx2_ASAP7_75t_L g451 ( .A(n_338), .Y(n_451) );
BUFx3_ASAP7_75t_L g465 ( .A(n_338), .Y(n_465) );
BUFx3_ASAP7_75t_L g514 ( .A(n_338), .Y(n_514) );
INVx1_ASAP7_75t_L g535 ( .A(n_338), .Y(n_535) );
BUFx2_ASAP7_75t_SL g565 ( .A(n_338), .Y(n_565) );
BUFx3_ASAP7_75t_L g597 ( .A(n_338), .Y(n_597) );
AND2x2_ASAP7_75t_L g593 ( .A(n_339), .B(n_352), .Y(n_593) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx5_ASAP7_75t_L g475 ( .A(n_342), .Y(n_475) );
INVx2_ASAP7_75t_L g526 ( .A(n_342), .Y(n_526) );
INVx4_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_SL g568 ( .A(n_345), .Y(n_568) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
BUFx2_ASAP7_75t_L g476 ( .A(n_346), .Y(n_476) );
BUFx2_ASAP7_75t_L g501 ( .A(n_346), .Y(n_501) );
BUFx4f_ASAP7_75t_L g527 ( .A(n_346), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_349), .B1(n_353), .B2(n_354), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_349), .A2(n_354), .B1(n_438), .B2(n_439), .Y(n_437) );
BUFx3_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_350), .A2(n_397), .B1(n_398), .B2(n_399), .Y(n_396) );
INVx4_ASAP7_75t_L g681 ( .A(n_350), .Y(n_681) );
NAND2x1p5_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
AND2x4_ASAP7_75t_L g363 ( .A(n_351), .B(n_364), .Y(n_363) );
AND2x4_ASAP7_75t_L g368 ( .A(n_351), .B(n_369), .Y(n_368) );
AND2x4_ASAP7_75t_L g479 ( .A(n_351), .B(n_480), .Y(n_479) );
BUFx2_ASAP7_75t_L g399 ( .A(n_354), .Y(n_399) );
CKINVDCx16_ASAP7_75t_R g684 ( .A(n_354), .Y(n_684) );
OR2x6_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x4_ASAP7_75t_L g481 ( .A(n_356), .B(n_358), .Y(n_481) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_SL g389 ( .A(n_360), .Y(n_389) );
INVx2_ASAP7_75t_L g751 ( .A(n_360), .Y(n_751) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx3_ASAP7_75t_L g435 ( .A(n_361), .Y(n_435) );
INVx2_ASAP7_75t_SL g490 ( .A(n_361), .Y(n_490) );
INVx4_ASAP7_75t_L g572 ( .A(n_361), .Y(n_572) );
INVx2_ASAP7_75t_L g581 ( .A(n_361), .Y(n_581) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_362), .Y(n_392) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx4f_ASAP7_75t_SL g483 ( .A(n_363), .Y(n_483) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_363), .Y(n_503) );
BUFx2_ASAP7_75t_L g575 ( .A(n_363), .Y(n_575) );
INVx1_ASAP7_75t_L g369 ( .A(n_365), .Y(n_369) );
BUFx4f_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g544 ( .A(n_367), .Y(n_544) );
BUFx12f_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_368), .Y(n_395) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_368), .Y(n_493) );
INVx1_ASAP7_75t_L g546 ( .A(n_372), .Y(n_546) );
XNOR2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_454), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B1(n_424), .B2(n_453), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g423 ( .A(n_377), .Y(n_423) );
AND2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_400), .Y(n_377) );
NOR3xp33_ASAP7_75t_L g378 ( .A(n_379), .B(n_388), .C(n_396), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_381), .B1(n_384), .B2(n_385), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_381), .A2(n_743), .B1(n_744), .B2(n_745), .Y(n_742) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_381), .A2(n_385), .B1(n_796), .B2(n_797), .Y(n_795) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx3_ASAP7_75t_L g429 ( .A(n_382), .Y(n_429) );
INVx2_ASAP7_75t_L g671 ( .A(n_382), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_385), .A2(n_669), .B1(n_670), .B2(n_672), .Y(n_668) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g431 ( .A(n_386), .Y(n_431) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx3_ASAP7_75t_L g747 ( .A(n_387), .Y(n_747) );
OAI221xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_390), .B1(n_391), .B2(n_393), .C(n_394), .Y(n_388) );
OAI21xp5_ASAP7_75t_SL g709 ( .A1(n_389), .A2(n_710), .B(n_711), .Y(n_709) );
INVx2_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_SL g675 ( .A(n_392), .Y(n_675) );
INVx1_ASAP7_75t_L g613 ( .A(n_395), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_399), .A2(n_803), .B1(n_804), .B2(n_805), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_401), .B(n_411), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_408), .Y(n_401) );
BUFx3_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx3_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx3_ASAP7_75t_L g463 ( .A(n_405), .Y(n_463) );
BUFx3_ASAP7_75t_L g510 ( .A(n_405), .Y(n_510) );
BUFx3_ASAP7_75t_L g532 ( .A(n_405), .Y(n_532) );
BUFx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx3_ASAP7_75t_L g448 ( .A(n_410), .Y(n_448) );
INVx2_ASAP7_75t_L g697 ( .A(n_410), .Y(n_697) );
INVx2_ASAP7_75t_L g810 ( .A(n_410), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_412), .B(n_415), .Y(n_411) );
INVx1_ASAP7_75t_L g629 ( .A(n_414), .Y(n_629) );
BUFx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx6f_ASAP7_75t_L g720 ( .A(n_417), .Y(n_720) );
INVx5_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g445 ( .A(n_418), .Y(n_445) );
INVx3_ASAP7_75t_L g471 ( .A(n_418), .Y(n_471) );
BUFx3_ASAP7_75t_L g518 ( .A(n_418), .Y(n_518) );
INVx4_ASAP7_75t_L g557 ( .A(n_418), .Y(n_557) );
INVx1_ASAP7_75t_L g622 ( .A(n_418), .Y(n_622) );
INVx8_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx2_ASAP7_75t_L g472 ( .A(n_421), .Y(n_472) );
BUFx2_ASAP7_75t_L g521 ( .A(n_421), .Y(n_521) );
BUFx4f_ASAP7_75t_SL g690 ( .A(n_421), .Y(n_690) );
INVx2_ASAP7_75t_SL g453 ( .A(n_424), .Y(n_453) );
XOR2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_452), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_440), .Y(n_425) );
NOR3xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_432), .C(n_437), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_429), .B1(n_430), .B2(n_431), .Y(n_427) );
OAI21xp33_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B(n_436), .Y(n_432) );
OAI21xp5_ASAP7_75t_SL g643 ( .A1(n_434), .A2(n_644), .B(n_645), .Y(n_643) );
OAI221xp5_ASAP7_75t_L g673 ( .A1(n_434), .A2(n_674), .B1(n_675), .B2(n_676), .C(n_677), .Y(n_673) );
INVx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_441), .B(n_446), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_444), .Y(n_441) );
INVx1_ASAP7_75t_L g761 ( .A(n_443), .Y(n_761) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_445), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_447), .B(n_449), .Y(n_446) );
BUFx2_ASAP7_75t_L g656 ( .A(n_450), .Y(n_656) );
XNOR2x1_ASAP7_75t_L g454 ( .A(n_455), .B(n_485), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
NAND4xp75_ASAP7_75t_SL g458 ( .A(n_459), .B(n_466), .C(n_473), .D(n_482), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_464), .Y(n_459) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_470), .Y(n_466) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_SL g473 ( .A(n_474), .B(n_477), .Y(n_473) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_475), .Y(n_499) );
BUFx6f_ASAP7_75t_L g732 ( .A(n_475), .Y(n_732) );
BUFx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g504 ( .A(n_479), .Y(n_504) );
BUFx3_ASAP7_75t_L g529 ( .A(n_479), .Y(n_529) );
INVx1_ASAP7_75t_L g650 ( .A(n_479), .Y(n_650) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_481), .Y(n_496) );
BUFx2_ASAP7_75t_SL g545 ( .A(n_481), .Y(n_545) );
BUFx2_ASAP7_75t_SL g584 ( .A(n_481), .Y(n_584) );
BUFx3_ASAP7_75t_L g651 ( .A(n_481), .Y(n_651) );
INVx1_ASAP7_75t_L g611 ( .A(n_483), .Y(n_611) );
INVx1_ASAP7_75t_L g749 ( .A(n_483), .Y(n_749) );
XOR2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_522), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_488), .B(n_505), .Y(n_487) );
NOR2xp33_ASAP7_75t_SL g488 ( .A(n_489), .B(n_497), .Y(n_488) );
OAI21xp5_ASAP7_75t_SL g489 ( .A1(n_490), .A2(n_491), .B(n_492), .Y(n_489) );
BUFx2_ASAP7_75t_L g646 ( .A(n_493), .Y(n_646) );
INVx2_ASAP7_75t_L g753 ( .A(n_493), .Y(n_753) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
NAND3xp33_ASAP7_75t_L g497 ( .A(n_498), .B(n_500), .C(n_502), .Y(n_497) );
NOR2x1_ASAP7_75t_L g505 ( .A(n_506), .B(n_515), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_511), .Y(n_506) );
BUFx4f_ASAP7_75t_SL g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g770 ( .A(n_510), .Y(n_770) );
INVx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_519), .Y(n_515) );
INVx3_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_520), .Y(n_813) );
NAND4xp75_ASAP7_75t_L g523 ( .A(n_524), .B(n_530), .C(n_536), .D(n_542), .Y(n_523) );
AND2x2_ASAP7_75t_SL g524 ( .A(n_525), .B(n_528), .Y(n_524) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_533), .Y(n_530) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_541), .Y(n_536) );
INVx4_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx3_ASAP7_75t_L g625 ( .A(n_539), .Y(n_625) );
INVx4_ASAP7_75t_L g661 ( .A(n_539), .Y(n_661) );
INVx2_ASAP7_75t_SL g724 ( .A(n_539), .Y(n_724) );
INVx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OAI22xp5_ASAP7_75t_SL g548 ( .A1(n_549), .A2(n_550), .B1(n_601), .B2(n_602), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_577), .B1(n_599), .B2(n_600), .Y(n_550) );
INVx2_ASAP7_75t_SL g599 ( .A(n_551), .Y(n_599) );
XOR2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_576), .Y(n_551) );
NOR4xp75_ASAP7_75t_L g552 ( .A(n_553), .B(n_558), .C(n_566), .D(n_570), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_554), .B(n_555), .Y(n_553) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2x1_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
INVx4_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OAI221xp5_ASAP7_75t_SL g760 ( .A1(n_563), .A2(n_761), .B1(n_762), .B2(n_763), .C(n_764), .Y(n_760) );
INVx4_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_567), .B(n_569), .Y(n_566) );
OAI21xp5_ASAP7_75t_SL g570 ( .A1(n_571), .A2(n_573), .B(n_574), .Y(n_570) );
OAI221xp5_ASAP7_75t_SL g798 ( .A1(n_571), .A2(n_611), .B1(n_799), .B2(n_800), .C(n_801), .Y(n_798) );
BUFx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx4_ASAP7_75t_L g609 ( .A(n_572), .Y(n_609) );
OAI21xp5_ASAP7_75t_SL g830 ( .A1(n_572), .A2(n_831), .B(n_832), .Y(n_830) );
INVx1_ASAP7_75t_L g600 ( .A(n_577), .Y(n_600) );
INVx2_ASAP7_75t_L g632 ( .A(n_577), .Y(n_632) );
XOR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_598), .Y(n_577) );
NAND2x1_ASAP7_75t_L g578 ( .A(n_579), .B(n_589), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_580), .B(n_585), .Y(n_579) );
OAI21xp5_ASAP7_75t_SL g580 ( .A1(n_581), .A2(n_582), .B(n_583), .Y(n_580) );
NAND3xp33_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .C(n_588), .Y(n_585) );
NOR2x1_ASAP7_75t_L g589 ( .A(n_590), .B(n_594), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
INVx1_ASAP7_75t_L g635 ( .A(n_600), .Y(n_635) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_631), .B1(n_633), .B2(n_634), .Y(n_602) );
INVx1_ASAP7_75t_L g633 ( .A(n_603), .Y(n_633) );
INVx2_ASAP7_75t_L g630 ( .A(n_605), .Y(n_630) );
NAND3x1_ASAP7_75t_L g605 ( .A(n_606), .B(n_618), .C(n_623), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_615), .Y(n_606) );
OAI222xp33_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_610), .B1(n_611), .B2(n_612), .C1(n_613), .C2(n_614), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g777 ( .A(n_637), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_701), .B1(n_774), .B2(n_775), .Y(n_637) );
INVx1_ASAP7_75t_L g774 ( .A(n_638), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_664), .B1(n_665), .B2(n_700), .Y(n_638) );
INVx1_ASAP7_75t_L g700 ( .A(n_639), .Y(n_700) );
INVx1_ASAP7_75t_SL g663 ( .A(n_641), .Y(n_663) );
NAND3x1_ASAP7_75t_L g641 ( .A(n_642), .B(n_653), .C(n_659), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_647), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_652), .Y(n_647) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_657), .Y(n_653) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_662), .Y(n_659) );
INVx1_ASAP7_75t_L g694 ( .A(n_661), .Y(n_694) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g699 ( .A(n_666), .Y(n_699) );
AND3x1_ASAP7_75t_L g666 ( .A(n_667), .B(n_685), .C(n_691), .Y(n_666) );
NOR3xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_673), .C(n_678), .Y(n_667) );
INVx1_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_680), .B1(n_682), .B2(n_683), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_680), .A2(n_756), .B1(n_757), .B2(n_758), .Y(n_755) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx3_ASAP7_75t_SL g804 ( .A(n_681), .Y(n_804) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g758 ( .A(n_684), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_690), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_694), .B1(n_695), .B2(n_696), .Y(n_692) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g775 ( .A(n_701), .Y(n_775) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_705), .B1(n_739), .B2(n_773), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
XNOR2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_725), .Y(n_705) );
NAND3xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_716), .C(n_721), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_709), .B(n_712), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .C(n_715), .Y(n_712) );
AND2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_719), .Y(n_716) );
AND2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
NAND4xp75_ASAP7_75t_L g726 ( .A(n_727), .B(n_730), .C(n_734), .D(n_738), .Y(n_726) );
AND2x2_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
AND2x2_ASAP7_75t_SL g730 ( .A(n_731), .B(n_733), .Y(n_730) );
AND2x2_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
INVx1_ASAP7_75t_L g773 ( .A(n_739), .Y(n_773) );
INVx1_ASAP7_75t_L g772 ( .A(n_740), .Y(n_772) );
AND2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_759), .Y(n_740) );
NOR3xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_748), .C(n_755), .Y(n_741) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OAI222xp33_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_750), .B1(n_751), .B2(n_752), .C1(n_753), .C2(n_754), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_766), .Y(n_759) );
NAND2xp5_ASAP7_75t_SL g766 ( .A(n_767), .B(n_768), .Y(n_766) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_SL g778 ( .A(n_779), .Y(n_778) );
NOR2x1_ASAP7_75t_L g779 ( .A(n_780), .B(n_784), .Y(n_779) );
OR2x2_ASAP7_75t_SL g846 ( .A(n_780), .B(n_785), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_781), .B(n_783), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_782), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_782), .B(n_821), .Y(n_824) );
CKINVDCx16_ASAP7_75t_R g821 ( .A(n_783), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_785), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_787), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_789), .B(n_790), .Y(n_788) );
OAI322xp33_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_817), .A3(n_818), .B1(n_822), .B2(n_825), .C1(n_826), .C2(n_844), .Y(n_791) );
INVx2_ASAP7_75t_L g816 ( .A(n_793), .Y(n_816) );
AND2x2_ASAP7_75t_SL g793 ( .A(n_794), .B(n_806), .Y(n_793) );
NOR3xp33_ASAP7_75t_L g794 ( .A(n_795), .B(n_798), .C(n_802), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_807), .B(n_811), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_812), .B(n_814), .Y(n_811) );
HB1xp67_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
HB1xp67_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
CKINVDCx20_ASAP7_75t_R g822 ( .A(n_823), .Y(n_822) );
INVx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
AND2x4_ASAP7_75t_L g828 ( .A(n_829), .B(n_837), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_830), .B(n_833), .Y(n_829) );
NAND3xp33_ASAP7_75t_L g833 ( .A(n_834), .B(n_835), .C(n_836), .Y(n_833) );
NOR2x1_ASAP7_75t_L g837 ( .A(n_838), .B(n_841), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_839), .B(n_840), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_842), .B(n_843), .Y(n_841) );
CKINVDCx20_ASAP7_75t_R g844 ( .A(n_845), .Y(n_844) );
CKINVDCx20_ASAP7_75t_R g845 ( .A(n_846), .Y(n_845) );
endmodule