module real_jpeg_2896_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_247;
wire n_146;
wire n_78;
wire n_249;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_205;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_244;
wire n_213;
wire n_128;
wire n_179;
wire n_216;
wire n_133;
wire n_202;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_48),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_45),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_45),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_3),
.A2(n_45),
.B1(n_57),
.B2(n_59),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_4),
.A2(n_39),
.B1(n_57),
.B2(n_59),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_4),
.A2(n_39),
.B1(n_67),
.B2(n_68),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_4),
.B(n_57),
.C(n_72),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_4),
.B(n_75),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_4),
.B(n_25),
.C(n_54),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_4),
.B(n_43),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_4),
.B(n_29),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_4),
.B(n_30),
.C(n_32),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_4),
.B(n_52),
.Y(n_213)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_23)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_6),
.A2(n_27),
.B1(n_57),
.B2(n_59),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_6),
.A2(n_27),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_6),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_138)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_236),
.B1(n_257),
.B2(n_258),
.Y(n_13)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_14),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_126),
.B(n_235),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_104),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_17),
.B(n_104),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_80),
.C(n_91),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_18),
.B(n_80),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_49),
.B2(n_50),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_19),
.B(n_51),
.C(n_79),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_40),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_21),
.A2(n_22),
.B1(n_40),
.B2(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_21),
.A2(n_22),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_21),
.A2(n_22),
.B1(n_186),
.B2(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_22),
.B(n_181),
.C(n_186),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_22),
.B(n_137),
.C(n_213),
.Y(n_218)
);

OA22x2_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_37),
.B2(n_38),
.Y(n_22)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_23),
.A2(n_28),
.B1(n_37),
.B2(n_38),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_25),
.B1(n_30),
.B2(n_35),
.Y(n_36)
);

AOI22x1_ASAP7_75t_L g53 ( 
.A1(n_24),
.A2(n_25),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_25),
.B(n_206),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_28),
.A2(n_37),
.B(n_38),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_28),
.B(n_37),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_36),
.Y(n_28)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_29),
.A2(n_89),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

AO22x1_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_29)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_32),
.B(n_199),
.Y(n_198)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_37),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_40),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_41),
.B(n_46),
.Y(n_83)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_42),
.B(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_42),
.A2(n_43),
.B1(n_96),
.B2(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_44),
.A2(n_46),
.B(n_95),
.Y(n_94)
);

OA21x2_ASAP7_75t_L g157 ( 
.A1(n_46),
.A2(n_95),
.B(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_47),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_64),
.B1(n_78),
.B2(n_79),
.Y(n_50)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_51),
.B(n_100),
.C(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_51),
.A2(n_78),
.B1(n_148),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_51),
.A2(n_78),
.B1(n_97),
.B2(n_98),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_51),
.B(n_97),
.C(n_221),
.Y(n_227)
);

AO21x1_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_56),
.B(n_60),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_52),
.A2(n_56),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_53),
.A2(n_61),
.B(n_62),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_53),
.A2(n_249),
.B(n_251),
.Y(n_248)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_59),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_57),
.Y(n_59)
);

AO22x1_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_59),
.B1(n_72),
.B2(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_57),
.B(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_60),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_64),
.A2(n_79),
.B1(n_121),
.B2(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_64),
.B(n_121),
.C(n_132),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_71),
.B1(n_75),
.B2(n_77),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OA21x2_ASAP7_75t_L g101 ( 
.A1(n_66),
.A2(n_102),
.B(n_103),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_67),
.A2(n_72),
.B(n_74),
.C(n_75),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_72),
.Y(n_74)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_68),
.B(n_135),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_77),
.Y(n_103)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_72),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_84),
.B1(n_85),
.B2(n_90),
.Y(n_80)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_85),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_81),
.A2(n_90),
.B1(n_112),
.B2(n_115),
.Y(n_111)
);

INVxp33_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_83),
.B(n_96),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_90),
.A2(n_108),
.B(n_115),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_91),
.B(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_99),
.C(n_100),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_92),
.A2(n_93),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_94),
.A2(n_97),
.B1(n_98),
.B2(n_145),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_94),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_97),
.A2(n_98),
.B1(n_205),
.B2(n_207),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_97),
.B(n_207),
.Y(n_215)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_99),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_100),
.A2(n_101),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_100),
.A2(n_101),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_102),
.B(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_125),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_116),
.B2(n_117),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_107),
.B(n_116),
.C(n_125),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_112),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_121),
.B(n_124),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_121),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g246 ( 
.A(n_120),
.B(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_156),
.C(n_157),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_121),
.A2(n_140),
.B1(n_182),
.B2(n_185),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_124),
.A2(n_241),
.B1(n_242),
.B2(n_253),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_124),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_230),
.B(n_234),
.Y(n_126)
);

OAI211xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_159),
.B(n_173),
.C(n_174),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_149),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_149),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_141),
.B2(n_142),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_144),
.C(n_146),
.Y(n_161)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_139),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_134),
.B1(n_136),
.B2(n_137),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_136),
.A2(n_137),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_137),
.B(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_137),
.B(n_201),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_148),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_154),
.C(n_155),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_155),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_157),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NAND3xp33_ASAP7_75t_SL g174 ( 
.A(n_160),
.B(n_175),
.C(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_162),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_163),
.B(n_165),
.C(n_171),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_170),
.B2(n_171),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21x1_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_192),
.B(n_229),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_178),
.B(n_180),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_182),
.Y(n_185)
);

NOR2xp67_ASAP7_75t_SL g203 ( 
.A(n_184),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_204),
.Y(n_208)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_187),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_223),
.B(n_228),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_217),
.B(n_222),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_209),
.B(n_216),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_203),
.B(n_208),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_200),
.B(n_202),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_205),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_215),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_215),
.Y(n_216)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_213),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_219),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_227),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_231),
.B(n_232),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_236),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_255),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_238),
.B(n_239),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_254),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_248),
.B2(n_252),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_248),
.Y(n_252)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);


endmodule