module fake_jpeg_4900_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_SL g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_24),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_25),
.B(n_28),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_31),
.A2(n_32),
.B1(n_19),
.B2(n_23),
.Y(n_44)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_34),
.B(n_36),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_17),
.B(n_11),
.C(n_19),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_35),
.A2(n_39),
.B1(n_26),
.B2(n_2),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_11),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g38 ( 
.A1(n_24),
.A2(n_15),
.B(n_16),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_17),
.B1(n_26),
.B2(n_24),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_15),
.B1(n_16),
.B2(n_13),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_22),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_42),
.B(n_14),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_47),
.B(n_55),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_11),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_53),
.Y(n_64)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_19),
.B(n_21),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_56),
.B(n_61),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_21),
.B1(n_20),
.B2(n_23),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_14),
.Y(n_53)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_1),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_59),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_45),
.B(n_1),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_60),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_46),
.B(n_43),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_72),
.Y(n_76)
);

AND2x6_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_46),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_69),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_47),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_79),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_56),
.C(n_55),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_67),
.C(n_70),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_52),
.B1(n_61),
.B2(n_53),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_77),
.A2(n_62),
.B1(n_65),
.B2(n_71),
.Y(n_82)
);

INVxp33_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_52),
.Y(n_79)
);

NOR3xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_4),
.C(n_5),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_80),
.B(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

AOI221xp5_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_76),
.B1(n_78),
.B2(n_40),
.C(n_9),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_62),
.B(n_70),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_75),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_76),
.C(n_41),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_83),
.B(n_41),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_89),
.A2(n_87),
.B(n_84),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_86),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_91),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_85),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_41),
.C(n_40),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_93),
.A2(n_96),
.B(n_92),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_94),
.B(n_88),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_95),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_4),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_98),
.A2(n_99),
.B(n_6),
.Y(n_101)
);

BUFx24_ASAP7_75t_SL g102 ( 
.A(n_100),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_101),
.C(n_7),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_10),
.Y(n_104)
);


endmodule