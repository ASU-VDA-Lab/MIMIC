module fake_netlist_6_124_n_489 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_489);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_489;

wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_209;
wire n_367;
wire n_465;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_148;
wire n_208;
wire n_161;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_350;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_372;
wire n_468;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_375;
wire n_338;
wire n_466;
wire n_360;
wire n_235;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_428;
wire n_432;
wire n_167;
wire n_174;
wire n_153;
wire n_156;
wire n_145;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_294;
wire n_302;
wire n_380;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_397;
wire n_155;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_172;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_460;
wire n_417;
wire n_446;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_456;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_455;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_152;
wire n_321;
wire n_331;
wire n_227;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_476;
wire n_291;
wire n_219;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_477;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_282;
wire n_436;
wire n_211;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_273;
wire n_311;
wire n_403;
wire n_253;
wire n_136;
wire n_249;
wire n_201;
wire n_386;
wire n_159;
wire n_157;
wire n_162;
wire n_487;
wire n_241;
wire n_275;
wire n_276;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_277;
wire n_418;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_453;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_347;
wire n_459;
wire n_328;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_205;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_288;
wire n_427;
wire n_479;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_187;
wire n_361;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

INVx1_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_2),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_40),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_97),
.Y(n_143)
);

INVxp67_ASAP7_75t_SL g144 ( 
.A(n_86),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_52),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_68),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_15),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_71),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_3),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

INVxp33_ASAP7_75t_SL g153 ( 
.A(n_122),
.Y(n_153)
);

INVxp67_ASAP7_75t_SL g154 ( 
.A(n_118),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_0),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_70),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_14),
.B(n_111),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_3),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_38),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_74),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

INVxp33_ASAP7_75t_SL g163 ( 
.A(n_121),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_69),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_96),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_81),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_95),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_83),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_92),
.Y(n_169)
);

INVx4_ASAP7_75t_R g170 ( 
.A(n_105),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_31),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_45),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_55),
.Y(n_173)
);

INVxp67_ASAP7_75t_SL g174 ( 
.A(n_98),
.Y(n_174)
);

BUFx2_ASAP7_75t_SL g175 ( 
.A(n_6),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_125),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_16),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_59),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_51),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_47),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_35),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_120),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_43),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_21),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_27),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_54),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_24),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_63),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_44),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_110),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_101),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_78),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_61),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_89),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_4),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_130),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_106),
.Y(n_198)
);

INVxp33_ASAP7_75t_SL g199 ( 
.A(n_126),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_32),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_84),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_133),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_5),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_6),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_2),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_64),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_119),
.Y(n_207)
);

INVxp67_ASAP7_75t_SL g208 ( 
.A(n_22),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_143),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_202),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_151),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_155),
.Y(n_213)
);

OA21x2_ASAP7_75t_L g214 ( 
.A1(n_159),
.A2(n_203),
.B(n_196),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_171),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_182),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_183),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_139),
.B(n_0),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_R g222 ( 
.A(n_160),
.B(n_1),
.Y(n_222)
);

INVxp33_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_145),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_134),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_206),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_135),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_137),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_147),
.B(n_1),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_165),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_180),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_138),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_177),
.B(n_4),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_150),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_207),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_185),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_139),
.B(n_5),
.Y(n_238)
);

INVxp67_ASAP7_75t_SL g239 ( 
.A(n_188),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_140),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_188),
.B(n_7),
.Y(n_241)
);

AND2x4_ASAP7_75t_L g242 ( 
.A(n_152),
.B(n_10),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_174),
.Y(n_243)
);

BUFx2_ASAP7_75t_SL g244 ( 
.A(n_187),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_141),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_153),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_163),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_199),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_211),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_174),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_226),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_234),
.A2(n_208),
.B1(n_204),
.B2(n_136),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_229),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_190),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_229),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_231),
.Y(n_259)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_190),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_235),
.Y(n_263)
);

AO22x2_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_208),
.B1(n_200),
.B2(n_201),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_235),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_245),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_233),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_221),
.B(n_192),
.Y(n_268)
);

AND2x4_ASAP7_75t_L g269 ( 
.A(n_232),
.B(n_144),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_192),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_232),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_214),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_214),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_214),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_210),
.Y(n_275)
);

AND2x4_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_154),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_209),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_212),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_221),
.B(n_244),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_210),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_222),
.B(n_142),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_217),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_225),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_212),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_215),
.B(n_146),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_217),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_259),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_216),
.Y(n_289)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_263),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_267),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_248),
.B(n_220),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_248),
.A2(n_246),
.B1(n_237),
.B2(n_236),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_227),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_250),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_260),
.B(n_224),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_260),
.B(n_224),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_283),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_275),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_278),
.Y(n_300)
);

NAND3xp33_ASAP7_75t_L g301 ( 
.A(n_268),
.B(n_213),
.C(n_223),
.Y(n_301)
);

AND2x4_ASAP7_75t_L g302 ( 
.A(n_269),
.B(n_276),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_260),
.B(n_218),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_273),
.A2(n_218),
.B(n_219),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_280),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_256),
.A2(n_222),
.B1(n_223),
.B2(n_219),
.Y(n_306)
);

AO22x1_ASAP7_75t_L g307 ( 
.A1(n_247),
.A2(n_198),
.B1(n_197),
.B2(n_195),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_277),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_277),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_263),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_282),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_261),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_260),
.B(n_148),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_249),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_278),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_286),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_278),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_285),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_265),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_263),
.Y(n_320)
);

INVx5_ASAP7_75t_L g321 ( 
.A(n_284),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_276),
.B(n_149),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_269),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_252),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_251),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_247),
.Y(n_326)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_284),
.Y(n_327)
);

NAND3xp33_ASAP7_75t_SL g328 ( 
.A(n_254),
.B(n_194),
.C(n_193),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_270),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g330 ( 
.A(n_281),
.B(n_156),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_291),
.Y(n_331)
);

BUFx4f_ASAP7_75t_SL g332 ( 
.A(n_298),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_324),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_272),
.Y(n_334)
);

AND2x4_ASAP7_75t_L g335 ( 
.A(n_300),
.B(n_251),
.Y(n_335)
);

INVx3_ASAP7_75t_SL g336 ( 
.A(n_308),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_296),
.A2(n_274),
.B(n_256),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_302),
.B(n_262),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_302),
.B(n_262),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_295),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_289),
.B(n_264),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_287),
.Y(n_342)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_323),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_297),
.A2(n_264),
.B(n_266),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_312),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_270),
.Y(n_346)
);

OR2x6_ASAP7_75t_L g347 ( 
.A(n_288),
.B(n_264),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_319),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_323),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_326),
.B(n_157),
.Y(n_350)
);

AND2x6_ASAP7_75t_L g351 ( 
.A(n_314),
.B(n_161),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_294),
.B(n_162),
.Y(n_352)
);

NOR2x1_ASAP7_75t_SL g353 ( 
.A(n_322),
.B(n_164),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_318),
.Y(n_354)
);

AO22x2_ASAP7_75t_L g355 ( 
.A1(n_328),
.A2(n_178),
.B1(n_166),
.B2(n_167),
.Y(n_355)
);

NAND2x1p5_ASAP7_75t_L g356 ( 
.A(n_315),
.B(n_253),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_301),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_299),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_306),
.B(n_255),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_317),
.Y(n_360)
);

OR2x6_ASAP7_75t_L g361 ( 
.A(n_307),
.B(n_293),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_292),
.B(n_168),
.Y(n_362)
);

A2O1A1Ixp33_ASAP7_75t_L g363 ( 
.A1(n_330),
.A2(n_158),
.B(n_179),
.C(n_191),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_330),
.Y(n_364)
);

OR2x6_ASAP7_75t_L g365 ( 
.A(n_309),
.B(n_169),
.Y(n_365)
);

OAI321xp33_ASAP7_75t_L g366 ( 
.A1(n_313),
.A2(n_181),
.A3(n_172),
.B1(n_189),
.B2(n_186),
.C(n_184),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_310),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_311),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_334),
.B(n_304),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_299),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_354),
.B(n_321),
.Y(n_371)
);

OAI21x1_ASAP7_75t_L g372 ( 
.A1(n_337),
.A2(n_303),
.B(n_320),
.Y(n_372)
);

OAI22xp33_ASAP7_75t_L g373 ( 
.A1(n_361),
.A2(n_327),
.B1(n_321),
.B2(n_316),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_342),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_359),
.B(n_305),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_361),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_335),
.B(n_327),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_335),
.B(n_327),
.Y(n_378)
);

CKINVDCx11_ASAP7_75t_R g379 ( 
.A(n_336),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g380 ( 
.A1(n_352),
.A2(n_316),
.B1(n_305),
.B2(n_173),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_338),
.A2(n_339),
.B(n_343),
.Y(n_381)
);

NAND2x1p5_ASAP7_75t_L g382 ( 
.A(n_343),
.B(n_290),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_358),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_332),
.Y(n_384)
);

OAI21x1_ASAP7_75t_L g385 ( 
.A1(n_344),
.A2(n_258),
.B(n_257),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_341),
.A2(n_176),
.B1(n_310),
.B2(n_290),
.Y(n_386)
);

O2A1O1Ixp33_ASAP7_75t_L g387 ( 
.A1(n_357),
.A2(n_170),
.B(n_8),
.C(n_9),
.Y(n_387)
);

AO31x2_ASAP7_75t_L g388 ( 
.A1(n_363),
.A2(n_7),
.A3(n_8),
.B(n_9),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_364),
.A2(n_331),
.B(n_368),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_349),
.A2(n_310),
.B(n_12),
.Y(n_390)
);

INVx6_ASAP7_75t_L g391 ( 
.A(n_360),
.Y(n_391)
);

AOI221xp5_ASAP7_75t_L g392 ( 
.A1(n_350),
.A2(n_11),
.B1(n_13),
.B2(n_17),
.C(n_18),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_333),
.B(n_19),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_347),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_340),
.Y(n_395)
);

AOI21xp33_ASAP7_75t_L g396 ( 
.A1(n_355),
.A2(n_20),
.B(n_23),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_345),
.Y(n_397)
);

OAI221xp5_ASAP7_75t_L g398 ( 
.A1(n_362),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.C(n_29),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_L g399 ( 
.A1(n_355),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_383),
.Y(n_400)
);

OA21x2_ASAP7_75t_L g401 ( 
.A1(n_385),
.A2(n_366),
.B(n_348),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_374),
.Y(n_402)
);

AOI21x1_ASAP7_75t_L g403 ( 
.A1(n_381),
.A2(n_353),
.B(n_365),
.Y(n_403)
);

OAI21x1_ASAP7_75t_L g404 ( 
.A1(n_372),
.A2(n_367),
.B(n_356),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_375),
.B(n_353),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_375),
.B(n_351),
.Y(n_406)
);

AOI221xp5_ASAP7_75t_L g407 ( 
.A1(n_387),
.A2(n_351),
.B1(n_365),
.B2(n_39),
.C(n_41),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_395),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_371),
.B(n_36),
.Y(n_409)
);

OAI221xp5_ASAP7_75t_L g410 ( 
.A1(n_394),
.A2(n_37),
.B1(n_42),
.B2(n_46),
.C(n_48),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_384),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_L g412 ( 
.A1(n_396),
.A2(n_399),
.B1(n_392),
.B2(n_398),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_370),
.B(n_49),
.Y(n_413)
);

OAI22xp33_ASAP7_75t_L g414 ( 
.A1(n_376),
.A2(n_132),
.B1(n_53),
.B2(n_56),
.Y(n_414)
);

OAI21x1_ASAP7_75t_L g415 ( 
.A1(n_369),
.A2(n_50),
.B(n_57),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_391),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_369),
.A2(n_60),
.B(n_62),
.Y(n_417)
);

AOI221xp5_ASAP7_75t_L g418 ( 
.A1(n_396),
.A2(n_65),
.B1(n_72),
.B2(n_73),
.C(n_76),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_397),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_L g420 ( 
.A1(n_370),
.A2(n_79),
.B1(n_82),
.B2(n_85),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_408),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_406),
.B(n_377),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_378),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_405),
.B(n_393),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_412),
.A2(n_407),
.B1(n_405),
.B2(n_413),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_418),
.A2(n_382),
.B(n_386),
.Y(n_426)
);

OAI221xp5_ASAP7_75t_L g427 ( 
.A1(n_412),
.A2(n_389),
.B1(n_384),
.B2(n_380),
.C(n_386),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_L g428 ( 
.A1(n_400),
.A2(n_393),
.B1(n_373),
.B2(n_391),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_408),
.Y(n_429)
);

AOI211xp5_ASAP7_75t_L g430 ( 
.A1(n_414),
.A2(n_390),
.B(n_379),
.C(n_388),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_419),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_403),
.Y(n_432)
);

AO21x2_ASAP7_75t_L g433 ( 
.A1(n_404),
.A2(n_388),
.B(n_382),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_411),
.B(n_131),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_409),
.Y(n_435)
);

OAI221xp5_ASAP7_75t_L g436 ( 
.A1(n_420),
.A2(n_87),
.B1(n_90),
.B2(n_91),
.C(n_93),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_421),
.Y(n_437)
);

OR2x2_ASAP7_75t_L g438 ( 
.A(n_422),
.B(n_402),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_422),
.B(n_416),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_423),
.B(n_420),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_431),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_433),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_423),
.B(n_415),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_429),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_435),
.B(n_424),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_434),
.B(n_415),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_432),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_428),
.B(n_404),
.Y(n_448)
);

NAND2x1_ASAP7_75t_L g449 ( 
.A(n_426),
.B(n_417),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g450 ( 
.A(n_427),
.B(n_401),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_425),
.B(n_401),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_433),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_445),
.B(n_430),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_439),
.B(n_433),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_441),
.B(n_426),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g456 ( 
.A(n_438),
.B(n_401),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_440),
.B(n_410),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_441),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_443),
.B(n_94),
.Y(n_459)
);

INVx3_ASAP7_75t_SL g460 ( 
.A(n_446),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_437),
.B(n_444),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_448),
.B(n_436),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_447),
.Y(n_463)
);

NAND2xp33_ASAP7_75t_R g464 ( 
.A(n_448),
.B(n_99),
.Y(n_464)
);

NAND4xp75_ASAP7_75t_L g465 ( 
.A(n_451),
.B(n_100),
.C(n_102),
.D(n_103),
.Y(n_465)
);

NOR2x1_ASAP7_75t_L g466 ( 
.A(n_465),
.B(n_455),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_453),
.A2(n_449),
.B1(n_450),
.B2(n_448),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_463),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_458),
.B(n_454),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_460),
.B(n_104),
.Y(n_470)
);

AOI221x1_ASAP7_75t_L g471 ( 
.A1(n_463),
.A2(n_452),
.B1(n_442),
.B2(n_107),
.C(n_108),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_452),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_469),
.B(n_456),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_468),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_472),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_466),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_474),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_475),
.B(n_467),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_476),
.A2(n_471),
.B(n_470),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_R g480 ( 
.A(n_478),
.B(n_464),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_477),
.B(n_473),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_479),
.A2(n_462),
.B1(n_459),
.B2(n_457),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_482),
.A2(n_481),
.B(n_480),
.Y(n_483)
);

CKINVDCx12_ASAP7_75t_R g484 ( 
.A(n_483),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_484),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_485),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_486),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_SL g488 ( 
.A1(n_487),
.A2(n_114),
.B1(n_115),
.B2(n_123),
.Y(n_488)
);

AOI221xp5_ASAP7_75t_L g489 ( 
.A1(n_488),
.A2(n_487),
.B1(n_124),
.B2(n_127),
.C(n_128),
.Y(n_489)
);


endmodule