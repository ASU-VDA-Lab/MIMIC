module fake_jpeg_2321_n_495 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_495);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_495;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_479;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVxp33_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_56),
.Y(n_146)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g178 ( 
.A(n_57),
.Y(n_178)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_58),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_59),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_64),
.Y(n_139)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_23),
.B(n_17),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_68),
.B(n_73),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_23),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_69),
.B(n_93),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_71),
.Y(n_149)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_72),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_0),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_32),
.B(n_0),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_106),
.Y(n_123)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_75),
.Y(n_169)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_76),
.Y(n_154)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_78),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_79),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_80),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_20),
.B(n_0),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_82),
.B(n_112),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_84),
.Y(n_189)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_86),
.Y(n_191)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g161 ( 
.A(n_87),
.Y(n_161)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_88),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_89),
.Y(n_168)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_90),
.Y(n_183)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_91),
.Y(n_194)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_92),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_54),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_96),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_98),
.Y(n_193)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_99),
.B(n_105),
.Y(n_141)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_102),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_103),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_104),
.Y(n_127)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_24),
.Y(n_106)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_24),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_107),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_20),
.B(n_0),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_114),
.Y(n_147)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_35),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_113),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_29),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_110),
.Y(n_173)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_111),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_37),
.B(n_1),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_42),
.Y(n_113)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_42),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_36),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_116),
.Y(n_143)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_36),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g117 ( 
.A(n_51),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_47),
.Y(n_151)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_50),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_53),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_28),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g195 ( 
.A1(n_119),
.A2(n_5),
.B(n_8),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_83),
.A2(n_34),
.B1(n_47),
.B2(n_44),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_121),
.A2(n_136),
.B1(n_138),
.B2(n_145),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_74),
.A2(n_25),
.B1(n_45),
.B2(n_43),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_89),
.A2(n_34),
.B1(n_47),
.B2(n_44),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_73),
.A2(n_25),
.B1(n_45),
.B2(n_43),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_151),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_68),
.B(n_37),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_153),
.B(n_164),
.Y(n_201)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_101),
.B(n_34),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_156),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_82),
.A2(n_42),
.B1(n_19),
.B2(n_41),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_159),
.A2(n_172),
.B1(n_177),
.B2(n_179),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_112),
.A2(n_31),
.B1(n_21),
.B2(n_41),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_162),
.A2(n_166),
.B1(n_87),
.B2(n_77),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_85),
.B(n_30),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_53),
.C(n_50),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_165),
.B(n_167),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_103),
.A2(n_30),
.B1(n_39),
.B2(n_21),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_60),
.B(n_39),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_SL g237 ( 
.A(n_171),
.B(n_189),
.C(n_139),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_100),
.A2(n_38),
.B1(n_22),
.B2(n_27),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_63),
.A2(n_31),
.B1(n_27),
.B2(n_19),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_114),
.A2(n_22),
.B1(n_38),
.B2(n_97),
.Y(n_179)
);

CKINVDCx12_ASAP7_75t_R g181 ( 
.A(n_67),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_102),
.A2(n_38),
.B1(n_22),
.B2(n_3),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_182),
.A2(n_184),
.B1(n_185),
.B2(n_188),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_104),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_70),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_110),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_113),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_192),
.A2(n_146),
.B1(n_168),
.B2(n_194),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_195),
.A2(n_91),
.B(n_96),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_111),
.B(n_14),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_10),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_143),
.A2(n_95),
.B1(n_79),
.B2(n_71),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_198),
.A2(n_202),
.B1(n_230),
.B2(n_243),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_199),
.Y(n_264)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_140),
.Y(n_203)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_203),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_205),
.B(n_214),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_141),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_206),
.B(n_223),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_207),
.B(n_237),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_147),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_208),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_L g209 ( 
.A1(n_179),
.A2(n_172),
.B1(n_138),
.B2(n_121),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_209),
.A2(n_211),
.B1(n_218),
.B2(n_204),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_123),
.B(n_11),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_210),
.B(n_216),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_133),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_150),
.Y(n_212)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_212),
.Y(n_304)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_213),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_152),
.B(n_14),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_152),
.B(n_133),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_215),
.B(n_255),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_165),
.B(n_156),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_184),
.A2(n_188),
.B1(n_192),
.B2(n_175),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_156),
.B(n_126),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_221),
.B(n_227),
.Y(n_271)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_154),
.Y(n_222)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_222),
.Y(n_283)
);

A2O1A1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_141),
.A2(n_144),
.B(n_130),
.C(n_128),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_132),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_224),
.B(n_253),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_190),
.A2(n_186),
.B1(n_160),
.B2(n_173),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_226),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_124),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_127),
.B(n_176),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_228),
.B(n_234),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_190),
.A2(n_186),
.B(n_182),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_229),
.A2(n_209),
.B(n_249),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_142),
.A2(n_169),
.B1(n_154),
.B2(n_149),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_142),
.Y(n_231)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_231),
.Y(n_275)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_169),
.Y(n_232)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_232),
.Y(n_277)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_122),
.Y(n_233)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_233),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_187),
.B(n_160),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_132),
.Y(n_235)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_235),
.Y(n_281)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_150),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_236),
.Y(n_303)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_122),
.Y(n_238)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_238),
.Y(n_287)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_120),
.Y(n_239)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_239),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_180),
.B(n_139),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_240),
.B(n_245),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_125),
.B(n_174),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_241),
.B(n_251),
.Y(n_289)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_125),
.Y(n_242)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_242),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_194),
.A2(n_196),
.B1(n_155),
.B2(n_149),
.Y(n_243)
);

INVx11_ASAP7_75t_L g244 ( 
.A(n_170),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_244),
.A2(n_256),
.B1(n_200),
.B2(n_199),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_180),
.B(n_157),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_129),
.A2(n_146),
.B1(n_157),
.B2(n_189),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_246),
.B(n_248),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_134),
.A2(n_137),
.B1(n_155),
.B2(n_135),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_247),
.A2(n_252),
.B1(n_243),
.B2(n_246),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_131),
.B(n_183),
.Y(n_248)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_120),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_250),
.B(n_254),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_174),
.B(n_129),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_134),
.A2(n_135),
.B1(n_137),
.B2(n_178),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_163),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_131),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_178),
.B(n_163),
.Y(n_255)
);

AND2x2_ASAP7_75t_SL g257 ( 
.A(n_191),
.B(n_196),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_200),
.C(n_248),
.Y(n_268)
);

A2O1A1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_148),
.A2(n_123),
.B(n_153),
.C(n_152),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_221),
.Y(n_279)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_191),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_260),
.Y(n_293)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_168),
.Y(n_260)
);

FAx1_ASAP7_75t_SL g261 ( 
.A(n_148),
.B(n_123),
.CI(n_152),
.CON(n_261),
.SN(n_261)
);

AOI32xp33_ASAP7_75t_L g306 ( 
.A1(n_261),
.A2(n_258),
.A3(n_211),
.B1(n_234),
.B2(n_251),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_142),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_262),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_263),
.A2(n_290),
.B1(n_291),
.B2(n_266),
.Y(n_322)
);

OR2x2_ASAP7_75t_SL g328 ( 
.A(n_268),
.B(n_279),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_203),
.A2(n_216),
.B1(n_220),
.B2(n_207),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_272),
.A2(n_284),
.B1(n_308),
.B2(n_310),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_276),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_280),
.A2(n_267),
.B(n_309),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_202),
.A2(n_206),
.B1(n_229),
.B2(n_261),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_282),
.A2(n_267),
.B1(n_269),
.B2(n_306),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_220),
.A2(n_225),
.B1(n_210),
.B2(n_218),
.Y(n_284)
);

OA22x2_ASAP7_75t_L g295 ( 
.A1(n_223),
.A2(n_217),
.B1(n_257),
.B2(n_261),
.Y(n_295)
);

AO22x2_ASAP7_75t_L g348 ( 
.A1(n_295),
.A2(n_296),
.B1(n_294),
.B2(n_275),
.Y(n_348)
);

OA22x2_ASAP7_75t_L g296 ( 
.A1(n_217),
.A2(n_257),
.B1(n_235),
.B2(n_220),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_227),
.B(n_228),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_311),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_254),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_301),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_201),
.B(n_213),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_307),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_231),
.B(n_232),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_241),
.A2(n_222),
.B1(n_242),
.B2(n_233),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_238),
.A2(n_253),
.B1(n_245),
.B2(n_240),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_240),
.B(n_245),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_280),
.A2(n_212),
.B1(n_236),
.B2(n_244),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_312),
.A2(n_321),
.B1(n_322),
.B2(n_294),
.Y(n_349)
);

AO22x1_ASAP7_75t_SL g313 ( 
.A1(n_284),
.A2(n_248),
.B1(n_259),
.B2(n_250),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_313),
.B(n_336),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_272),
.B(n_260),
.C(n_239),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_316),
.B(n_329),
.C(n_332),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_300),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_317),
.B(n_323),
.Y(n_359)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_273),
.Y(n_318)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_318),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_270),
.B(n_219),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_319),
.B(n_324),
.C(n_328),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_290),
.A2(n_219),
.B1(n_289),
.B2(n_270),
.Y(n_321)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_292),
.Y(n_323)
);

MAJx2_ASAP7_75t_L g324 ( 
.A(n_279),
.B(n_271),
.C(n_292),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_325),
.A2(n_337),
.B(n_340),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_265),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_326),
.B(n_330),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_297),
.B(n_278),
.Y(n_327)
);

NAND3xp33_ASAP7_75t_L g368 ( 
.A(n_327),
.B(n_305),
.C(n_331),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_265),
.B(n_271),
.C(n_296),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_286),
.B(n_299),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_278),
.C(n_268),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_273),
.Y(n_333)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_333),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_293),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_334),
.B(n_335),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_303),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_289),
.B(n_296),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_266),
.A2(n_267),
.B1(n_309),
.B2(n_291),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_281),
.Y(n_338)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_338),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_304),
.Y(n_339)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_339),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_295),
.B(n_281),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_341),
.B(n_347),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_295),
.B(n_294),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_342),
.B(n_348),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_264),
.B(n_288),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_343),
.B(n_345),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_274),
.A2(n_309),
.B1(n_295),
.B2(n_310),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_344),
.A2(n_275),
.B1(n_277),
.B2(n_287),
.Y(n_350)
);

INVx8_ASAP7_75t_L g345 ( 
.A(n_303),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_311),
.B(n_288),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_349),
.A2(n_350),
.B1(n_362),
.B2(n_365),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_314),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_352),
.B(n_356),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_347),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_341),
.A2(n_285),
.B(n_277),
.Y(n_358)
);

XNOR2x1_ASAP7_75t_L g383 ( 
.A(n_358),
.B(n_360),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_342),
.A2(n_298),
.B(n_264),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_346),
.A2(n_298),
.B1(n_304),
.B2(n_302),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_346),
.A2(n_287),
.B1(n_302),
.B2(n_283),
.Y(n_365)
);

OAI21xp33_ASAP7_75t_L g367 ( 
.A1(n_320),
.A2(n_305),
.B(n_283),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_367),
.B(n_368),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_332),
.B(n_328),
.C(n_329),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_369),
.B(n_337),
.C(n_313),
.Y(n_386)
);

O2A1O1Ixp33_ASAP7_75t_L g371 ( 
.A1(n_336),
.A2(n_348),
.B(n_340),
.C(n_312),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_371),
.B(n_375),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_321),
.A2(n_315),
.B1(n_344),
.B2(n_331),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_374),
.A2(n_377),
.B1(n_348),
.B2(n_318),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_327),
.B(n_315),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_376),
.B(n_319),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_325),
.A2(n_316),
.B1(n_317),
.B2(n_313),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_334),
.B(n_313),
.Y(n_378)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_378),
.Y(n_380)
);

XOR2x2_ASAP7_75t_L g381 ( 
.A(n_376),
.B(n_324),
.Y(n_381)
);

XNOR2x1_ASAP7_75t_L g408 ( 
.A(n_381),
.B(n_364),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_361),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_382),
.B(n_388),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_384),
.B(n_386),
.C(n_390),
.Y(n_409)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_372),
.Y(n_385)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_385),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_361),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_372),
.Y(n_389)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_389),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_369),
.B(n_348),
.C(n_335),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_370),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_391),
.B(n_399),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_369),
.B(n_348),
.C(n_333),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_392),
.B(n_400),
.C(n_351),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_393),
.A2(n_396),
.B1(n_402),
.B2(n_353),
.Y(n_410)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_354),
.Y(n_394)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_394),
.Y(n_424)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_354),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_395),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_377),
.A2(n_338),
.B1(n_339),
.B2(n_345),
.Y(n_396)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_373),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_364),
.B(n_339),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_373),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_401),
.B(n_403),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_350),
.A2(n_349),
.B1(n_378),
.B2(n_374),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_370),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_402),
.A2(n_380),
.B1(n_398),
.B2(n_393),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_404),
.A2(n_410),
.B1(n_419),
.B2(n_398),
.Y(n_436)
);

INVx4_ASAP7_75t_L g406 ( 
.A(n_391),
.Y(n_406)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_406),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_408),
.B(n_381),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_400),
.B(n_364),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_411),
.B(n_412),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_384),
.B(n_355),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_385),
.Y(n_413)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_413),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_403),
.B(n_360),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_417),
.A2(n_383),
.B(n_388),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_380),
.A2(n_375),
.B1(n_353),
.B2(n_356),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_379),
.B(n_368),
.Y(n_420)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_420),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_379),
.B(n_363),
.Y(n_421)
);

NAND3xp33_ASAP7_75t_L g432 ( 
.A(n_421),
.B(n_425),
.C(n_359),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_392),
.B(n_358),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_422),
.B(n_351),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_423),
.B(n_390),
.C(n_386),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_382),
.B(n_363),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_426),
.A2(n_417),
.B(n_418),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_428),
.B(n_435),
.C(n_440),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_407),
.A2(n_397),
.B(n_352),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_429),
.B(n_432),
.Y(n_449)
);

BUFx24_ASAP7_75t_SL g431 ( 
.A(n_414),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_431),
.B(n_441),
.Y(n_446)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_414),
.Y(n_433)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_433),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_434),
.B(n_439),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_411),
.B(n_383),
.C(n_355),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_436),
.A2(n_404),
.B1(n_387),
.B2(n_406),
.Y(n_443)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_418),
.Y(n_438)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_438),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_409),
.B(n_396),
.C(n_366),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_409),
.B(n_366),
.C(n_387),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_443),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_441),
.B(n_359),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_447),
.B(n_452),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_442),
.B(n_423),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_450),
.B(n_442),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_437),
.B(n_416),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_451),
.Y(n_463)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_437),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_436),
.B(n_416),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_454),
.B(n_417),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_455),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_457),
.B(n_450),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_453),
.B(n_440),
.C(n_428),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_460),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_451),
.Y(n_460)
);

INVxp33_ASAP7_75t_L g461 ( 
.A(n_449),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_461),
.B(n_466),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_449),
.A2(n_430),
.B1(n_420),
.B2(n_426),
.Y(n_462)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_462),
.B(n_464),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_446),
.B(n_427),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_467),
.B(n_468),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_456),
.A2(n_445),
.B1(n_448),
.B2(n_454),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_458),
.B(n_453),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_469),
.B(n_472),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_463),
.B(n_445),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_465),
.A2(n_455),
.B(n_435),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_473),
.B(n_471),
.C(n_470),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_448),
.Y(n_475)
);

MAJx2_ASAP7_75t_L g479 ( 
.A(n_475),
.B(n_459),
.C(n_460),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_474),
.B(n_457),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_478),
.B(n_480),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_479),
.B(n_481),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_471),
.B(n_475),
.C(n_456),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_472),
.B(n_424),
.Y(n_482)
);

AOI21xp33_ASAP7_75t_L g484 ( 
.A1(n_482),
.A2(n_399),
.B(n_401),
.Y(n_484)
);

NAND4xp25_ASAP7_75t_L g483 ( 
.A(n_477),
.B(n_452),
.C(n_415),
.D(n_405),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_483),
.A2(n_413),
.B(n_357),
.Y(n_490)
);

OAI321xp33_ASAP7_75t_L g488 ( 
.A1(n_484),
.A2(n_485),
.A3(n_395),
.B1(n_394),
.B2(n_389),
.C(n_486),
.Y(n_488)
);

AO21x1_ASAP7_75t_L g487 ( 
.A1(n_479),
.A2(n_439),
.B(n_422),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_487),
.B(n_434),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_488),
.A2(n_489),
.B(n_476),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_490),
.B(n_443),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_491),
.B(n_492),
.C(n_408),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_493),
.A2(n_444),
.B1(n_412),
.B2(n_371),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_494),
.B(n_444),
.Y(n_495)
);


endmodule