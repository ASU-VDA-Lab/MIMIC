module fake_jpeg_23764_n_242 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_242);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_242;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_4),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_30),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_61),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_29),
.B1(n_35),
.B2(n_21),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_51),
.A2(n_68),
.B(n_34),
.Y(n_82)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_32),
.B(n_18),
.C(n_22),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_58),
.B(n_72),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_29),
.B1(n_35),
.B2(n_22),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_27),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_16),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_16),
.Y(n_67)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

NAND2xp33_ASAP7_75t_SL g68 ( 
.A(n_43),
.B(n_27),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_42),
.B(n_30),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_75),
.Y(n_93)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_36),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_40),
.B(n_25),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_79),
.B(n_31),
.Y(n_107)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_84),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_82),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_51),
.A2(n_33),
.B(n_17),
.C(n_25),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_83),
.A2(n_71),
.B1(n_56),
.B2(n_49),
.Y(n_126)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_44),
.C(n_40),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_92),
.Y(n_117)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_23),
.Y(n_88)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_74),
.B(n_24),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_90),
.B(n_91),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_52),
.Y(n_91)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_4),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_27),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_104),
.Y(n_113)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_59),
.Y(n_128)
);

AO22x1_ASAP7_75t_SL g101 ( 
.A1(n_49),
.A2(n_44),
.B1(n_37),
.B2(n_2),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_101),
.A2(n_71),
.B1(n_70),
.B2(n_37),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_23),
.Y(n_102)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

OAI32xp33_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_19),
.A3(n_31),
.B1(n_34),
.B2(n_24),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_70),
.B(n_17),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_106),
.B(n_107),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_53),
.B(n_19),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_108),
.B(n_48),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_76),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_111),
.B(n_6),
.Y(n_157)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_122),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_132),
.B1(n_134),
.B2(n_104),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_119),
.B(n_120),
.Y(n_158)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_127),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_96),
.B1(n_98),
.B2(n_93),
.Y(n_141)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_80),
.B(n_59),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_129),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_59),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_133),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_136),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_89),
.B(n_107),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_89),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_145),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_92),
.Y(n_140)
);

XOR2x2_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_113),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_148),
.B1(n_153),
.B2(n_122),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_146),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_97),
.Y(n_145)
);

BUFx4f_ASAP7_75t_SL g146 ( 
.A(n_114),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_127),
.A2(n_97),
.B1(n_93),
.B2(n_109),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_109),
.B(n_94),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_149),
.A2(n_116),
.B(n_112),
.Y(n_181)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_151),
.B(n_156),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_95),
.B1(n_103),
.B2(n_84),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_113),
.A2(n_94),
.B1(n_95),
.B2(n_103),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_154),
.A2(n_110),
.B(n_112),
.Y(n_180)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_157),
.B(n_160),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_115),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_123),
.Y(n_178)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_133),
.B(n_123),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_161),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_111),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_172),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_144),
.C(n_116),
.Y(n_197)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_166),
.B(n_169),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_167),
.A2(n_156),
.B1(n_160),
.B2(n_139),
.Y(n_188)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_120),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_110),
.Y(n_173)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_175),
.Y(n_184)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_100),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_180),
.B(n_181),
.Y(n_196)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_178),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_155),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_187),
.Y(n_203)
);

A2O1A1O1Ixp25_ASAP7_75t_L g183 ( 
.A1(n_171),
.A2(n_150),
.B(n_149),
.C(n_157),
.D(n_161),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_197),
.C(n_144),
.Y(n_202)
);

NAND2x1_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_148),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_186),
.A2(n_189),
.B(n_177),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_142),
.Y(n_187)
);

AOI221xp5_ASAP7_75t_L g201 ( 
.A1(n_188),
.A2(n_192),
.B1(n_170),
.B2(n_167),
.C(n_164),
.Y(n_201)
);

OA21x2_ASAP7_75t_L g189 ( 
.A1(n_163),
.A2(n_141),
.B(n_146),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_168),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_190),
.Y(n_204)
);

AOI21xp33_ASAP7_75t_L g192 ( 
.A1(n_172),
.A2(n_159),
.B(n_151),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_169),
.A2(n_139),
.B1(n_152),
.B2(n_158),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_195),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_209)
);

BUFx12f_ASAP7_75t_SL g198 ( 
.A(n_186),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_198),
.A2(n_189),
.B1(n_196),
.B2(n_183),
.Y(n_217)
);

AOI322xp5_ASAP7_75t_L g199 ( 
.A1(n_196),
.A2(n_176),
.A3(n_164),
.B1(n_180),
.B2(n_179),
.C1(n_166),
.C2(n_174),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_202),
.C(n_208),
.Y(n_218)
);

NOR3xp33_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_181),
.C(n_175),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_200),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_201),
.Y(n_214)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_185),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_206),
.Y(n_213)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_207),
.A2(n_189),
.B1(n_195),
.B2(n_194),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_62),
.C(n_13),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_209),
.A2(n_197),
.B1(n_187),
.B2(n_10),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_184),
.B(n_11),
.Y(n_210)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_210),
.Y(n_215)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_207),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_212),
.A2(n_217),
.B(n_220),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_202),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_220),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_198),
.A2(n_182),
.B1(n_11),
.B2(n_10),
.Y(n_220)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_213),
.C(n_206),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_226),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_211),
.B(n_204),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_223),
.B(n_225),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_215),
.B(n_205),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_203),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_203),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_231),
.A2(n_232),
.B(n_214),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_213),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_233),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_229),
.A2(n_221),
.B1(n_222),
.B2(n_219),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_235),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_228),
.A2(n_218),
.B(n_208),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_230),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_232),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_9),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_241),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_238),
.A2(n_10),
.B(n_237),
.Y(n_241)
);


endmodule