module fake_jpeg_16361_n_92 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_92);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_92;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_11),
.B(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_7),
.B(n_2),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_0),
.B(n_5),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_12),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_24),
.B(n_31),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_16),
.A2(n_10),
.B1(n_9),
.B2(n_2),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_25),
.A2(n_26),
.B1(n_29),
.B2(n_6),
.Y(n_42)
);

OAI32xp33_ASAP7_75t_L g26 ( 
.A1(n_12),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_27),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_16),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_15),
.A2(n_5),
.B(n_6),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_14),
.C(n_13),
.Y(n_49)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_31),
.Y(n_34)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_23),
.A2(n_16),
.B1(n_20),
.B2(n_21),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_35),
.A2(n_37),
.B1(n_41),
.B2(n_10),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_21),
.B1(n_20),
.B2(n_19),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_15),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_40),
.C(n_46),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_17),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_19),
.B1(n_18),
.B2(n_14),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_47),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_22),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_18),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_19),
.B(n_7),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_13),
.B(n_18),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_33),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_50),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_13),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_49),
.C(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_61),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_34),
.A2(n_7),
.B(n_9),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_59),
.A2(n_63),
.B(n_39),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_45),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_42),
.B1(n_35),
.B2(n_46),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_39),
.B(n_48),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_54),
.B(n_52),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_53),
.C(n_51),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_56),
.A2(n_35),
.B1(n_37),
.B2(n_47),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_70),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_43),
.B1(n_44),
.B2(n_50),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_43),
.B1(n_44),
.B2(n_36),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_59),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_63),
.B(n_61),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_74),
.A2(n_79),
.B(n_72),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_70),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_54),
.C(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_76),
.B(n_78),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_52),
.C(n_62),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_80),
.B(n_65),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_82),
.A2(n_84),
.B(n_73),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_77),
.A2(n_67),
.B1(n_72),
.B2(n_69),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_73),
.B(n_74),
.Y(n_88)
);

AO221x1_ASAP7_75t_L g91 ( 
.A1(n_88),
.A2(n_83),
.B1(n_81),
.B2(n_65),
.C(n_55),
.Y(n_91)
);

NAND4xp25_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_86),
.C(n_90),
.D(n_89),
.Y(n_92)
);


endmodule