module fake_jpeg_15415_n_256 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_256);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

BUFx12_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_17),
.A2(n_0),
.B(n_1),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_25),
.Y(n_38)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_25),
.Y(n_40)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_22),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_48),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_21),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_14),
.B1(n_16),
.B2(n_21),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_36),
.B1(n_33),
.B2(n_14),
.Y(n_65)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_14),
.B1(n_36),
.B2(n_16),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_55),
.A2(n_65),
.B1(n_74),
.B2(n_15),
.Y(n_95)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_61),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_24),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_21),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_28),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_70),
.Y(n_86)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_56),
.Y(n_91)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_44),
.A2(n_14),
.B1(n_33),
.B2(n_22),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_17),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_75),
.B(n_19),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_28),
.B(n_34),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_76),
.A2(n_28),
.B(n_34),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_77),
.A2(n_94),
.B1(n_52),
.B2(n_47),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_71),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_85),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_30),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_34),
.C(n_29),
.Y(n_116)
);

NAND2xp33_ASAP7_75t_SL g82 ( 
.A(n_61),
.B(n_34),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_92),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_84),
.B(n_15),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_57),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_63),
.Y(n_114)
);

AO22x2_ASAP7_75t_L g94 ( 
.A1(n_58),
.A2(n_34),
.B1(n_28),
.B2(n_33),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_95),
.A2(n_46),
.B1(n_52),
.B2(n_65),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_69),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_30),
.B1(n_19),
.B2(n_17),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_97),
.A2(n_46),
.B1(n_52),
.B2(n_30),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_98),
.B(n_105),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_94),
.A2(n_77),
.B1(n_82),
.B2(n_95),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_83),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_88),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_108),
.B1(n_53),
.B2(n_39),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_103),
.A2(n_112),
.B(n_81),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_68),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_86),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_92),
.A2(n_94),
.B1(n_80),
.B2(n_76),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_94),
.A2(n_46),
.B1(n_18),
.B2(n_27),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_119),
.B1(n_113),
.B2(n_24),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_94),
.A2(n_39),
.B1(n_53),
.B2(n_47),
.Y(n_112)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_34),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_116),
.C(n_117),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_29),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_63),
.B1(n_73),
.B2(n_66),
.Y(n_119)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_135),
.B1(n_119),
.B2(n_51),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_83),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_124),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_125),
.A2(n_127),
.B(n_98),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_93),
.B(n_79),
.Y(n_127)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_133),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_99),
.A2(n_66),
.B1(n_87),
.B2(n_89),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_130),
.A2(n_140),
.B1(n_109),
.B2(n_100),
.Y(n_146)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_132),
.Y(n_158)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_35),
.C(n_31),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_137),
.C(n_90),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_101),
.A2(n_87),
.B1(n_39),
.B2(n_51),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_96),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_136),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_35),
.C(n_31),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_104),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_139),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_112),
.A2(n_103),
.B1(n_107),
.B2(n_118),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_118),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_145),
.C(n_153),
.Y(n_175)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_129),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_161),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_147),
.A2(n_152),
.B(n_159),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_102),
.C(n_110),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_148),
.B(n_139),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_141),
.A2(n_51),
.B1(n_15),
.B2(n_24),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_102),
.Y(n_153)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_123),
.A2(n_18),
.B1(n_27),
.B2(n_23),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_157),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_127),
.A2(n_54),
.B1(n_90),
.B2(n_35),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_160),
.B1(n_162),
.B2(n_132),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_125),
.A2(n_0),
.B(n_1),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_128),
.A2(n_13),
.B(n_23),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_121),
.A2(n_140),
.B(n_131),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_138),
.Y(n_162)
);

AOI21x1_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_26),
.B(n_31),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_135),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_137),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_182),
.C(n_157),
.Y(n_185)
);

MAJx2_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_120),
.C(n_128),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_167),
.A2(n_171),
.B1(n_177),
.B2(n_178),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_134),
.B1(n_131),
.B2(n_133),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_179),
.A2(n_154),
.B1(n_159),
.B2(n_156),
.Y(n_190)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_180),
.Y(n_197)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_181),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_147),
.B(n_124),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_184),
.Y(n_196)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_142),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_167),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_153),
.C(n_142),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_194),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_164),
.B1(n_151),
.B2(n_158),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_178),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_172),
.A2(n_160),
.B1(n_144),
.B2(n_155),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_144),
.C(n_90),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_26),
.C(n_13),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_198),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_26),
.C(n_13),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_165),
.A2(n_7),
.B(n_12),
.C(n_11),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_199),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_186),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_202),
.B(n_214),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_177),
.B(n_179),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_203),
.A2(n_2),
.B(n_3),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_205),
.B(n_1),
.Y(n_224)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_207),
.Y(n_215)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_192),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_182),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_210),
.C(n_204),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_197),
.A2(n_173),
.B(n_169),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_209),
.A2(n_212),
.B(n_11),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_211),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_173),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_193),
.A2(n_7),
.B(n_12),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_193),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_201),
.A2(n_200),
.B1(n_188),
.B2(n_194),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_217),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_195),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_218),
.B(n_208),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_189),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_222),
.C(n_26),
.Y(n_233)
);

OAI221xp5_ASAP7_75t_L g220 ( 
.A1(n_213),
.A2(n_191),
.B1(n_199),
.B2(n_198),
.C(n_13),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_220),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_223),
.A2(n_225),
.B1(n_212),
.B2(n_4),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_205),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_229),
.Y(n_241)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_227),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_231),
.C(n_232),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_219),
.A2(n_203),
.B1(n_4),
.B2(n_5),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_215),
.A2(n_221),
.B(n_216),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_13),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_225),
.Y(n_236)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_236),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_234),
.B(n_230),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_238),
.B(n_239),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_3),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_233),
.B(n_7),
.Y(n_240)
);

BUFx24_ASAP7_75t_SL g243 ( 
.A(n_240),
.Y(n_243)
);

OAI21x1_ASAP7_75t_L g244 ( 
.A1(n_237),
.A2(n_229),
.B(n_232),
.Y(n_244)
);

AOI21xp33_ASAP7_75t_L g249 ( 
.A1(n_244),
.A2(n_8),
.B(n_5),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_235),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_245),
.A2(n_8),
.B(n_4),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_239),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_248),
.Y(n_250)
);

A2O1A1O1Ixp25_ASAP7_75t_L g251 ( 
.A1(n_249),
.A2(n_243),
.B(n_5),
.C(n_6),
.D(n_3),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_246),
.C(n_26),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_252),
.A2(n_250),
.B(n_8),
.Y(n_253)
);

NAND3xp33_ASAP7_75t_SL g254 ( 
.A(n_253),
.B(n_3),
.C(n_5),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_254),
.A2(n_6),
.B(n_26),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_6),
.Y(n_256)
);


endmodule