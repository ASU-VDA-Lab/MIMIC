module real_jpeg_11662_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_65;
wire n_33;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g86 ( 
.A(n_2),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_3),
.A2(n_30),
.B1(n_45),
.B2(n_46),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_3),
.A2(n_30),
.B1(n_61),
.B2(n_62),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_3),
.A2(n_30),
.B1(n_37),
.B2(n_38),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_5),
.B(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_5),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_5),
.B(n_139),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_5),
.A2(n_37),
.B1(n_38),
.B2(n_103),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_5),
.B(n_62),
.C(n_86),
.Y(n_157)
);

NAND2x1_ASAP7_75t_SL g161 ( 
.A(n_5),
.B(n_36),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g183 ( 
.A1(n_5),
.A2(n_66),
.B(n_167),
.Y(n_183)
);

O2A1O1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_5),
.A2(n_27),
.B(n_35),
.C(n_194),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_103),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_6),
.A2(n_61),
.B1(n_62),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_6),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_7),
.A2(n_61),
.B1(n_62),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_7),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_9),
.A2(n_61),
.B1(n_62),
.B2(n_65),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_9),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_9),
.A2(n_37),
.B1(n_38),
.B2(n_65),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_47),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_10),
.A2(n_37),
.B1(n_38),
.B2(n_47),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_10),
.A2(n_47),
.B1(n_61),
.B2(n_62),
.Y(n_173)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_12),
.A2(n_37),
.B1(n_38),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_12),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_83),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_12),
.A2(n_61),
.B1(n_62),
.B2(n_83),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_14),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_14),
.A2(n_37),
.B1(n_38),
.B2(n_42),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_14),
.A2(n_42),
.B1(n_61),
.B2(n_62),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_15),
.A2(n_61),
.B1(n_62),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_15),
.A2(n_37),
.B1(n_38),
.B2(n_71),
.Y(n_110)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_125),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_20),
.B(n_105),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_77),
.C(n_91),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_21),
.A2(n_22),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_58),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_43),
.B2(n_57),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_24),
.B(n_57),
.C(n_58),
.Y(n_124)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B(n_40),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_26),
.A2(n_31),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_27),
.A2(n_28),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

AOI32xp33_ASAP7_75t_L g74 ( 
.A1(n_27),
.A2(n_46),
.A3(n_50),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g76 ( 
.A(n_28),
.B(n_49),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_31),
.A2(n_40),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_32),
.B(n_41),
.Y(n_122)
);

NOR2x1_ASAP7_75t_R g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

AO22x1_ASAP7_75t_SL g36 ( 
.A1(n_34),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_34),
.A2(n_37),
.B(n_103),
.Y(n_194)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g85 ( 
.A1(n_37),
.A2(n_38),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_38),
.B(n_157),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_48),
.B(n_51),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_44),
.A2(n_48),
.B1(n_53),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_54)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_46),
.A2(n_53),
.B(n_103),
.C(n_104),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_48),
.B(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_56),
.Y(n_101)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_48),
.Y(n_139)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_73),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_59),
.A2(n_73),
.B1(n_74),
.B2(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_66),
.B1(n_69),
.B2(n_72),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_60),
.A2(n_66),
.B1(n_72),
.B2(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_61),
.B(n_68),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_61),
.A2(n_62),
.B1(n_86),
.B2(n_87),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_61),
.B(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_66),
.A2(n_72),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_66),
.A2(n_166),
.B(n_167),
.Y(n_165)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_68),
.B1(n_70),
.B2(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_67),
.A2(n_68),
.B1(n_172),
.B2(n_174),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_67),
.B(n_168),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_68),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_68),
.B(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_72),
.A2(n_173),
.B(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_72),
.B(n_103),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_72),
.A2(n_141),
.B(n_181),
.Y(n_195)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_77),
.B(n_91),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_78),
.B(n_81),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_79),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B1(n_89),
.B2(n_90),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_84),
.B(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_89),
.B1(n_90),
.B2(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_84),
.A2(n_90),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_88),
.A2(n_94),
.B(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_88),
.B(n_103),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_90),
.B(n_95),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.C(n_99),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_92),
.B(n_96),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_97),
.A2(n_98),
.B(n_122),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_98),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_100),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_124),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_116),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_123),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_120),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_145),
.B(n_225),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_142),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_129),
.B(n_142),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.C(n_135),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_130),
.B(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_133),
.B(n_135),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.C(n_140),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_136),
.B(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_137),
.A2(n_138),
.B1(n_140),
.B2(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_140),
.Y(n_211)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_220),
.B(n_224),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_205),
.B(n_219),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_189),
.B(n_204),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_169),
.B(n_188),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_158),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_150),
.B(n_158),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_156),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_151),
.A2(n_152),
.B1(n_156),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B(n_155),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_154),
.A2(n_155),
.B(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_165),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_163),
.C(n_165),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_177),
.B(n_187),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_171),
.B(n_175),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_182),
.B(n_186),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_179),
.B(n_180),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_190),
.B(n_191),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_196),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_199),
.C(n_203),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_195),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_199),
.B1(n_202),
.B2(n_203),
.Y(n_196)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_199),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_206),
.B(n_207),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_212),
.B2(n_213),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_215),
.C(n_217),
.Y(n_221)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_214),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_221),
.B(n_222),
.Y(n_224)
);


endmodule