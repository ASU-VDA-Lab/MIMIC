module fake_netlist_6_3787_n_904 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_904);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_904;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_671;
wire n_607;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_893;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_222;
wire n_718;
wire n_248;
wire n_517;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_758;
wire n_516;
wire n_720;
wire n_631;
wire n_525;
wire n_842;
wire n_611;
wire n_491;
wire n_878;
wire n_772;
wire n_656;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_600;
wire n_464;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_598;
wire n_496;
wire n_422;
wire n_696;
wire n_722;
wire n_688;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_663;
wire n_508;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_678;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_122),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_100),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_167),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_38),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_142),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_64),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_80),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_16),
.Y(n_211)
);

BUFx8_ASAP7_75t_SL g212 ( 
.A(n_111),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_30),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_114),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_28),
.Y(n_215)
);

BUFx8_ASAP7_75t_SL g216 ( 
.A(n_200),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_25),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_48),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_63),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_42),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_1),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_0),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_96),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_136),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g225 ( 
.A(n_156),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_116),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_174),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_25),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_172),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_78),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_95),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_171),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_0),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_183),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_29),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_69),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_74),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_201),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_31),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_181),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_132),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_47),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_159),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_151),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_193),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_110),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_147),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_6),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_84),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_203),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_71),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_130),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_126),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_152),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_6),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_154),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_139),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_108),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_40),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_199),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_105),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_166),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_32),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_93),
.Y(n_265)
);

BUFx5_ASAP7_75t_L g266 ( 
.A(n_173),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_62),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_109),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_123),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_103),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_198),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_7),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_12),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_178),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_118),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_141),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_125),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_20),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_4),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_56),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_153),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_180),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_120),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_192),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_170),
.Y(n_285)
);

AND2x4_ASAP7_75t_L g286 ( 
.A(n_237),
.B(n_33),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_1),
.Y(n_287)
);

AND2x4_ASAP7_75t_L g288 ( 
.A(n_237),
.B(n_2),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_2),
.Y(n_289)
);

AND2x4_ASAP7_75t_L g290 ( 
.A(n_241),
.B(n_3),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_263),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_241),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_263),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_228),
.Y(n_294)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_263),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_3),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_228),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_4),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_266),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_266),
.Y(n_300)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_263),
.Y(n_301)
);

AND2x4_ASAP7_75t_L g302 ( 
.A(n_246),
.B(n_34),
.Y(n_302)
);

AND2x4_ASAP7_75t_L g303 ( 
.A(n_246),
.B(n_35),
.Y(n_303)
);

BUFx12f_ASAP7_75t_L g304 ( 
.A(n_225),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_264),
.B(n_5),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_264),
.Y(n_306)
);

AND2x4_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_208),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_277),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_209),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_225),
.B(n_5),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_225),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_211),
.B(n_7),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_222),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_217),
.B(n_8),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_221),
.B(n_8),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_272),
.Y(n_316)
);

AND2x4_ASAP7_75t_L g317 ( 
.A(n_213),
.B(n_219),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_223),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_229),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_234),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_235),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_266),
.B(n_9),
.Y(n_322)
);

AND2x4_ASAP7_75t_L g323 ( 
.A(n_238),
.B(n_36),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_266),
.B(n_239),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_233),
.B(n_9),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_266),
.B(n_10),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_240),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_212),
.B(n_10),
.Y(n_328)
);

BUFx12f_ASAP7_75t_L g329 ( 
.A(n_249),
.Y(n_329)
);

INVx5_ASAP7_75t_L g330 ( 
.A(n_212),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_256),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_227),
.B(n_11),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_243),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_266),
.B(n_11),
.Y(n_334)
);

BUFx8_ASAP7_75t_L g335 ( 
.A(n_266),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_280),
.B(n_247),
.Y(n_336)
);

AND2x4_ASAP7_75t_L g337 ( 
.A(n_261),
.B(n_12),
.Y(n_337)
);

AND2x4_ASAP7_75t_L g338 ( 
.A(n_286),
.B(n_267),
.Y(n_338)
);

OAI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_298),
.A2(n_279),
.B1(n_278),
.B2(n_273),
.Y(n_339)
);

AO22x2_ASAP7_75t_L g340 ( 
.A1(n_325),
.A2(n_268),
.B1(n_271),
.B2(n_281),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_293),
.Y(n_341)
);

OA22x2_ASAP7_75t_L g342 ( 
.A1(n_331),
.A2(n_283),
.B1(n_282),
.B2(n_276),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_204),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_293),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_328),
.A2(n_218),
.B1(n_250),
.B2(n_252),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_330),
.B(n_205),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_293),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_292),
.B(n_13),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_325),
.A2(n_244),
.B1(n_274),
.B2(n_269),
.Y(n_349)
);

AO22x2_ASAP7_75t_L g350 ( 
.A1(n_310),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_350)
);

OAI22xp33_ASAP7_75t_L g351 ( 
.A1(n_287),
.A2(n_275),
.B1(n_265),
.B2(n_262),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_296),
.A2(n_260),
.B1(n_259),
.B2(n_258),
.Y(n_352)
);

OA22x2_ASAP7_75t_L g353 ( 
.A1(n_313),
.A2(n_257),
.B1(n_255),
.B2(n_254),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_329),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_296),
.A2(n_253),
.B1(n_251),
.B2(n_248),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_332),
.A2(n_224),
.B1(n_242),
.B2(n_236),
.Y(n_356)
);

AND2x2_ASAP7_75t_SL g357 ( 
.A(n_305),
.B(n_216),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_330),
.B(n_206),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_293),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_306),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_306),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_312),
.A2(n_245),
.B1(n_232),
.B2(n_231),
.Y(n_362)
);

AO22x2_ASAP7_75t_L g363 ( 
.A1(n_288),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_L g364 ( 
.A1(n_311),
.A2(n_230),
.B1(n_226),
.B2(n_220),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_330),
.B(n_207),
.Y(n_365)
);

OAI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_336),
.A2(n_322),
.B1(n_326),
.B2(n_334),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_332),
.A2(n_215),
.B1(n_214),
.B2(n_210),
.Y(n_367)
);

OAI22xp33_ASAP7_75t_L g368 ( 
.A1(n_311),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_368)
);

OAI22xp33_ASAP7_75t_L g369 ( 
.A1(n_304),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_369)
);

OAI22xp33_ASAP7_75t_L g370 ( 
.A1(n_304),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_306),
.Y(n_371)
);

OAI22xp33_ASAP7_75t_R g372 ( 
.A1(n_336),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_292),
.B(n_37),
.Y(n_373)
);

OAI22xp33_ASAP7_75t_L g374 ( 
.A1(n_289),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_307),
.B(n_39),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_289),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_307),
.B(n_41),
.Y(n_377)
);

OAI22xp33_ASAP7_75t_L g378 ( 
.A1(n_329),
.A2(n_27),
.B1(n_43),
.B2(n_44),
.Y(n_378)
);

OAI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_288),
.A2(n_45),
.B1(n_46),
.B2(n_49),
.Y(n_379)
);

OAI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_290),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_314),
.A2(n_315),
.B1(n_302),
.B2(n_303),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_307),
.B(n_53),
.Y(n_382)
);

OAI22xp33_ASAP7_75t_L g383 ( 
.A1(n_324),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_317),
.B(n_306),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_308),
.B(n_58),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_308),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_308),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_308),
.Y(n_388)
);

AND2x2_ASAP7_75t_SL g389 ( 
.A(n_290),
.B(n_59),
.Y(n_389)
);

OAI22xp33_ASAP7_75t_L g390 ( 
.A1(n_316),
.A2(n_60),
.B1(n_61),
.B2(n_65),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_309),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_286),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_361),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_361),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_345),
.B(n_286),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_360),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_386),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_387),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_345),
.Y(n_399)
);

XOR2x2_ASAP7_75t_L g400 ( 
.A(n_362),
.B(n_337),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_366),
.B(n_317),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_381),
.A2(n_323),
.B(n_303),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_389),
.B(n_302),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_388),
.Y(n_404)
);

XNOR2x2_ASAP7_75t_L g405 ( 
.A(n_350),
.B(n_320),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_391),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_391),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_349),
.B(n_302),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_357),
.B(n_356),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_347),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_338),
.A2(n_321),
.B(n_333),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_349),
.B(n_303),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_371),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_341),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_341),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_344),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_344),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_371),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_371),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_359),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_359),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_385),
.Y(n_422)
);

XOR2x2_ASAP7_75t_L g423 ( 
.A(n_339),
.B(n_337),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_348),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_375),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_377),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_382),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_354),
.B(n_323),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_338),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_342),
.B(n_323),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_373),
.Y(n_431)
);

INVxp33_ASAP7_75t_L g432 ( 
.A(n_367),
.Y(n_432)
);

NOR2xp67_ASAP7_75t_L g433 ( 
.A(n_356),
.B(n_295),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_353),
.Y(n_434)
);

AND2x6_ASAP7_75t_L g435 ( 
.A(n_376),
.B(n_343),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_340),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_340),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_346),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_352),
.B(n_327),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_352),
.B(n_294),
.Y(n_440)
);

NOR2xp67_ASAP7_75t_L g441 ( 
.A(n_355),
.B(n_295),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_358),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_365),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_379),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_363),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_380),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_363),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_350),
.B(n_66),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_390),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_376),
.B(n_294),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_378),
.B(n_297),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_351),
.B(n_67),
.Y(n_452)
);

XNOR2x2_ASAP7_75t_L g453 ( 
.A(n_372),
.B(n_299),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_364),
.B(n_68),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_374),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_368),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_383),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_369),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_370),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_356),
.B(n_295),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_347),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_440),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_401),
.A2(n_300),
.B(n_299),
.Y(n_463)
);

NOR2xp67_ASAP7_75t_L g464 ( 
.A(n_431),
.B(n_291),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_422),
.B(n_297),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_392),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_392),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_429),
.B(n_70),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_436),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_424),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_429),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_410),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_410),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_439),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_438),
.B(n_300),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_442),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_461),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_461),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_408),
.B(n_412),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_421),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_408),
.B(n_309),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_420),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_443),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_412),
.B(n_402),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_426),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_421),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_420),
.Y(n_487)
);

AND2x2_ASAP7_75t_SL g488 ( 
.A(n_409),
.B(n_291),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_402),
.B(n_309),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_435),
.A2(n_319),
.B1(n_318),
.B2(n_309),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_435),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_406),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_434),
.B(n_72),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_426),
.Y(n_494)
);

INVx4_ASAP7_75t_L g495 ( 
.A(n_426),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_407),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_414),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_415),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_435),
.A2(n_319),
.B1(n_318),
.B2(n_335),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_454),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_450),
.B(n_318),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_450),
.B(n_318),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_418),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_403),
.B(n_319),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_426),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_403),
.B(n_319),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_416),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_417),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_428),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_419),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_425),
.B(n_335),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_437),
.B(n_295),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_444),
.B(n_73),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_401),
.A2(n_301),
.B(n_76),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_427),
.B(n_301),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_399),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_433),
.B(n_301),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_396),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_446),
.B(n_75),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_397),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_445),
.B(n_301),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_413),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_398),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_404),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_460),
.B(n_77),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_435),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_445),
.B(n_79),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_393),
.Y(n_528)
);

INVx1_ASAP7_75t_SL g529 ( 
.A(n_430),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_423),
.Y(n_530)
);

NOR2xp67_ASAP7_75t_L g531 ( 
.A(n_394),
.B(n_81),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_447),
.B(n_82),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_457),
.A2(n_83),
.B(n_85),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_478),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_471),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_476),
.B(n_451),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_478),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_476),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_471),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_501),
.B(n_451),
.Y(n_540)
);

NAND2x1p5_ASAP7_75t_L g541 ( 
.A(n_485),
.B(n_413),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_474),
.B(n_395),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_479),
.B(n_432),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_467),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_465),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_484),
.B(n_435),
.Y(n_546)
);

INVx5_ASAP7_75t_L g547 ( 
.A(n_467),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_462),
.B(n_432),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_465),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_470),
.B(n_458),
.Y(n_550)
);

BUFx4f_ASAP7_75t_L g551 ( 
.A(n_493),
.Y(n_551)
);

OR2x6_ASAP7_75t_L g552 ( 
.A(n_491),
.B(n_447),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_467),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_501),
.B(n_449),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_484),
.B(n_411),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_481),
.B(n_411),
.Y(n_556)
);

NAND2x1p5_ASAP7_75t_L g557 ( 
.A(n_485),
.B(n_441),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_502),
.B(n_458),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_530),
.B(n_459),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_487),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_SL g561 ( 
.A(n_500),
.B(n_455),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_483),
.B(n_456),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_467),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_502),
.B(n_86),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_473),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_487),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_483),
.B(n_405),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_466),
.B(n_87),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_516),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_SL g570 ( 
.A(n_500),
.B(n_488),
.Y(n_570)
);

OR2x6_ASAP7_75t_L g571 ( 
.A(n_491),
.B(n_448),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_466),
.B(n_88),
.Y(n_572)
);

NOR2x1_ASAP7_75t_L g573 ( 
.A(n_485),
.B(n_452),
.Y(n_573)
);

BUFx12f_ASAP7_75t_L g574 ( 
.A(n_493),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_469),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_SL g576 ( 
.A(n_488),
.B(n_400),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_481),
.B(n_480),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_L g578 ( 
.A(n_467),
.B(n_453),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_486),
.B(n_89),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_486),
.B(n_90),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_473),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_468),
.Y(n_582)
);

NOR2x1_ASAP7_75t_R g583 ( 
.A(n_493),
.B(n_91),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_468),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_489),
.B(n_92),
.Y(n_585)
);

AND2x6_ASAP7_75t_L g586 ( 
.A(n_499),
.B(n_94),
.Y(n_586)
);

OR2x6_ASAP7_75t_L g587 ( 
.A(n_526),
.B(n_97),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_468),
.B(n_98),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_492),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_SL g590 ( 
.A(n_488),
.B(n_99),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_489),
.B(n_101),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_477),
.Y(n_592)
);

INVxp67_ASAP7_75t_SL g593 ( 
.A(n_582),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_534),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_569),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_582),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_543),
.B(n_526),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_534),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_537),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_537),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g601 ( 
.A1(n_551),
.A2(n_499),
.B1(n_504),
.B2(n_490),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_582),
.Y(n_602)
);

INVx3_ASAP7_75t_SL g603 ( 
.A(n_587),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_538),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_584),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_584),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_584),
.Y(n_607)
);

BUFx6f_ASAP7_75t_SL g608 ( 
.A(n_536),
.Y(n_608)
);

CKINVDCx6p67_ASAP7_75t_R g609 ( 
.A(n_574),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_544),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_544),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_545),
.Y(n_612)
);

INVx8_ASAP7_75t_L g613 ( 
.A(n_586),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_565),
.Y(n_614)
);

BUFx2_ASAP7_75t_SL g615 ( 
.A(n_547),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_581),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_592),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_547),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_558),
.B(n_527),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_560),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_544),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_566),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_589),
.Y(n_623)
);

BUFx10_ASAP7_75t_L g624 ( 
.A(n_548),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_552),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_552),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_577),
.B(n_475),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_554),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_536),
.Y(n_629)
);

INVx5_ASAP7_75t_L g630 ( 
.A(n_553),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_553),
.Y(n_631)
);

CKINVDCx14_ASAP7_75t_R g632 ( 
.A(n_559),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_553),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_554),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_563),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_535),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_587),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_539),
.Y(n_638)
);

BUFx4_ASAP7_75t_SL g639 ( 
.A(n_571),
.Y(n_639)
);

CKINVDCx16_ASAP7_75t_R g640 ( 
.A(n_570),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_540),
.Y(n_641)
);

OAI22xp33_ASAP7_75t_L g642 ( 
.A1(n_640),
.A2(n_576),
.B1(n_590),
.B2(n_561),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_632),
.A2(n_542),
.B1(n_573),
.B2(n_578),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_623),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_598),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_623),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_618),
.Y(n_647)
);

INVx6_ASAP7_75t_L g648 ( 
.A(n_629),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_622),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_597),
.A2(n_529),
.B1(n_546),
.B2(n_540),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_622),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_620),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_619),
.A2(n_551),
.B1(n_567),
.B2(n_562),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_620),
.Y(n_654)
);

INVx4_ASAP7_75t_L g655 ( 
.A(n_630),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_611),
.Y(n_656)
);

BUFx2_ASAP7_75t_SL g657 ( 
.A(n_604),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_598),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_600),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_600),
.Y(n_660)
);

CKINVDCx11_ASAP7_75t_R g661 ( 
.A(n_609),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_SL g662 ( 
.A1(n_640),
.A2(n_586),
.B1(n_588),
.B2(n_571),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_594),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_595),
.Y(n_664)
);

BUFx12f_ASAP7_75t_L g665 ( 
.A(n_595),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_619),
.A2(n_586),
.B1(n_533),
.B2(n_555),
.Y(n_666)
);

INVx1_ASAP7_75t_SL g667 ( 
.A(n_604),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_594),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_SL g669 ( 
.A1(n_613),
.A2(n_586),
.B1(n_588),
.B2(n_513),
.Y(n_669)
);

BUFx10_ASAP7_75t_L g670 ( 
.A(n_608),
.Y(n_670)
);

OAI22xp33_ASAP7_75t_L g671 ( 
.A1(n_603),
.A2(n_490),
.B1(n_549),
.B2(n_556),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_599),
.Y(n_672)
);

OAI22xp5_ASAP7_75t_L g673 ( 
.A1(n_601),
.A2(n_557),
.B1(n_547),
.B2(n_564),
.Y(n_673)
);

CKINVDCx6p67_ASAP7_75t_R g674 ( 
.A(n_609),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_599),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_626),
.Y(n_676)
);

INVx6_ASAP7_75t_L g677 ( 
.A(n_629),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_613),
.A2(n_514),
.B1(n_519),
.B2(n_513),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_625),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_630),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_627),
.B(n_550),
.Y(n_681)
);

INVx6_ASAP7_75t_L g682 ( 
.A(n_629),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_616),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_625),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_684),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_643),
.B(n_624),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_664),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_642),
.A2(n_603),
.B1(n_637),
.B2(n_634),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_645),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_642),
.A2(n_624),
.B1(n_613),
.B2(n_637),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g691 ( 
.A1(n_678),
.A2(n_603),
.B1(n_634),
.B2(n_628),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_645),
.Y(n_692)
);

OAI21xp33_ASAP7_75t_L g693 ( 
.A1(n_681),
.A2(n_511),
.B(n_628),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_662),
.B(n_624),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_SL g695 ( 
.A1(n_653),
.A2(n_613),
.B1(n_624),
.B2(n_516),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_649),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_662),
.A2(n_613),
.B1(n_513),
.B2(n_519),
.Y(n_697)
);

OAI21xp33_ASAP7_75t_L g698 ( 
.A1(n_650),
.A2(n_666),
.B(n_678),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_676),
.B(n_636),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_644),
.B(n_612),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_666),
.A2(n_513),
.B1(n_519),
.B2(n_496),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_667),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_669),
.A2(n_492),
.B1(n_496),
.B2(n_564),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_646),
.B(n_612),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_663),
.Y(n_705)
);

OAI222xp33_ASAP7_75t_L g706 ( 
.A1(n_669),
.A2(n_638),
.B1(n_636),
.B2(n_509),
.C1(n_580),
.C2(n_579),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_647),
.Y(n_707)
);

BUFx12f_ASAP7_75t_L g708 ( 
.A(n_661),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_671),
.A2(n_638),
.B1(n_614),
.B2(n_608),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_671),
.A2(n_652),
.B1(n_654),
.B2(n_651),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g711 ( 
.A1(n_673),
.A2(n_641),
.B1(n_593),
.B2(n_608),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_679),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_672),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_661),
.Y(n_714)
);

NAND3xp33_ASAP7_75t_L g715 ( 
.A(n_675),
.B(n_464),
.C(n_520),
.Y(n_715)
);

INVx5_ASAP7_75t_SL g716 ( 
.A(n_674),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_663),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_658),
.A2(n_614),
.B1(n_520),
.B2(n_523),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_647),
.Y(n_719)
);

OAI21xp5_ASAP7_75t_SL g720 ( 
.A1(n_668),
.A2(n_525),
.B(n_591),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_656),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_668),
.B(n_575),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_659),
.B(n_641),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_679),
.B(n_527),
.Y(n_724)
);

OAI22xp33_ASAP7_75t_L g725 ( 
.A1(n_660),
.A2(n_585),
.B1(n_616),
.B2(n_617),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_L g726 ( 
.A1(n_657),
.A2(n_568),
.B1(n_572),
.B2(n_605),
.Y(n_726)
);

AOI222xp33_ASAP7_75t_L g727 ( 
.A1(n_665),
.A2(n_583),
.B1(n_475),
.B2(n_532),
.C1(n_463),
.C2(n_572),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_683),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_683),
.A2(n_523),
.B1(n_507),
.B2(n_498),
.Y(n_729)
);

CKINVDCx11_ASAP7_75t_R g730 ( 
.A(n_670),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_656),
.Y(n_731)
);

OAI22xp33_ASAP7_75t_L g732 ( 
.A1(n_648),
.A2(n_617),
.B1(n_596),
.B2(n_605),
.Y(n_732)
);

AOI211xp5_ASAP7_75t_L g733 ( 
.A1(n_656),
.A2(n_532),
.B(n_568),
.C(n_464),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_670),
.A2(n_507),
.B1(n_508),
.B2(n_498),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_722),
.B(n_648),
.Y(n_735)
);

OAI221xp5_ASAP7_75t_L g736 ( 
.A1(n_693),
.A2(n_506),
.B1(n_605),
.B2(n_518),
.C(n_497),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_705),
.B(n_656),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_697),
.A2(n_733),
.B1(n_690),
.B2(n_701),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_713),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_696),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_698),
.A2(n_508),
.B1(n_497),
.B2(n_518),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_SL g742 ( 
.A1(n_686),
.A2(n_682),
.B1(n_648),
.B2(n_677),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_727),
.A2(n_510),
.B1(n_503),
.B2(n_494),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_697),
.A2(n_682),
.B1(n_677),
.B2(n_596),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_690),
.A2(n_701),
.B1(n_695),
.B2(n_703),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_694),
.A2(n_510),
.B1(n_503),
.B2(n_494),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_691),
.A2(n_494),
.B1(n_682),
.B2(n_677),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_705),
.B(n_610),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_702),
.B(n_602),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_717),
.B(n_610),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_728),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_688),
.A2(n_528),
.B1(n_596),
.B2(n_602),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_709),
.A2(n_528),
.B1(n_602),
.B2(n_606),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_689),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_709),
.A2(n_703),
.B1(n_711),
.B2(n_724),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_685),
.A2(n_602),
.B1(n_606),
.B2(n_607),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_SL g757 ( 
.A1(n_726),
.A2(n_615),
.B1(n_680),
.B2(n_602),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_730),
.A2(n_710),
.B1(n_708),
.B2(n_734),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_710),
.B(n_610),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_SL g760 ( 
.A1(n_712),
.A2(n_615),
.B1(n_680),
.B2(n_607),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_699),
.B(n_606),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_692),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_734),
.A2(n_606),
.B1(n_607),
.B2(n_495),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_SL g764 ( 
.A1(n_716),
.A2(n_607),
.B1(n_606),
.B2(n_639),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_SL g765 ( 
.A1(n_716),
.A2(n_607),
.B1(n_635),
.B2(n_655),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_715),
.A2(n_505),
.B1(n_495),
.B2(n_524),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_723),
.A2(n_718),
.B1(n_732),
.B2(n_725),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_687),
.A2(n_563),
.B1(n_495),
.B2(n_505),
.Y(n_768)
);

NAND2xp33_ASAP7_75t_SL g769 ( 
.A(n_700),
.B(n_655),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_718),
.A2(n_505),
.B1(n_524),
.B2(n_522),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_729),
.A2(n_635),
.B1(n_618),
.B2(n_621),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_729),
.A2(n_635),
.B1(n_618),
.B2(n_621),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_739),
.B(n_731),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_735),
.B(n_704),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_761),
.B(n_725),
.Y(n_775)
);

OAI21xp33_ASAP7_75t_L g776 ( 
.A1(n_758),
.A2(n_720),
.B(n_515),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_740),
.B(n_721),
.Y(n_777)
);

OAI221xp5_ASAP7_75t_SL g778 ( 
.A1(n_755),
.A2(n_732),
.B1(n_706),
.B2(n_719),
.C(n_707),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_737),
.B(n_721),
.Y(n_779)
);

OA21x2_ASAP7_75t_L g780 ( 
.A1(n_767),
.A2(n_531),
.B(n_517),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_737),
.B(n_707),
.Y(n_781)
);

OAI221xp5_ASAP7_75t_L g782 ( 
.A1(n_745),
.A2(n_714),
.B1(n_719),
.B2(n_531),
.C(n_524),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_749),
.B(n_716),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_751),
.B(n_631),
.Y(n_784)
);

NAND3xp33_ASAP7_75t_L g785 ( 
.A(n_738),
.B(n_742),
.C(n_743),
.Y(n_785)
);

NAND2xp33_ASAP7_75t_L g786 ( 
.A(n_747),
.B(n_630),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_759),
.B(n_754),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_764),
.A2(n_630),
.B1(n_631),
.B2(n_633),
.Y(n_788)
);

AOI221xp5_ASAP7_75t_L g789 ( 
.A1(n_769),
.A2(n_512),
.B1(n_522),
.B2(n_521),
.C(n_477),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_762),
.B(n_754),
.Y(n_790)
);

NAND3xp33_ASAP7_75t_L g791 ( 
.A(n_741),
.B(n_633),
.C(n_611),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_SL g792 ( 
.A1(n_768),
.A2(n_631),
.B(n_512),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_759),
.B(n_611),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_757),
.B(n_611),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_769),
.B(n_760),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_750),
.B(n_611),
.Y(n_796)
);

NOR2xp67_ASAP7_75t_L g797 ( 
.A(n_736),
.B(n_630),
.Y(n_797)
);

OAI221xp5_ASAP7_75t_L g798 ( 
.A1(n_746),
.A2(n_541),
.B1(n_482),
.B2(n_633),
.C(n_472),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_SL g799 ( 
.A1(n_753),
.A2(n_633),
.B(n_521),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_748),
.B(n_633),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_748),
.B(n_102),
.Y(n_801)
);

NAND3xp33_ASAP7_75t_L g802 ( 
.A(n_752),
.B(n_482),
.C(n_630),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_782),
.B(n_795),
.Y(n_803)
);

NAND3xp33_ASAP7_75t_L g804 ( 
.A(n_785),
.B(n_756),
.C(n_765),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_787),
.B(n_750),
.Y(n_805)
);

AOI211xp5_ASAP7_75t_L g806 ( 
.A1(n_778),
.A2(n_744),
.B(n_771),
.C(n_772),
.Y(n_806)
);

AO21x2_ASAP7_75t_L g807 ( 
.A1(n_795),
.A2(n_766),
.B(n_763),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_773),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_780),
.A2(n_770),
.B1(n_472),
.B2(n_107),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_787),
.B(n_104),
.Y(n_810)
);

NAND3xp33_ASAP7_75t_L g811 ( 
.A(n_776),
.B(n_472),
.C(n_112),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_779),
.B(n_106),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_774),
.B(n_113),
.Y(n_813)
);

NOR3xp33_ASAP7_75t_L g814 ( 
.A(n_792),
.B(n_115),
.C(n_117),
.Y(n_814)
);

NAND3xp33_ASAP7_75t_L g815 ( 
.A(n_789),
.B(n_119),
.C(n_121),
.Y(n_815)
);

NAND3xp33_ASAP7_75t_L g816 ( 
.A(n_775),
.B(n_124),
.C(n_127),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_780),
.A2(n_128),
.B1(n_129),
.B2(n_131),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_797),
.A2(n_133),
.B(n_134),
.Y(n_818)
);

AO21x2_ASAP7_75t_L g819 ( 
.A1(n_794),
.A2(n_135),
.B(n_137),
.Y(n_819)
);

NAND3xp33_ASAP7_75t_SL g820 ( 
.A(n_783),
.B(n_138),
.C(n_140),
.Y(n_820)
);

AO21x2_ASAP7_75t_L g821 ( 
.A1(n_794),
.A2(n_143),
.B(n_144),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_780),
.A2(n_145),
.B1(n_146),
.B2(n_148),
.Y(n_822)
);

NAND4xp75_ASAP7_75t_SL g823 ( 
.A(n_803),
.B(n_801),
.C(n_800),
.D(n_777),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_805),
.B(n_779),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_808),
.B(n_781),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_808),
.B(n_773),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_803),
.B(n_777),
.Y(n_827)
);

XNOR2xp5_ASAP7_75t_L g828 ( 
.A(n_812),
.B(n_793),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_812),
.Y(n_829)
);

XNOR2x1_ASAP7_75t_L g830 ( 
.A(n_804),
.B(n_788),
.Y(n_830)
);

INVx4_ASAP7_75t_L g831 ( 
.A(n_819),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_810),
.B(n_790),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_807),
.B(n_796),
.Y(n_833)
);

INVx1_ASAP7_75t_SL g834 ( 
.A(n_833),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_824),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_826),
.Y(n_836)
);

XNOR2xp5_ASAP7_75t_L g837 ( 
.A(n_828),
.B(n_806),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_830),
.A2(n_822),
.B1(n_817),
.B2(n_811),
.Y(n_838)
);

XNOR2x1_ASAP7_75t_L g839 ( 
.A(n_830),
.B(n_813),
.Y(n_839)
);

OA22x2_ASAP7_75t_L g840 ( 
.A1(n_837),
.A2(n_829),
.B1(n_827),
.B2(n_831),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_838),
.A2(n_839),
.B1(n_822),
.B2(n_817),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_834),
.Y(n_842)
);

BUFx2_ASAP7_75t_L g843 ( 
.A(n_835),
.Y(n_843)
);

OA22x2_ASAP7_75t_L g844 ( 
.A1(n_834),
.A2(n_829),
.B1(n_827),
.B2(n_831),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_842),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_843),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_844),
.Y(n_847)
);

NOR2x1_ASAP7_75t_L g848 ( 
.A(n_841),
.B(n_831),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_846),
.Y(n_849)
);

OA22x2_ASAP7_75t_L g850 ( 
.A1(n_847),
.A2(n_840),
.B1(n_836),
.B2(n_818),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_848),
.A2(n_845),
.B1(n_814),
.B2(n_819),
.Y(n_851)
);

INVx1_ASAP7_75t_SL g852 ( 
.A(n_849),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_850),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_851),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_849),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_855),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_853),
.B(n_832),
.Y(n_857)
);

NOR3xp33_ASAP7_75t_L g858 ( 
.A(n_854),
.B(n_820),
.C(n_816),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_852),
.A2(n_855),
.B1(n_821),
.B2(n_807),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_855),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_853),
.A2(n_821),
.B1(n_815),
.B2(n_832),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_853),
.B(n_826),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_860),
.Y(n_863)
);

NOR3xp33_ASAP7_75t_SL g864 ( 
.A(n_857),
.B(n_799),
.C(n_798),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_858),
.A2(n_786),
.B1(n_809),
.B2(n_784),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_862),
.Y(n_866)
);

INVxp67_ASAP7_75t_SL g867 ( 
.A(n_856),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_859),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_861),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_867),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_866),
.A2(n_809),
.B1(n_786),
.B2(n_825),
.Y(n_871)
);

NAND4xp25_ASAP7_75t_L g872 ( 
.A(n_869),
.B(n_823),
.C(n_802),
.D(n_791),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_863),
.Y(n_873)
);

AO22x1_ASAP7_75t_L g874 ( 
.A1(n_868),
.A2(n_149),
.B1(n_150),
.B2(n_155),
.Y(n_874)
);

AO22x2_ASAP7_75t_L g875 ( 
.A1(n_864),
.A2(n_865),
.B1(n_158),
.B2(n_160),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_863),
.Y(n_876)
);

INVxp67_ASAP7_75t_SL g877 ( 
.A(n_870),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_876),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_873),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_875),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_874),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_872),
.A2(n_157),
.B1(n_161),
.B2(n_162),
.Y(n_882)
);

INVxp67_ASAP7_75t_SL g883 ( 
.A(n_871),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_870),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_881),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_880),
.A2(n_168),
.B1(n_169),
.B2(n_175),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_877),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_878),
.A2(n_176),
.B1(n_177),
.B2(n_179),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_877),
.Y(n_889)
);

OAI22x1_ASAP7_75t_L g890 ( 
.A1(n_883),
.A2(n_884),
.B1(n_882),
.B2(n_879),
.Y(n_890)
);

OAI22x1_ASAP7_75t_L g891 ( 
.A1(n_881),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_887),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_889),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_890),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_891),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_885),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_SL g897 ( 
.A1(n_894),
.A2(n_888),
.B1(n_886),
.B2(n_188),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_895),
.A2(n_186),
.B1(n_187),
.B2(n_189),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_897),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_898),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_899),
.A2(n_896),
.B1(n_893),
.B2(n_892),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_901),
.Y(n_902)
);

AOI221xp5_ASAP7_75t_L g903 ( 
.A1(n_902),
.A2(n_900),
.B1(n_191),
.B2(n_194),
.C(n_195),
.Y(n_903)
);

AOI31xp33_ASAP7_75t_L g904 ( 
.A1(n_903),
.A2(n_190),
.A3(n_196),
.B(n_197),
.Y(n_904)
);


endmodule