module fake_jpeg_2928_n_229 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_229);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_0),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g71 ( 
.A(n_9),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_6),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_17),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_8),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_1),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_6),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_24),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_11),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_0),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_71),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_1),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_88),
.Y(n_94)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_53),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_59),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_2),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_84),
.Y(n_92)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_101),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_103),
.Y(n_117)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVxp67_ASAP7_75t_SL g118 ( 
.A(n_98),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_86),
.A2(n_77),
.B1(n_78),
.B2(n_76),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_67),
.B1(n_76),
.B2(n_86),
.Y(n_114)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_62),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_110),
.B(n_119),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_87),
.Y(n_111)
);

XNOR2x1_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_63),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_101),
.A2(n_77),
.B1(n_59),
.B2(n_61),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_93),
.C(n_68),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_118),
.C(n_105),
.Y(n_138)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_81),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_120),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_81),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_95),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_67),
.B1(n_61),
.B2(n_79),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_121),
.A2(n_73),
.B1(n_74),
.B2(n_58),
.Y(n_134)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_80),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_57),
.Y(n_143)
);

AO21x2_ASAP7_75t_SL g127 ( 
.A1(n_119),
.A2(n_56),
.B(n_71),
.Y(n_127)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_56),
.B(n_63),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_131),
.B(n_136),
.Y(n_147)
);

AO22x1_ASAP7_75t_SL g132 ( 
.A1(n_111),
.A2(n_74),
.B1(n_63),
.B2(n_90),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_4),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_64),
.B1(n_109),
.B2(n_75),
.Y(n_152)
);

OAI32xp33_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_60),
.A3(n_64),
.B1(n_58),
.B2(n_5),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_139),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_124),
.A2(n_117),
.B(n_113),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_66),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_141),
.B(n_143),
.Y(n_157)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_2),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_146),
.B(n_27),
.Y(n_154)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_137),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_154),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_160),
.B1(n_170),
.B2(n_30),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_75),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_156),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_60),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_28),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_3),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_161),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_26),
.B1(n_51),
.B2(n_50),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_3),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_162),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_52),
.Y(n_163)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_163),
.A2(n_166),
.B(n_168),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_133),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_164),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_131),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_127),
.B(n_5),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_7),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_10),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_125),
.A2(n_23),
.B1(n_48),
.B2(n_47),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_129),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_171),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_165),
.A2(n_129),
.B(n_132),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_147),
.C(n_158),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_184),
.B1(n_190),
.B2(n_170),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_179),
.B(n_147),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_182),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_12),
.Y(n_181)
);

OAI322xp33_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_157),
.A3(n_163),
.B1(n_16),
.B2(n_17),
.C1(n_18),
.C2(n_19),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_153),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_166),
.A2(n_49),
.B(n_22),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_186),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_148),
.A2(n_12),
.B(n_13),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_188),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_46),
.B(n_31),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_189),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_150),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_190)
);

NOR3xp33_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_197),
.C(n_14),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_193),
.A2(n_175),
.B1(n_190),
.B2(n_188),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_202),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_183),
.C(n_187),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_198),
.C(n_186),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_155),
.C(n_160),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_181),
.B(n_150),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_203),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_206),
.C(n_208),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_176),
.C(n_191),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_178),
.C(n_177),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_174),
.C(n_180),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_209),
.B(n_198),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_41),
.B(n_44),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_20),
.Y(n_218)
);

NOR3xp33_ASAP7_75t_SL g213 ( 
.A(n_212),
.B(n_194),
.C(n_202),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_213),
.B(n_215),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_211),
.B(n_15),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_218),
.C(n_207),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_221),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_212),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_218),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_221),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_223),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_217),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_32),
.B(n_42),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_43),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_45),
.Y(n_229)
);


endmodule