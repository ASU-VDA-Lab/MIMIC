module real_jpeg_18064_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_17;
wire n_21;
wire n_10;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_22;
wire n_18;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_16;
wire n_15;
wire n_13;

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_4),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_0),
.B(n_4),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_1),
.B(n_5),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_3),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_2),
.B(n_3),
.Y(n_13)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_4),
.B(n_18),
.C(n_20),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_5),
.B(n_19),
.Y(n_18)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_6),
.B(n_7),
.C(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_17),
.C(n_21),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_8),
.A2(n_15),
.B1(n_22),
.B2(n_23),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_14),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_12),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B(n_28),
.Y(n_25)
);


endmodule