module fake_jpeg_12209_n_509 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_509);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_509;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx2_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx12f_ASAP7_75t_SL g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_51),
.B(n_64),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_54),
.B(n_97),
.Y(n_105)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_16),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_56),
.B(n_75),
.Y(n_118)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

HAxp5_ASAP7_75t_SL g58 ( 
.A(n_33),
.B(n_0),
.CON(n_58),
.SN(n_58)
);

NAND3xp33_ASAP7_75t_SL g143 ( 
.A(n_58),
.B(n_24),
.C(n_41),
.Y(n_143)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_61),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_66),
.B(n_79),
.Y(n_124)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_67),
.Y(n_144)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_69),
.Y(n_123)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_72),
.Y(n_158)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_74),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_33),
.B(n_16),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_48),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_82),
.Y(n_148)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_48),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_84),
.B(n_85),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_48),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_48),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_87),
.B(n_91),
.Y(n_147)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

BUFx16f_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_33),
.B(n_15),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_93),
.B(n_96),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_39),
.B(n_15),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_49),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_93),
.A2(n_42),
.B1(n_47),
.B2(n_18),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_102),
.A2(n_134),
.B1(n_35),
.B2(n_44),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_103),
.B(n_69),
.Y(n_159)
);

AOI21xp33_ASAP7_75t_SL g119 ( 
.A1(n_58),
.A2(n_67),
.B(n_19),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_119),
.A2(n_143),
.B(n_24),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_67),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_125),
.B(n_146),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_65),
.B(n_20),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_126),
.B(n_138),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_73),
.A2(n_42),
.B1(n_47),
.B2(n_18),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_130),
.A2(n_49),
.B1(n_42),
.B2(n_47),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_51),
.A2(n_23),
.B1(n_26),
.B2(n_18),
.Y(n_134)
);

INVx6_ASAP7_75t_SL g137 ( 
.A(n_92),
.Y(n_137)
);

INVx6_ASAP7_75t_SL g176 ( 
.A(n_137),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_80),
.B(n_20),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_68),
.B(n_37),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_139),
.B(n_154),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_57),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_60),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_149),
.B(n_152),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_92),
.B(n_41),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_59),
.B(n_37),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_159),
.B(n_168),
.Y(n_224)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_161),
.Y(n_225)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_162),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_119),
.A2(n_23),
.B1(n_26),
.B2(n_46),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_163),
.Y(n_239)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_105),
.B(n_46),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_165),
.B(n_167),
.Y(n_235)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_112),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_166),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_25),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_124),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_169),
.B(n_173),
.Y(n_214)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_171),
.Y(n_222)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_172),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_145),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_147),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_193),
.Y(n_217)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_177),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_103),
.B(n_76),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_178),
.B(n_123),
.C(n_114),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_133),
.B(n_34),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_179),
.B(n_187),
.Y(n_241)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_181),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_144),
.A2(n_26),
.B1(n_23),
.B2(n_34),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_182),
.A2(n_196),
.B1(n_201),
.B2(n_202),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_184),
.Y(n_226)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_118),
.B(n_36),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_150),
.Y(n_188)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_188),
.Y(n_253)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_122),
.Y(n_189)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_189),
.Y(n_255)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_107),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_190),
.Y(n_215)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_107),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_192),
.Y(n_247)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_131),
.Y(n_193)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_113),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_194),
.B(n_195),
.Y(n_236)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_113),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_134),
.A2(n_99),
.B1(n_53),
.B2(n_52),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_111),
.B(n_36),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_197),
.B(n_203),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_136),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_198),
.Y(n_223)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_151),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_199),
.B(n_200),
.Y(n_242)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_141),
.Y(n_200)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_140),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_106),
.A2(n_63),
.B1(n_62),
.B2(n_89),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_108),
.B(n_77),
.Y(n_203)
);

OA22x2_ASAP7_75t_L g254 ( 
.A1(n_204),
.A2(n_129),
.B1(n_121),
.B2(n_158),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_116),
.Y(n_205)
);

BUFx8_ASAP7_75t_L g237 ( 
.A(n_205),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_143),
.B(n_35),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_206),
.B(n_208),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_135),
.A2(n_95),
.B1(n_94),
.B2(n_98),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_209),
.B1(n_211),
.B2(n_212),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_151),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_144),
.A2(n_29),
.B1(n_43),
.B2(n_50),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_114),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_213),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_L g212 ( 
.A1(n_135),
.A2(n_101),
.B1(n_88),
.B2(n_74),
.Y(n_212)
);

CKINVDCx12_ASAP7_75t_R g213 ( 
.A(n_123),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_211),
.A2(n_117),
.B1(n_116),
.B2(n_156),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_227),
.A2(n_243),
.B1(n_207),
.B2(n_202),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_228),
.B(n_230),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_185),
.B(n_109),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_245),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_168),
.B(n_128),
.C(n_155),
.Y(n_230)
);

OAI32xp33_ASAP7_75t_L g231 ( 
.A1(n_191),
.A2(n_121),
.A3(n_110),
.B1(n_128),
.B2(n_142),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_231),
.B(n_248),
.Y(n_274)
);

AND2x4_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_142),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_234),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_180),
.A2(n_156),
.B1(n_117),
.B2(n_157),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_240),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_170),
.A2(n_100),
.B1(n_72),
.B2(n_81),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_190),
.A2(n_157),
.B1(n_42),
.B2(n_47),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_244),
.B(n_251),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_178),
.B(n_159),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_159),
.B(n_155),
.C(n_148),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_192),
.A2(n_158),
.B1(n_90),
.B2(n_86),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_254),
.A2(n_176),
.B1(n_186),
.B2(n_208),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_178),
.B(n_50),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_208),
.Y(n_270)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_216),
.Y(n_261)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_261),
.Y(n_302)
);

INVx13_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_262),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_263),
.A2(n_264),
.B1(n_297),
.B2(n_219),
.Y(n_321)
);

BUFx12f_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_265),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_241),
.B(n_176),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_266),
.B(n_271),
.Y(n_317)
);

AND2x6_ASAP7_75t_L g267 ( 
.A(n_224),
.B(n_212),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_267),
.B(n_268),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_217),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_249),
.A2(n_166),
.B1(n_194),
.B2(n_195),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_269),
.A2(n_277),
.B1(n_282),
.B2(n_284),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_270),
.B(n_276),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_258),
.B(n_199),
.Y(n_271)
);

AND2x6_ASAP7_75t_L g272 ( 
.A(n_224),
.B(n_161),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_272),
.B(n_280),
.Y(n_328)
);

A2O1A1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_224),
.A2(n_43),
.B(n_29),
.C(n_50),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_273),
.B(n_283),
.Y(n_306)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_275),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_235),
.B(n_172),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_239),
.A2(n_164),
.B1(n_171),
.B2(n_200),
.Y(n_277)
);

INVx13_ASAP7_75t_L g279 ( 
.A(n_233),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_279),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_242),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_239),
.A2(n_201),
.B1(n_181),
.B2(n_183),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_229),
.B(n_210),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_230),
.A2(n_205),
.B1(n_160),
.B2(n_177),
.Y(n_284)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_221),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_285),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_214),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_286),
.B(n_287),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_43),
.Y(n_287)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_225),
.Y(n_288)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_288),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_227),
.A2(n_129),
.B1(n_115),
.B2(n_174),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_289),
.B(n_293),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_245),
.B(n_110),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_290),
.A2(n_237),
.B(n_61),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_218),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_291),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_234),
.A2(n_82),
.B1(n_115),
.B2(n_49),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_292),
.A2(n_215),
.B1(n_247),
.B2(n_259),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_256),
.B(n_188),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_216),
.Y(n_294)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_294),
.Y(n_319)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_255),
.Y(n_295)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_295),
.Y(n_324)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_226),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_296),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_243),
.A2(n_232),
.B1(n_234),
.B2(n_254),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_220),
.B(n_184),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_301),
.Y(n_316)
);

INVx13_ASAP7_75t_L g301 ( 
.A(n_226),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_300),
.A2(n_218),
.B(n_228),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_303),
.A2(n_301),
.B(n_296),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_274),
.A2(n_234),
.B1(n_254),
.B2(n_248),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_305),
.A2(n_318),
.B1(n_327),
.B2(n_264),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_220),
.C(n_250),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_308),
.B(n_333),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_250),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_310),
.B(n_303),
.Y(n_343)
);

OAI32xp33_ASAP7_75t_L g311 ( 
.A1(n_260),
.A2(n_231),
.A3(n_254),
.B1(n_236),
.B2(n_219),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_311),
.B(n_291),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_313),
.A2(n_321),
.B1(n_330),
.B2(n_335),
.Y(n_351)
);

FAx1_ASAP7_75t_SL g314 ( 
.A(n_260),
.B(n_223),
.CI(n_215),
.CON(n_314),
.SN(n_314)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_314),
.B(n_287),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_278),
.A2(n_247),
.B1(n_259),
.B2(n_252),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_278),
.A2(n_252),
.B1(n_225),
.B2(n_246),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_275),
.Y(n_329)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_329),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_300),
.A2(n_246),
.B1(n_238),
.B2(n_222),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_295),
.Y(n_332)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_332),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_298),
.B(n_253),
.C(n_238),
.Y(n_333)
);

XOR2x2_ASAP7_75t_L g334 ( 
.A(n_270),
.B(n_253),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_334),
.B(n_292),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_284),
.A2(n_222),
.B1(n_29),
.B2(n_237),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_261),
.Y(n_336)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_336),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_338),
.Y(n_361)
);

INVxp33_ASAP7_75t_L g340 ( 
.A(n_317),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_340),
.B(n_358),
.Y(n_384)
);

AND2x6_ASAP7_75t_L g341 ( 
.A(n_328),
.B(n_272),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_341),
.B(n_353),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_342),
.A2(n_355),
.B1(n_363),
.B2(n_318),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_343),
.B(n_333),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_315),
.B(n_283),
.Y(n_346)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_346),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_348),
.B(n_313),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_331),
.B(n_286),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_350),
.B(n_354),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_310),
.B(n_290),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_352),
.B(n_324),
.C(n_329),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_316),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_331),
.B(n_266),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_304),
.A2(n_307),
.B1(n_326),
.B2(n_305),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_356),
.B(n_359),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_326),
.A2(n_290),
.B(n_280),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_357),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_316),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_320),
.B(n_268),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_314),
.B(n_273),
.Y(n_360)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_360),
.Y(n_377)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_309),
.Y(n_362)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_362),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_307),
.A2(n_267),
.B1(n_281),
.B2(n_269),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_314),
.B(n_288),
.Y(n_364)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_364),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_365),
.B(n_368),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_334),
.A2(n_282),
.B1(n_277),
.B2(n_271),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_366),
.A2(n_335),
.B1(n_332),
.B2(n_339),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_316),
.B(n_294),
.Y(n_367)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_367),
.Y(n_388)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_309),
.Y(n_369)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_369),
.Y(n_396)
);

OAI32xp33_ASAP7_75t_L g370 ( 
.A1(n_306),
.A2(n_285),
.A3(n_296),
.B1(n_301),
.B2(n_279),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_370),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_308),
.B(n_221),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_371),
.B(n_325),
.Y(n_392)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_324),
.Y(n_372)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_372),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_374),
.A2(n_393),
.B1(n_397),
.B2(n_351),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_375),
.B(n_380),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_357),
.A2(n_306),
.B(n_338),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_378),
.A2(n_368),
.B(n_360),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_379),
.B(n_385),
.C(n_395),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_344),
.B(n_311),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_346),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_381),
.B(n_392),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_344),
.B(n_330),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_391),
.A2(n_348),
.B1(n_366),
.B2(n_361),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_343),
.B(n_312),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_342),
.A2(n_339),
.B1(n_327),
.B2(n_312),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_367),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_399),
.B(n_354),
.Y(n_414)
);

AO22x1_ASAP7_75t_L g400 ( 
.A1(n_364),
.A2(n_337),
.B1(n_336),
.B2(n_319),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_400),
.A2(n_372),
.B(n_345),
.Y(n_417)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_345),
.Y(n_401)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_401),
.Y(n_404)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_349),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_402),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_403),
.B(n_411),
.Y(n_429)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_384),
.Y(n_405)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_405),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_406),
.B(n_415),
.Y(n_445)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_402),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_407),
.B(n_413),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_383),
.A2(n_353),
.B(n_358),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_409),
.A2(n_417),
.B(n_422),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_410),
.A2(n_412),
.B1(n_419),
.B2(n_423),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_375),
.B(n_395),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_391),
.A2(n_390),
.B1(n_383),
.B2(n_386),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_382),
.Y(n_413)
);

CKINVDCx14_ASAP7_75t_R g440 ( 
.A(n_414),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_374),
.A2(n_355),
.B1(n_363),
.B2(n_352),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_376),
.B(n_369),
.Y(n_418)
);

NOR2x1_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_421),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_374),
.A2(n_341),
.B1(n_370),
.B2(n_365),
.Y(n_419)
);

FAx1_ASAP7_75t_SL g421 ( 
.A(n_378),
.B(n_362),
.CI(n_347),
.CON(n_421),
.SN(n_421)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_389),
.A2(n_322),
.B(n_337),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_396),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_398),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_424),
.A2(n_347),
.B1(n_373),
.B2(n_349),
.Y(n_436)
);

BUFx24_ASAP7_75t_SL g425 ( 
.A(n_389),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_425),
.A2(n_387),
.B(n_373),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_385),
.B(n_379),
.C(n_380),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_427),
.B(n_394),
.C(n_377),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_430),
.B(n_435),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_408),
.B(n_394),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_431),
.B(n_433),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_411),
.B(n_397),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_408),
.B(n_388),
.C(n_393),
.Y(n_435)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_436),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_437),
.B(n_438),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_427),
.B(n_390),
.C(n_400),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_426),
.B(n_400),
.C(n_319),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_441),
.B(n_447),
.C(n_265),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_412),
.A2(n_302),
.B1(n_323),
.B2(n_285),
.Y(n_442)
);

OAI22xp33_ASAP7_75t_SL g460 ( 
.A1(n_442),
.A2(n_265),
.B1(n_1),
.B2(n_2),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_426),
.B(n_302),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_49),
.Y(n_461)
);

AOI22x1_ASAP7_75t_L g444 ( 
.A1(n_403),
.A2(n_323),
.B1(n_279),
.B2(n_262),
.Y(n_444)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_444),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_415),
.B(n_419),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_428),
.A2(n_406),
.B1(n_438),
.B2(n_439),
.Y(n_448)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_448),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_432),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_449),
.B(n_452),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_445),
.A2(n_409),
.B1(n_416),
.B2(n_421),
.Y(n_452)
);

NOR3xp33_ASAP7_75t_SL g455 ( 
.A(n_440),
.B(n_422),
.C(n_421),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_455),
.A2(n_49),
.B1(n_3),
.B2(n_4),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_445),
.A2(n_417),
.B1(n_420),
.B2(n_423),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_456),
.B(n_458),
.Y(n_472)
);

AO221x1_ASAP7_75t_L g457 ( 
.A1(n_446),
.A2(n_407),
.B1(n_434),
.B2(n_424),
.C(n_404),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_457),
.A2(n_434),
.B(n_441),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_435),
.A2(n_420),
.B1(n_265),
.B2(n_262),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_459),
.B(n_460),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_461),
.B(n_444),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_447),
.B(n_0),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_463),
.B(n_1),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_462),
.B(n_431),
.C(n_430),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_464),
.B(n_466),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_462),
.B(n_443),
.C(n_433),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_467),
.B(n_468),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_429),
.Y(n_468)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_469),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_459),
.B(n_429),
.C(n_78),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_470),
.A2(n_476),
.B(n_463),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_473),
.A2(n_463),
.B1(n_4),
.B2(n_5),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_474),
.B(n_477),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_454),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_452),
.B(n_1),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_478),
.B(n_483),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_465),
.B(n_450),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_479),
.B(n_487),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_475),
.A2(n_451),
.B(n_455),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_480),
.A2(n_485),
.B(n_477),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_456),
.C(n_458),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_484),
.B(n_474),
.Y(n_491)
);

MAJx2_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_466),
.C(n_472),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_470),
.A2(n_3),
.B(n_4),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_482),
.B(n_465),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_489),
.B(n_493),
.C(n_488),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_490),
.B(n_491),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_483),
.B(n_6),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_481),
.B(n_6),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_494),
.B(n_486),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_496),
.B(n_497),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_495),
.B(n_485),
.C(n_488),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_499),
.B(n_7),
.Y(n_502)
);

AOI31xp33_ASAP7_75t_L g501 ( 
.A1(n_498),
.A2(n_492),
.A3(n_489),
.B(n_493),
.Y(n_501)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_501),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_502),
.B(n_8),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_504),
.A2(n_500),
.B(n_9),
.Y(n_505)
);

AOI322xp5_ASAP7_75t_L g506 ( 
.A1(n_505),
.A2(n_503),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_13),
.Y(n_506)
);

OAI32xp33_ASAP7_75t_L g507 ( 
.A1(n_506),
.A2(n_8),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_507),
.B(n_11),
.Y(n_508)
);

A2O1A1Ixp33_ASAP7_75t_SL g509 ( 
.A1(n_508),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_509)
);


endmodule