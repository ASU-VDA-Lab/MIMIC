module fake_jpeg_1970_n_309 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_309);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_309;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_19),
.B(n_1),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_52),
.B(n_53),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_19),
.B(n_3),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_56),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_32),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_21),
.B(n_3),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_58),
.B(n_69),
.Y(n_124)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_60),
.Y(n_151)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_20),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_65),
.B(n_88),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_21),
.B(n_5),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_23),
.B(n_8),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_70),
.B(n_81),
.Y(n_131)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_23),
.B(n_8),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_78),
.B(n_89),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_28),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_79),
.A2(n_36),
.B1(n_47),
.B2(n_45),
.Y(n_123)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_26),
.B(n_10),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_26),
.B(n_10),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_90),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_29),
.B(n_11),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_92),
.Y(n_136)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_94),
.Y(n_138)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

BUFx16f_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_29),
.B(n_30),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_99),
.Y(n_139)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_97),
.Y(n_104)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_98),
.A2(n_39),
.B1(n_20),
.B2(n_51),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_35),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_18),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_54),
.A2(n_30),
.B1(n_36),
.B2(n_33),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_101),
.A2(n_120),
.B1(n_127),
.B2(n_128),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_102),
.A2(n_98),
.B1(n_87),
.B2(n_82),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_65),
.A2(n_20),
.B1(n_51),
.B2(n_43),
.Y(n_120)
);

AO22x2_ASAP7_75t_L g122 ( 
.A1(n_59),
.A2(n_40),
.B1(n_48),
.B2(n_43),
.Y(n_122)
);

AO22x2_ASAP7_75t_L g168 ( 
.A1(n_122),
.A2(n_149),
.B1(n_148),
.B2(n_105),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_142),
.B1(n_57),
.B2(n_64),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_66),
.A2(n_47),
.B1(n_45),
.B2(n_41),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_61),
.A2(n_33),
.B1(n_41),
.B2(n_50),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_67),
.A2(n_50),
.B1(n_48),
.B2(n_40),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_130),
.A2(n_148),
.B1(n_139),
.B2(n_128),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_141),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_80),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_95),
.B(n_12),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_145),
.B(n_131),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_90),
.B(n_18),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_86),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_73),
.A2(n_13),
.B1(n_17),
.B2(n_75),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_97),
.A2(n_17),
.B1(n_74),
.B2(n_76),
.Y(n_149)
);

OAI31xp33_ASAP7_75t_L g162 ( 
.A1(n_149),
.A2(n_82),
.A3(n_72),
.B(n_85),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_138),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_152),
.B(n_156),
.Y(n_198)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_153),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_132),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_154),
.Y(n_208)
);

BUFx2_ASAP7_75t_SL g155 ( 
.A(n_114),
.Y(n_155)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_155),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_103),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_158),
.A2(n_162),
.B1(n_182),
.B2(n_183),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_159),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_160),
.Y(n_201)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_164),
.Y(n_194)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_110),
.Y(n_166)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_106),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_167),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_168),
.B(n_171),
.Y(n_212)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_105),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_173),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_107),
.B(n_137),
.Y(n_171)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_118),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_132),
.A2(n_145),
.B(n_139),
.Y(n_174)
);

FAx1_ASAP7_75t_SL g209 ( 
.A(n_174),
.B(n_172),
.CI(n_154),
.CON(n_209),
.SN(n_209)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_112),
.B(n_116),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_180),
.C(n_181),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_114),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_176),
.A2(n_179),
.B1(n_187),
.B2(n_189),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_136),
.A2(n_149),
.B1(n_104),
.B2(n_140),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_177),
.A2(n_178),
.B1(n_133),
.B2(n_143),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_111),
.A2(n_134),
.B1(n_118),
.B2(n_124),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_134),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_102),
.A2(n_151),
.B1(n_117),
.B2(n_125),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_108),
.A2(n_115),
.B1(n_119),
.B2(n_129),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_184),
.A2(n_186),
.B1(n_173),
.B2(n_179),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_109),
.B(n_113),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_175),
.C(n_188),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_108),
.A2(n_115),
.B1(n_119),
.B2(n_133),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_129),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_121),
.Y(n_188)
);

OAI32xp33_ASAP7_75t_L g191 ( 
.A1(n_188),
.A2(n_121),
.A3(n_146),
.B1(n_144),
.B2(n_143),
.Y(n_191)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_121),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_190),
.A2(n_202),
.B1(n_166),
.B2(n_153),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_191),
.B(n_190),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_161),
.A2(n_165),
.B1(n_177),
.B2(n_158),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_170),
.A2(n_168),
.B1(n_162),
.B2(n_174),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_204),
.A2(n_208),
.B1(n_216),
.B2(n_206),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_168),
.A2(n_178),
.B1(n_186),
.B2(n_184),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_206),
.A2(n_167),
.B1(n_169),
.B2(n_187),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_209),
.A2(n_212),
.B(n_194),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_185),
.Y(n_219)
);

FAx1_ASAP7_75t_SL g216 ( 
.A(n_168),
.B(n_181),
.CI(n_175),
.CON(n_216),
.SN(n_216)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_192),
.Y(n_224)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_210),
.Y(n_217)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_218),
.A2(n_222),
.B1(n_211),
.B2(n_197),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_229),
.C(n_209),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_220),
.A2(n_232),
.B1(n_238),
.B2(n_208),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_185),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_221),
.B(n_225),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_163),
.B1(n_189),
.B2(n_205),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_223),
.Y(n_253)
);

NOR3xp33_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_237),
.C(n_215),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_200),
.B(n_205),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_226),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_199),
.B(n_209),
.Y(n_243)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_228),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_212),
.C(n_200),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_193),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_233),
.Y(n_250)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_203),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_193),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_236),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_213),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_192),
.B(n_191),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_244),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_243),
.A2(n_251),
.B(n_235),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_237),
.A2(n_216),
.B1(n_196),
.B2(n_215),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_199),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_249),
.C(n_226),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_248),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_230),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_233),
.Y(n_268)
);

XOR2x1_ASAP7_75t_SL g255 ( 
.A(n_227),
.B(n_211),
.Y(n_255)
);

OAI322xp33_ASAP7_75t_L g257 ( 
.A1(n_255),
.A2(n_224),
.A3(n_219),
.B1(n_217),
.B2(n_223),
.C1(n_232),
.C2(n_225),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_219),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_259),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_257),
.A2(n_269),
.B(n_250),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_245),
.B(n_234),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_258),
.B(n_264),
.Y(n_271)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_254),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

A2O1A1Ixp33_ASAP7_75t_SL g263 ( 
.A1(n_244),
.A2(n_220),
.B(n_222),
.C(n_218),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_268),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_228),
.C(n_231),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_266),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_255),
.C(n_240),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_267),
.B(n_250),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_213),
.B(n_235),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_262),
.A2(n_242),
.B1(n_240),
.B2(n_253),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_274),
.B1(n_239),
.B2(n_263),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_269),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_274),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_262),
.A2(n_253),
.B1(n_248),
.B2(n_235),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_276),
.A2(n_278),
.B1(n_279),
.B2(n_271),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_241),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_266),
.C(n_259),
.Y(n_281)
);

OA21x2_ASAP7_75t_SL g286 ( 
.A1(n_279),
.A2(n_260),
.B(n_280),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_286),
.C(n_275),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_280),
.A2(n_264),
.B(n_260),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_284),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_277),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_285),
.A2(n_287),
.B(n_288),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_247),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_270),
.C(n_275),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_281),
.C(n_265),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_247),
.C(n_263),
.Y(n_299)
);

NOR3xp33_ASAP7_75t_SL g293 ( 
.A(n_287),
.B(n_245),
.C(n_273),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_293),
.A2(n_292),
.B1(n_294),
.B2(n_239),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_291),
.A2(n_283),
.B(n_285),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_295),
.B(n_297),
.Y(n_302)
);

NOR2x1_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_299),
.Y(n_300)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_293),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_298),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_302),
.B(n_296),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_304),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_289),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_300),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_305),
.B(n_263),
.C(n_195),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_307),
.B(n_305),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_306),
.Y(n_309)
);


endmodule