module real_aes_6322_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_119;
wire n_310;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_183;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_393;
wire n_294;
wire n_84;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
A2O1A1Ixp33_ASAP7_75t_L g101 ( .A1(n_0), .A2(n_99), .B(n_102), .C(n_105), .Y(n_101) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_1), .A2(n_125), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_2), .B(n_148), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_3), .A2(n_25), .B1(n_397), .B2(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_3), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_4), .A2(n_406), .B1(n_504), .B2(n_528), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_4), .Y(n_528) );
AND2x6_ASAP7_75t_L g99 ( .A(n_5), .B(n_100), .Y(n_99) );
INVx1_ASAP7_75t_L g516 ( .A(n_5), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_5), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g132 ( .A(n_6), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g110 ( .A(n_7), .B(n_111), .Y(n_110) );
AO22x2_ASAP7_75t_L g425 ( .A1(n_8), .A2(n_28), .B1(n_417), .B2(n_422), .Y(n_425) );
INVx1_ASAP7_75t_L g91 ( .A(n_9), .Y(n_91) );
A2O1A1Ixp33_ASAP7_75t_L g142 ( .A1(n_10), .A2(n_133), .B(n_143), .C(n_146), .Y(n_142) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_11), .A2(n_56), .B1(n_434), .B2(n_438), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_12), .B(n_148), .Y(n_147) );
AO22x2_ASAP7_75t_L g427 ( .A1(n_13), .A2(n_30), .B1(n_417), .B2(n_418), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_14), .B(n_189), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g153 ( .A1(n_15), .A2(n_154), .B(n_155), .C(n_157), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_16), .B(n_111), .Y(n_211) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_17), .A2(n_71), .B1(n_411), .B2(n_428), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_18), .B(n_111), .Y(n_198) );
CKINVDCx16_ASAP7_75t_R g207 ( .A(n_19), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_19), .A2(n_207), .B1(n_406), .B2(n_504), .Y(n_518) );
INVx1_ASAP7_75t_L g197 ( .A(n_20), .Y(n_197) );
BUFx6f_ASAP7_75t_L g98 ( .A(n_21), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_22), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_23), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g184 ( .A(n_24), .Y(n_184) );
INVx1_ASAP7_75t_L g397 ( .A(n_25), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_26), .A2(n_32), .B1(n_444), .B2(n_448), .Y(n_443) );
INVx2_ASAP7_75t_L g97 ( .A(n_27), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_29), .Y(n_116) );
OAI221xp5_ASAP7_75t_L g508 ( .A1(n_30), .A2(n_45), .B1(n_55), .B2(n_509), .C(n_510), .Y(n_508) );
INVxp67_ASAP7_75t_L g511 ( .A(n_30), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g166 ( .A1(n_31), .A2(n_154), .B(n_167), .C(n_169), .Y(n_166) );
INVxp67_ASAP7_75t_L g186 ( .A(n_33), .Y(n_186) );
CKINVDCx14_ASAP7_75t_R g165 ( .A(n_34), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g195 ( .A1(n_35), .A2(n_102), .B(n_196), .C(n_200), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_36), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g129 ( .A1(n_37), .A2(n_113), .B(n_130), .C(n_131), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_38), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_39), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_40), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_41), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_42), .Y(n_500) );
INVx1_ASAP7_75t_L g152 ( .A(n_43), .Y(n_152) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_44), .A2(n_50), .B1(n_455), .B2(n_459), .Y(n_454) );
AO22x2_ASAP7_75t_L g416 ( .A1(n_45), .A2(n_67), .B1(n_417), .B2(n_418), .Y(n_416) );
INVxp67_ASAP7_75t_L g512 ( .A(n_45), .Y(n_512) );
CKINVDCx14_ASAP7_75t_R g127 ( .A(n_46), .Y(n_127) );
INVx1_ASAP7_75t_L g100 ( .A(n_47), .Y(n_100) );
INVx1_ASAP7_75t_L g90 ( .A(n_48), .Y(n_90) );
INVx1_ASAP7_75t_SL g168 ( .A(n_49), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_51), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_52), .B(n_148), .Y(n_159) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_53), .A2(n_76), .B1(n_400), .B2(n_401), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_53), .Y(n_401) );
INVx1_ASAP7_75t_L g210 ( .A(n_54), .Y(n_210) );
AO22x2_ASAP7_75t_L g421 ( .A1(n_55), .A2(n_72), .B1(n_417), .B2(n_422), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g124 ( .A1(n_57), .A2(n_125), .B(n_126), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_58), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g214 ( .A(n_59), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_60), .A2(n_125), .B(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g405 ( .A(n_60), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_61), .A2(n_179), .B(n_180), .Y(n_178) );
INVx1_ASAP7_75t_L g141 ( .A(n_62), .Y(n_141) );
CKINVDCx16_ASAP7_75t_R g194 ( .A(n_63), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_64), .A2(n_125), .B(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g144 ( .A(n_65), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_66), .Y(n_495) );
INVx2_ASAP7_75t_L g88 ( .A(n_68), .Y(n_88) );
INVx1_ASAP7_75t_L g106 ( .A(n_69), .Y(n_106) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_70), .A2(n_102), .B(n_209), .C(n_212), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_73), .B(n_118), .Y(n_135) );
INVx1_ASAP7_75t_L g417 ( .A(n_74), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_74), .Y(n_419) );
INVx2_ASAP7_75t_L g156 ( .A(n_75), .Y(n_156) );
INVx1_ASAP7_75t_L g400 ( .A(n_76), .Y(n_400) );
AOI221xp5_ASAP7_75t_SL g77 ( .A1(n_78), .A2(n_389), .B1(n_393), .B2(n_505), .C(n_517), .Y(n_77) );
OR2x2_ASAP7_75t_SL g78 ( .A(n_79), .B(n_344), .Y(n_78) );
NAND5xp2_ASAP7_75t_L g79 ( .A(n_80), .B(n_256), .C(n_294), .D(n_315), .E(n_332), .Y(n_79) );
NOR3xp33_ASAP7_75t_L g80 ( .A(n_81), .B(n_228), .C(n_249), .Y(n_80) );
OAI221xp5_ASAP7_75t_SL g81 ( .A1(n_82), .A2(n_160), .B1(n_191), .B2(n_215), .C(n_219), .Y(n_81) );
NAND2xp5_ASAP7_75t_L g82 ( .A(n_83), .B(n_120), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_84), .B(n_217), .Y(n_236) );
OR2x2_ASAP7_75t_L g263 ( .A(n_84), .B(n_137), .Y(n_263) );
AND2x2_ASAP7_75t_L g277 ( .A(n_84), .B(n_137), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_84), .B(n_123), .Y(n_291) );
AND2x2_ASAP7_75t_L g329 ( .A(n_84), .B(n_293), .Y(n_329) );
AND2x2_ASAP7_75t_L g358 ( .A(n_84), .B(n_268), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_84), .B(n_240), .Y(n_375) );
INVx4_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
AND2x2_ASAP7_75t_L g255 ( .A(n_85), .B(n_136), .Y(n_255) );
BUFx3_ASAP7_75t_L g280 ( .A(n_85), .Y(n_280) );
AND2x2_ASAP7_75t_L g309 ( .A(n_85), .B(n_137), .Y(n_309) );
AND3x2_ASAP7_75t_L g322 ( .A(n_85), .B(n_323), .C(n_324), .Y(n_322) );
AO21x2_ASAP7_75t_L g85 ( .A1(n_86), .A2(n_92), .B(n_115), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
OA21x2_ASAP7_75t_L g123 ( .A1(n_87), .A2(n_124), .B(n_135), .Y(n_123) );
INVx2_ASAP7_75t_L g190 ( .A(n_87), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_87), .A2(n_94), .B(n_194), .C(n_195), .Y(n_193) );
AND2x2_ASAP7_75t_SL g87 ( .A(n_88), .B(n_89), .Y(n_87) );
AND2x2_ASAP7_75t_L g119 ( .A(n_88), .B(n_89), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g89 ( .A(n_90), .B(n_91), .Y(n_89) );
OAI21xp5_ASAP7_75t_L g92 ( .A1(n_93), .A2(n_94), .B(n_101), .Y(n_92) );
OAI21xp5_ASAP7_75t_L g206 ( .A1(n_94), .A2(n_207), .B(n_208), .Y(n_206) );
NAND2x1p5_ASAP7_75t_L g94 ( .A(n_95), .B(n_99), .Y(n_94) );
AND2x4_ASAP7_75t_L g125 ( .A(n_95), .B(n_99), .Y(n_125) );
AND2x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_98), .Y(n_95) );
INVx1_ASAP7_75t_L g187 ( .A(n_96), .Y(n_187) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx2_ASAP7_75t_L g103 ( .A(n_97), .Y(n_103) );
INVx1_ASAP7_75t_L g158 ( .A(n_97), .Y(n_158) );
INVx1_ASAP7_75t_L g104 ( .A(n_98), .Y(n_104) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_98), .Y(n_109) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_98), .Y(n_111) );
INVx3_ASAP7_75t_L g133 ( .A(n_98), .Y(n_133) );
INVx4_ASAP7_75t_SL g134 ( .A(n_99), .Y(n_134) );
BUFx3_ASAP7_75t_L g200 ( .A(n_99), .Y(n_200) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_100), .Y(n_514) );
INVx5_ASAP7_75t_L g128 ( .A(n_102), .Y(n_128) );
AND2x6_ASAP7_75t_L g102 ( .A(n_103), .B(n_104), .Y(n_102) );
BUFx3_ASAP7_75t_L g114 ( .A(n_103), .Y(n_114) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_103), .Y(n_170) );
O2A1O1Ixp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_107), .B(n_110), .C(n_112), .Y(n_105) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_107), .A2(n_112), .B(n_210), .C(n_211), .Y(n_209) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_107), .Y(n_392) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx4_ASAP7_75t_L g145 ( .A(n_109), .Y(n_145) );
INVx2_ASAP7_75t_L g130 ( .A(n_111), .Y(n_130) );
INVx4_ASAP7_75t_L g154 ( .A(n_111), .Y(n_154) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g146 ( .A(n_114), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
INVx3_ASAP7_75t_L g148 ( .A(n_117), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_117), .B(n_202), .Y(n_201) );
AO21x2_ASAP7_75t_L g205 ( .A1(n_117), .A2(n_206), .B(n_213), .Y(n_205) );
INVx4_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_118), .Y(n_138) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g177 ( .A(n_119), .Y(n_177) );
INVx1_ASAP7_75t_L g245 ( .A(n_120), .Y(n_245) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_136), .Y(n_120) );
AOI32xp33_ASAP7_75t_L g300 ( .A1(n_121), .A2(n_252), .A3(n_301), .B1(n_304), .B2(n_305), .Y(n_300) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g227 ( .A(n_122), .B(n_136), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_122), .B(n_255), .Y(n_298) );
AND2x2_ASAP7_75t_L g305 ( .A(n_122), .B(n_277), .Y(n_305) );
OR2x2_ASAP7_75t_L g311 ( .A(n_122), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_122), .B(n_266), .Y(n_336) );
OR2x2_ASAP7_75t_L g354 ( .A(n_122), .B(n_173), .Y(n_354) );
BUFx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g218 ( .A(n_123), .B(n_149), .Y(n_218) );
INVx2_ASAP7_75t_L g240 ( .A(n_123), .Y(n_240) );
OR2x2_ASAP7_75t_L g262 ( .A(n_123), .B(n_149), .Y(n_262) );
AND2x2_ASAP7_75t_L g267 ( .A(n_123), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_123), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g323 ( .A(n_123), .B(n_217), .Y(n_323) );
BUFx2_ASAP7_75t_L g179 ( .A(n_125), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_128), .B(n_129), .C(n_134), .Y(n_126) );
O2A1O1Ixp33_ASAP7_75t_SL g140 ( .A1(n_128), .A2(n_134), .B(n_141), .C(n_142), .Y(n_140) );
O2A1O1Ixp33_ASAP7_75t_SL g151 ( .A1(n_128), .A2(n_134), .B(n_152), .C(n_153), .Y(n_151) );
O2A1O1Ixp33_ASAP7_75t_L g164 ( .A1(n_128), .A2(n_134), .B(n_165), .C(n_166), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_SL g180 ( .A1(n_128), .A2(n_134), .B(n_181), .C(n_182), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
INVx5_ASAP7_75t_L g185 ( .A(n_133), .Y(n_185) );
INVx1_ASAP7_75t_L g212 ( .A(n_134), .Y(n_212) );
INVx1_ASAP7_75t_SL g374 ( .A(n_136), .Y(n_374) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_149), .Y(n_136) );
INVx1_ASAP7_75t_SL g217 ( .A(n_137), .Y(n_217) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_137), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_137), .B(n_303), .Y(n_302) );
NAND3xp33_ASAP7_75t_L g369 ( .A(n_137), .B(n_240), .C(n_358), .Y(n_369) );
OA21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_139), .B(n_147), .Y(n_137) );
OA21x2_ASAP7_75t_L g149 ( .A1(n_138), .A2(n_150), .B(n_159), .Y(n_149) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_138), .A2(n_163), .B(n_171), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_145), .B(n_156), .Y(n_155) );
OAI22xp33_ASAP7_75t_L g183 ( .A1(n_145), .A2(n_184), .B1(n_185), .B2(n_186), .Y(n_183) );
INVx2_ASAP7_75t_L g268 ( .A(n_149), .Y(n_268) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_149), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_154), .B(n_168), .Y(n_167) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_161), .B(n_172), .Y(n_160) );
INVx1_ASAP7_75t_L g304 ( .A(n_161), .Y(n_304) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g222 ( .A(n_162), .B(n_204), .Y(n_222) );
INVx2_ASAP7_75t_L g239 ( .A(n_162), .Y(n_239) );
AND2x2_ASAP7_75t_L g244 ( .A(n_162), .B(n_205), .Y(n_244) );
AND2x2_ASAP7_75t_L g259 ( .A(n_162), .B(n_192), .Y(n_259) );
AND2x2_ASAP7_75t_L g271 ( .A(n_162), .B(n_243), .Y(n_271) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_172), .B(n_287), .Y(n_286) );
NAND2x1p5_ASAP7_75t_L g343 ( .A(n_172), .B(n_244), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_172), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_172), .B(n_238), .Y(n_366) );
BUFx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
OR2x2_ASAP7_75t_L g203 ( .A(n_173), .B(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_173), .B(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g248 ( .A(n_173), .B(n_192), .Y(n_248) );
AND2x2_ASAP7_75t_L g274 ( .A(n_173), .B(n_204), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_173), .B(n_314), .Y(n_313) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_178), .B(n_188), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AO21x2_ASAP7_75t_L g232 ( .A1(n_175), .A2(n_233), .B(n_234), .Y(n_232) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g233 ( .A(n_178), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_183), .B(n_187), .Y(n_182) );
O2A1O1Ixp33_ASAP7_75t_L g196 ( .A1(n_185), .A2(n_197), .B(n_198), .C(n_199), .Y(n_196) );
INVx2_ASAP7_75t_L g199 ( .A(n_187), .Y(n_199) );
INVx1_ASAP7_75t_L g234 ( .A(n_188), .Y(n_234) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_190), .B(n_214), .Y(n_213) );
OR2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_203), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_192), .B(n_225), .Y(n_224) );
AND2x4_ASAP7_75t_L g238 ( .A(n_192), .B(n_239), .Y(n_238) );
INVx3_ASAP7_75t_SL g243 ( .A(n_192), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_192), .B(n_230), .Y(n_296) );
OR2x2_ASAP7_75t_L g306 ( .A(n_192), .B(n_232), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_192), .B(n_274), .Y(n_334) );
OR2x2_ASAP7_75t_L g364 ( .A(n_192), .B(n_204), .Y(n_364) );
AND2x2_ASAP7_75t_L g368 ( .A(n_192), .B(n_205), .Y(n_368) );
NAND2xp5_ASAP7_75t_SL g381 ( .A(n_192), .B(n_244), .Y(n_381) );
AND2x2_ASAP7_75t_L g388 ( .A(n_192), .B(n_270), .Y(n_388) );
OR2x6_ASAP7_75t_L g192 ( .A(n_193), .B(n_201), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_199), .B(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_200), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_SL g331 ( .A(n_203), .Y(n_331) );
AND2x2_ASAP7_75t_L g270 ( .A(n_204), .B(n_232), .Y(n_270) );
AND2x2_ASAP7_75t_L g284 ( .A(n_204), .B(n_239), .Y(n_284) );
AND2x2_ASAP7_75t_L g287 ( .A(n_204), .B(n_243), .Y(n_287) );
INVx1_ASAP7_75t_L g314 ( .A(n_204), .Y(n_314) );
INVx2_ASAP7_75t_SL g204 ( .A(n_205), .Y(n_204) );
BUFx2_ASAP7_75t_L g226 ( .A(n_205), .Y(n_226) );
OAI322xp33_ASAP7_75t_L g517 ( .A1(n_210), .A2(n_518), .A3(n_519), .B1(n_523), .B2(n_524), .C1(n_527), .C2(n_529), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_218), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g385 ( .A1(n_216), .A2(n_262), .B(n_386), .C(n_387), .Y(n_385) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g292 ( .A(n_217), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_218), .B(n_235), .Y(n_250) );
AND2x2_ASAP7_75t_L g276 ( .A(n_218), .B(n_277), .Y(n_276) );
OAI21xp5_ASAP7_75t_SL g219 ( .A1(n_220), .A2(n_223), .B(n_227), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_221), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g247 ( .A(n_222), .B(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_222), .B(n_243), .Y(n_288) );
AND2x2_ASAP7_75t_L g379 ( .A(n_222), .B(n_230), .Y(n_379) );
INVxp67_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g252 ( .A(n_226), .B(n_239), .Y(n_252) );
OR2x2_ASAP7_75t_L g253 ( .A(n_226), .B(n_237), .Y(n_253) );
OAI322xp33_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_236), .A3(n_237), .B1(n_240), .B2(n_241), .C1(n_245), .C2(n_246), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_235), .Y(n_229) );
AND2x2_ASAP7_75t_L g340 ( .A(n_230), .B(n_252), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_230), .B(n_304), .Y(n_386) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_SL g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g283 ( .A(n_232), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g349 ( .A(n_236), .B(n_262), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_237), .B(n_331), .Y(n_330) );
INVx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_238), .B(n_270), .Y(n_327) );
AND2x2_ASAP7_75t_L g273 ( .A(n_239), .B(n_243), .Y(n_273) );
AND2x2_ASAP7_75t_L g281 ( .A(n_240), .B(n_282), .Y(n_281) );
A2O1A1Ixp33_ASAP7_75t_L g378 ( .A1(n_240), .A2(n_319), .B(n_379), .C(n_380), .Y(n_378) );
AOI21xp33_ASAP7_75t_L g351 ( .A1(n_241), .A2(n_254), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_SL g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_243), .B(n_270), .Y(n_310) );
AND2x2_ASAP7_75t_L g316 ( .A(n_243), .B(n_284), .Y(n_316) );
AND2x2_ASAP7_75t_L g350 ( .A(n_243), .B(n_252), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_244), .B(n_259), .Y(n_258) );
INVx2_ASAP7_75t_SL g360 ( .A(n_244), .Y(n_360) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g275 ( .A1(n_248), .A2(n_276), .B1(n_278), .B2(n_283), .Y(n_275) );
OAI22xp5_ASAP7_75t_SL g249 ( .A1(n_250), .A2(n_251), .B1(n_253), .B2(n_254), .Y(n_249) );
OAI22xp33_ASAP7_75t_L g285 ( .A1(n_250), .A2(n_286), .B1(n_288), .B2(n_289), .Y(n_285) );
INVxp67_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
AOI221xp5_ASAP7_75t_L g356 ( .A1(n_255), .A2(n_357), .B1(n_359), .B2(n_361), .C(n_365), .Y(n_356) );
AOI211xp5_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_260), .B(n_264), .C(n_285), .Y(n_256) );
INVxp67_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
OR2x2_ASAP7_75t_L g326 ( .A(n_262), .B(n_279), .Y(n_326) );
INVx1_ASAP7_75t_L g377 ( .A(n_262), .Y(n_377) );
OAI221xp5_ASAP7_75t_L g264 ( .A1(n_263), .A2(n_265), .B1(n_269), .B2(n_272), .C(n_275), .Y(n_264) );
INVx2_ASAP7_75t_SL g319 ( .A(n_263), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx1_ASAP7_75t_L g384 ( .A(n_266), .Y(n_384) );
AND2x2_ASAP7_75t_L g308 ( .A(n_267), .B(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g293 ( .A(n_268), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx1_ASAP7_75t_L g355 ( .A(n_271), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_279), .B(n_381), .Y(n_380) );
CKINVDCx16_ASAP7_75t_R g279 ( .A(n_280), .Y(n_279) );
INVxp67_ASAP7_75t_L g324 ( .A(n_282), .Y(n_324) );
O2A1O1Ixp33_ASAP7_75t_L g294 ( .A1(n_283), .A2(n_295), .B(n_297), .C(n_299), .Y(n_294) );
INVx1_ASAP7_75t_L g372 ( .A(n_286), .Y(n_372) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_290), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx2_ASAP7_75t_L g303 ( .A(n_293), .Y(n_303) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OAI222xp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_306), .B1(n_307), .B2(n_310), .C1(n_311), .C2(n_313), .Y(n_299) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_SL g339 ( .A(n_303), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_306), .B(n_360), .Y(n_359) );
NAND2xp33_ASAP7_75t_SL g337 ( .A(n_307), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_SL g312 ( .A(n_309), .Y(n_312) );
AND2x2_ASAP7_75t_L g376 ( .A(n_309), .B(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g342 ( .A(n_312), .B(n_339), .Y(n_342) );
INVx1_ASAP7_75t_L g371 ( .A(n_313), .Y(n_371) );
AOI211xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B(n_320), .C(n_325), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_319), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
AOI322xp5_ASAP7_75t_L g370 ( .A1(n_322), .A2(n_350), .A3(n_355), .B1(n_371), .B2(n_372), .C1(n_373), .C2(n_376), .Y(n_370) );
AND2x2_ASAP7_75t_L g357 ( .A(n_323), .B(n_358), .Y(n_357) );
OAI22xp33_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_327), .B1(n_328), .B2(n_330), .Y(n_325) );
INVxp33_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AOI221xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .B1(n_337), .B2(n_340), .C(n_341), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
NAND5xp2_ASAP7_75t_L g344 ( .A(n_345), .B(n_356), .C(n_370), .D(n_378), .E(n_382), .Y(n_344) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_350), .B(n_351), .Y(n_345) );
INVxp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVxp33_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
A2O1A1Ixp33_ASAP7_75t_L g382 ( .A1(n_358), .A2(n_383), .B(n_384), .C(n_385), .Y(n_382) );
AOI31xp33_ASAP7_75t_L g365 ( .A1(n_360), .A2(n_366), .A3(n_367), .B(n_369), .Y(n_365) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_L g383 ( .A(n_381), .Y(n_383) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g389 ( .A(n_390), .Y(n_389) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_391), .A2(n_513), .B(n_526), .Y(n_525) );
XNOR2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_403), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B1(n_399), .B2(n_402), .Y(n_394) );
CKINVDCx20_ASAP7_75t_R g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g402 ( .A(n_399), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B1(n_406), .B2(n_504), .Y(n_403) );
CKINVDCx20_ASAP7_75t_R g404 ( .A(n_405), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_406), .Y(n_504) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_SL g407 ( .A(n_408), .B(n_463), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_409), .B(n_442), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_433), .Y(n_409) );
BUFx3_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_423), .Y(n_413) );
AND2x6_ASAP7_75t_L g430 ( .A(n_414), .B(n_431), .Y(n_430) );
AND2x4_ASAP7_75t_L g446 ( .A(n_414), .B(n_447), .Y(n_446) );
AND2x6_ASAP7_75t_L g481 ( .A(n_414), .B(n_476), .Y(n_481) );
AND2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_420), .Y(n_414) );
AND2x2_ASAP7_75t_L g437 ( .A(n_415), .B(n_421), .Y(n_437) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_416), .B(n_421), .Y(n_441) );
AND2x2_ASAP7_75t_L g452 ( .A(n_416), .B(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g469 ( .A(n_416), .B(n_425), .Y(n_469) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g422 ( .A(n_419), .Y(n_422) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g453 ( .A(n_421), .Y(n_453) );
INVx1_ASAP7_75t_L g487 ( .A(n_421), .Y(n_487) );
AND2x4_ASAP7_75t_L g436 ( .A(n_423), .B(n_437), .Y(n_436) );
AND2x4_ASAP7_75t_L g439 ( .A(n_423), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g451 ( .A(n_423), .B(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_426), .Y(n_423) );
OR2x2_ASAP7_75t_L g432 ( .A(n_424), .B(n_427), .Y(n_432) );
AND2x2_ASAP7_75t_L g447 ( .A(n_424), .B(n_427), .Y(n_447) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g476 ( .A(n_425), .B(n_427), .Y(n_476) );
INVx1_ASAP7_75t_L g470 ( .A(n_426), .Y(n_470) );
AND2x2_ASAP7_75t_L g486 ( .A(n_426), .B(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g462 ( .A(n_427), .Y(n_462) );
INVx4_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx11_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g498 ( .A(n_432), .B(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx3_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g499 ( .A(n_437), .Y(n_499) );
NAND2x1p5_ASAP7_75t_L g503 ( .A(n_437), .B(n_447), .Y(n_503) );
BUFx3_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OR2x6_ASAP7_75t_L g461 ( .A(n_441), .B(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_454), .Y(n_442) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx6_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g458 ( .A(n_447), .B(n_452), .Y(n_458) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
BUFx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g478 ( .A(n_453), .Y(n_478) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx4_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx8_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx4f_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
INVx6_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
NOR3xp33_ASAP7_75t_SL g463 ( .A(n_464), .B(n_479), .C(n_494), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B1(n_471), .B2(n_472), .Y(n_464) );
INVx3_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
INVx4_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NAND2x1p5_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
AND2x4_ASAP7_75t_L g485 ( .A(n_469), .B(n_486), .Y(n_485) );
AND2x4_ASAP7_75t_L g492 ( .A(n_469), .B(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g473 ( .A(n_474), .Y(n_473) );
OR2x6_ASAP7_75t_L g474 ( .A(n_475), .B(n_477), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
OAI221xp5_ASAP7_75t_SL g479 ( .A1(n_480), .A2(n_482), .B1(n_483), .B2(n_488), .C(n_489), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g493 ( .A(n_487), .Y(n_493) );
BUFx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B1(n_500), .B2(n_501), .Y(n_494) );
INVx1_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
AND3x1_ASAP7_75t_SL g507 ( .A(n_508), .B(n_513), .C(n_515), .Y(n_507) );
INVxp67_ASAP7_75t_L g522 ( .A(n_508), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
CKINVDCx16_ASAP7_75t_R g523 ( .A(n_513), .Y(n_523) );
INVx1_ASAP7_75t_L g532 ( .A(n_513), .Y(n_532) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_514), .B(n_516), .Y(n_526) );
OR2x2_ASAP7_75t_SL g531 ( .A(n_515), .B(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_520), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_530), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_531), .Y(n_530) );
endmodule