module fake_aes_9025_n_16 (n_3, n_1, n_2, n_0, n_16);
input n_3;
input n_1;
input n_2;
input n_0;
output n_16;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
CKINVDCx20_ASAP7_75t_R g4 ( .A(n_0), .Y(n_4) );
CKINVDCx5p33_ASAP7_75t_R g5 ( .A(n_2), .Y(n_5) );
INVx2_ASAP7_75t_L g6 ( .A(n_1), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_6), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_7), .B(n_5), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
INVx2_ASAP7_75t_SL g10 ( .A(n_8), .Y(n_10) );
INVxp67_ASAP7_75t_SL g11 ( .A(n_10), .Y(n_11) );
AOI22xp5_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_10), .B1(n_9), .B2(n_4), .Y(n_12) );
INVx2_ASAP7_75t_SL g13 ( .A(n_12), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_13), .Y(n_14) );
BUFx6f_ASAP7_75t_L g15 ( .A(n_13), .Y(n_15) );
AOI22xp33_ASAP7_75t_SL g16 ( .A1(n_15), .A2(n_3), .B1(n_14), .B2(n_13), .Y(n_16) );
endmodule