module real_aes_10337_n_14 (n_13, n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_12, n_1, n_10, n_11, n_14);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_10;
input n_11;
output n_14;
wire n_28;
wire n_17;
wire n_22;
wire n_24;
wire n_41;
wire n_34;
wire n_19;
wire n_40;
wire n_46;
wire n_25;
wire n_43;
wire n_32;
wire n_30;
wire n_16;
wire n_37;
wire n_35;
wire n_42;
wire n_45;
wire n_39;
wire n_15;
wire n_27;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_44;
wire n_26;
wire n_18;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_0), .Y(n_23) );
NOR4xp25_ASAP7_75t_SL g34 ( .A(n_0), .B(n_27), .C(n_35), .D(n_36), .Y(n_34) );
NOR3xp33_ASAP7_75t_SL g20 ( .A(n_1), .B(n_11), .C(n_21), .Y(n_20) );
NOR3xp33_ASAP7_75t_SL g25 ( .A(n_1), .B(n_7), .C(n_26), .Y(n_25) );
NOR2xp33_ASAP7_75t_R g22 ( .A(n_2), .B(n_5), .Y(n_22) );
NAND2xp33_ASAP7_75t_R g26 ( .A(n_3), .B(n_22), .Y(n_26) );
CKINVDCx5p33_ASAP7_75t_R g27 ( .A(n_4), .Y(n_27) );
CKINVDCx5p33_ASAP7_75t_R g29 ( .A(n_6), .Y(n_29) );
NOR2xp33_ASAP7_75t_R g33 ( .A(n_6), .B(n_12), .Y(n_33) );
NOR2xp33_ASAP7_75t_R g39 ( .A(n_6), .B(n_28), .Y(n_39) );
NAND2xp33_ASAP7_75t_SL g43 ( .A(n_6), .B(n_28), .Y(n_43) );
NAND2xp33_ASAP7_75t_R g46 ( .A(n_6), .B(n_12), .Y(n_46) );
AOI22xp33_ASAP7_75t_SL g30 ( .A1(n_8), .A2(n_9), .B1(n_31), .B2(n_37), .Y(n_30) );
AOI22xp33_ASAP7_75t_L g40 ( .A1(n_10), .A2(n_13), .B1(n_41), .B2(n_45), .Y(n_40) );
CKINVDCx5p33_ASAP7_75t_R g36 ( .A(n_11), .Y(n_36) );
CKINVDCx5p33_ASAP7_75t_R g28 ( .A(n_12), .Y(n_28) );
NAND3xp33_ASAP7_75t_L g14 ( .A(n_15), .B(n_30), .C(n_40), .Y(n_14) );
NAND2xp33_ASAP7_75t_R g15 ( .A(n_16), .B(n_29), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_17), .Y(n_16) );
NAND2xp33_ASAP7_75t_R g17 ( .A(n_18), .B(n_28), .Y(n_17) );
NOR2xp33_ASAP7_75t_R g18 ( .A(n_19), .B(n_24), .Y(n_18) );
NAND2xp33_ASAP7_75t_R g19 ( .A(n_20), .B(n_23), .Y(n_19) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_22), .Y(n_21) );
NAND2xp33_ASAP7_75t_R g24 ( .A(n_25), .B(n_27), .Y(n_24) );
CKINVDCx5p33_ASAP7_75t_R g35 ( .A(n_25), .Y(n_35) );
CKINVDCx5p33_ASAP7_75t_R g31 ( .A(n_32), .Y(n_31) );
NAND2xp33_ASAP7_75t_R g32 ( .A(n_33), .B(n_34), .Y(n_32) );
NAND2xp33_ASAP7_75t_R g38 ( .A(n_34), .B(n_39), .Y(n_38) );
CKINVDCx5p33_ASAP7_75t_R g44 ( .A(n_34), .Y(n_44) );
CKINVDCx5p33_ASAP7_75t_R g37 ( .A(n_38), .Y(n_37) );
HB1xp67_ASAP7_75t_L g41 ( .A(n_42), .Y(n_41) );
NOR2xp33_ASAP7_75t_R g42 ( .A(n_43), .B(n_44), .Y(n_42) );
NOR2xp33_ASAP7_75t_R g45 ( .A(n_44), .B(n_46), .Y(n_45) );
endmodule