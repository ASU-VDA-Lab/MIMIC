module real_aes_6502_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_725;
wire n_119;
wire n_504;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g468 ( .A1(n_0), .A2(n_148), .B(n_469), .C(n_472), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_1), .B(n_463), .Y(n_473) );
INVx1_ASAP7_75t_L g424 ( .A(n_2), .Y(n_424) );
INVx1_ASAP7_75t_L g146 ( .A(n_3), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_4), .B(n_149), .Y(n_453) );
AOI222xp33_ASAP7_75t_L g432 ( .A1(n_5), .A2(n_433), .B1(n_719), .B2(n_720), .C1(n_726), .C2(n_727), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_6), .A2(n_458), .B(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_7), .B(n_430), .Y(n_429) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_8), .A2(n_171), .B(n_539), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_9), .A2(n_41), .B1(n_136), .B2(n_194), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_10), .A2(n_11), .B1(n_723), .B2(n_724), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_10), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_11), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_12), .B(n_171), .Y(n_179) );
AND2x6_ASAP7_75t_L g151 ( .A(n_13), .B(n_152), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_14), .A2(n_151), .B(n_449), .C(n_513), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_15), .B(n_42), .Y(n_425) );
INVx1_ASAP7_75t_L g736 ( .A(n_15), .Y(n_736) );
INVx1_ASAP7_75t_L g130 ( .A(n_16), .Y(n_130) );
INVx1_ASAP7_75t_L g127 ( .A(n_17), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_18), .B(n_132), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_19), .B(n_149), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_20), .B(n_123), .Y(n_181) );
AO32x2_ASAP7_75t_L g232 ( .A1(n_21), .A2(n_122), .A3(n_165), .B1(n_171), .B2(n_233), .Y(n_232) );
OAI22xp5_ASAP7_75t_SL g111 ( .A1(n_22), .A2(n_33), .B1(n_112), .B2(n_113), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_22), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_23), .B(n_136), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_24), .B(n_123), .Y(n_153) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_25), .A2(n_56), .B1(n_136), .B2(n_194), .Y(n_235) );
AOI22xp33_ASAP7_75t_SL g196 ( .A1(n_26), .A2(n_83), .B1(n_132), .B2(n_136), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_27), .B(n_136), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_28), .A2(n_165), .B(n_449), .C(n_480), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_29), .A2(n_165), .B(n_449), .C(n_542), .Y(n_541) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_30), .Y(n_141) );
OAI22xp5_ASAP7_75t_SL g720 ( .A1(n_31), .A2(n_721), .B1(n_722), .B2(n_725), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_31), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_32), .B(n_167), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_33), .Y(n_113) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_33), .A2(n_113), .B1(n_114), .B2(n_115), .Y(n_437) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_34), .A2(n_458), .B(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_35), .B(n_167), .Y(n_209) );
INVx2_ASAP7_75t_L g134 ( .A(n_36), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_37), .A2(n_455), .B(n_498), .C(n_499), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_38), .B(n_136), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_39), .B(n_167), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_40), .B(n_216), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_42), .B(n_736), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_43), .B(n_478), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_44), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_45), .B(n_149), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_46), .B(n_458), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_47), .A2(n_455), .B(n_498), .C(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_48), .B(n_136), .Y(n_174) );
INVx1_ASAP7_75t_L g470 ( .A(n_49), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_50), .A2(n_91), .B1(n_194), .B2(n_195), .Y(n_193) );
INVx1_ASAP7_75t_L g523 ( .A(n_51), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_52), .B(n_136), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_53), .B(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_54), .B(n_458), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_55), .B(n_144), .Y(n_178) );
AOI22xp33_ASAP7_75t_SL g185 ( .A1(n_57), .A2(n_61), .B1(n_132), .B2(n_136), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_58), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_59), .B(n_136), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_60), .B(n_136), .Y(n_213) );
INVx1_ASAP7_75t_L g152 ( .A(n_62), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_63), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_64), .B(n_463), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_65), .A2(n_138), .B(n_144), .C(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_66), .B(n_136), .Y(n_147) );
INVx1_ASAP7_75t_L g126 ( .A(n_67), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_68), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_69), .B(n_149), .Y(n_501) );
AO32x2_ASAP7_75t_L g191 ( .A1(n_70), .A2(n_165), .A3(n_171), .B1(n_192), .B2(n_197), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_71), .B(n_150), .Y(n_514) );
INVx1_ASAP7_75t_L g161 ( .A(n_72), .Y(n_161) );
INVx1_ASAP7_75t_L g204 ( .A(n_73), .Y(n_204) );
CKINVDCx16_ASAP7_75t_R g466 ( .A(n_74), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_75), .B(n_482), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_76), .A2(n_449), .B(n_451), .C(n_455), .Y(n_448) );
OAI321xp33_ASAP7_75t_L g108 ( .A1(n_77), .A2(n_109), .A3(n_419), .B1(n_426), .B2(n_427), .C(n_429), .Y(n_108) );
INVx1_ASAP7_75t_L g426 ( .A(n_77), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_78), .B(n_132), .Y(n_205) );
CKINVDCx16_ASAP7_75t_R g532 ( .A(n_79), .Y(n_532) );
INVx1_ASAP7_75t_L g740 ( .A(n_80), .Y(n_740) );
AOI22xp33_ASAP7_75t_SL g104 ( .A1(n_81), .A2(n_105), .B1(n_733), .B2(n_741), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_82), .B(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_84), .B(n_194), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_85), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_86), .B(n_132), .Y(n_208) );
INVx2_ASAP7_75t_L g124 ( .A(n_87), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_88), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_89), .B(n_164), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_90), .B(n_132), .Y(n_175) );
OR2x2_ASAP7_75t_L g421 ( .A(n_92), .B(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g436 ( .A(n_92), .B(n_423), .Y(n_436) );
INVx2_ASAP7_75t_L g440 ( .A(n_92), .Y(n_440) );
NAND3xp33_ASAP7_75t_SL g737 ( .A(n_92), .B(n_424), .C(n_738), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g184 ( .A1(n_93), .A2(n_103), .B1(n_132), .B2(n_133), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_94), .B(n_458), .Y(n_496) );
INVx1_ASAP7_75t_L g500 ( .A(n_95), .Y(n_500) );
INVxp67_ASAP7_75t_L g535 ( .A(n_96), .Y(n_535) );
XNOR2xp5_ASAP7_75t_L g109 ( .A(n_97), .B(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_98), .B(n_132), .Y(n_159) );
INVx1_ASAP7_75t_L g452 ( .A(n_99), .Y(n_452) );
INVx1_ASAP7_75t_L g510 ( .A(n_100), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_101), .B(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g525 ( .A(n_102), .B(n_167), .Y(n_525) );
OA21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_108), .B(n_431), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g732 ( .A(n_107), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_109), .B(n_428), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_114), .B1(n_115), .B2(n_418), .Y(n_110) );
INVx1_ASAP7_75t_L g418 ( .A(n_111), .Y(n_418) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OR5x1_ASAP7_75t_L g115 ( .A(n_116), .B(n_309), .C(n_367), .D(n_403), .E(n_410), .Y(n_115) );
NAND3xp33_ASAP7_75t_SL g116 ( .A(n_117), .B(n_255), .C(n_279), .Y(n_116) );
AOI221xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_187), .B1(n_221), .B2(n_226), .C(n_236), .Y(n_117) );
OAI21xp5_ASAP7_75t_SL g389 ( .A1(n_118), .A2(n_390), .B(n_392), .Y(n_389) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_168), .Y(n_118) );
NAND2x1p5_ASAP7_75t_L g379 ( .A(n_119), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_154), .Y(n_119) );
INVx2_ASAP7_75t_L g225 ( .A(n_120), .Y(n_225) );
AND2x2_ASAP7_75t_L g238 ( .A(n_120), .B(n_170), .Y(n_238) );
AND2x2_ASAP7_75t_L g292 ( .A(n_120), .B(n_169), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_120), .B(n_155), .Y(n_307) );
OA21x2_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_128), .B(n_153), .Y(n_120) );
OA21x2_ASAP7_75t_L g155 ( .A1(n_121), .A2(n_156), .B(n_166), .Y(n_155) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_122), .B(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_123), .Y(n_171) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_124), .B(n_125), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
OAI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_142), .B(n_151), .Y(n_128) );
O2A1O1Ixp33_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_131), .B(n_135), .C(n_138), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_131), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_131), .A2(n_543), .B(n_544), .Y(n_542) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g137 ( .A(n_134), .Y(n_137) );
INVx1_ASAP7_75t_L g145 ( .A(n_134), .Y(n_145) );
INVx3_ASAP7_75t_L g203 ( .A(n_136), .Y(n_203) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_136), .Y(n_454) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g194 ( .A(n_137), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_137), .Y(n_195) );
AND2x6_ASAP7_75t_L g449 ( .A(n_137), .B(n_450), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_L g451 ( .A1(n_138), .A2(n_452), .B(n_453), .C(n_454), .Y(n_451) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_139), .A2(n_207), .B(n_208), .Y(n_206) );
INVx4_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g482 ( .A(n_140), .Y(n_482) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx3_ASAP7_75t_L g150 ( .A(n_141), .Y(n_150) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_141), .Y(n_164) );
INVx1_ASAP7_75t_L g216 ( .A(n_141), .Y(n_216) );
INVx1_ASAP7_75t_L g450 ( .A(n_141), .Y(n_450) );
AND2x2_ASAP7_75t_L g459 ( .A(n_141), .B(n_145), .Y(n_459) );
O2A1O1Ixp33_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_146), .B(n_147), .C(n_148), .Y(n_142) );
O2A1O1Ixp5_ASAP7_75t_L g160 ( .A1(n_143), .A2(n_161), .B(n_162), .C(n_163), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_143), .A2(n_481), .B(n_483), .Y(n_480) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_148), .A2(n_177), .B(n_178), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g183 ( .A1(n_148), .A2(n_164), .B1(n_184), .B2(n_185), .Y(n_183) );
OAI22xp5_ASAP7_75t_L g233 ( .A1(n_148), .A2(n_164), .B1(n_234), .B2(n_235), .Y(n_233) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_149), .A2(n_158), .B(n_159), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_149), .A2(n_174), .B(n_175), .Y(n_173) );
O2A1O1Ixp5_ASAP7_75t_SL g202 ( .A1(n_149), .A2(n_203), .B(n_204), .C(n_205), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_149), .B(n_535), .Y(n_534) );
INVx5_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OAI22xp5_ASAP7_75t_SL g192 ( .A1(n_150), .A2(n_164), .B1(n_193), .B2(n_196), .Y(n_192) );
BUFx3_ASAP7_75t_L g165 ( .A(n_151), .Y(n_165) );
OAI21xp5_ASAP7_75t_L g172 ( .A1(n_151), .A2(n_173), .B(n_176), .Y(n_172) );
OAI21xp5_ASAP7_75t_L g201 ( .A1(n_151), .A2(n_202), .B(n_206), .Y(n_201) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_151), .A2(n_212), .B(n_217), .Y(n_211) );
INVx4_ASAP7_75t_SL g456 ( .A(n_151), .Y(n_456) );
AND2x4_ASAP7_75t_L g458 ( .A(n_151), .B(n_459), .Y(n_458) );
NAND2x1p5_ASAP7_75t_L g511 ( .A(n_151), .B(n_459), .Y(n_511) );
AND2x2_ASAP7_75t_L g325 ( .A(n_154), .B(n_266), .Y(n_325) );
AND2x2_ASAP7_75t_L g358 ( .A(n_154), .B(n_170), .Y(n_358) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
OR2x2_ASAP7_75t_L g265 ( .A(n_155), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g278 ( .A(n_155), .B(n_170), .Y(n_278) );
AND2x2_ASAP7_75t_L g285 ( .A(n_155), .B(n_266), .Y(n_285) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_155), .Y(n_294) );
AND2x2_ASAP7_75t_L g301 ( .A(n_155), .B(n_169), .Y(n_301) );
INVx1_ASAP7_75t_L g332 ( .A(n_155), .Y(n_332) );
OAI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_160), .B(n_165), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_163), .A2(n_218), .B(n_219), .Y(n_217) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx4_ASAP7_75t_L g471 ( .A(n_164), .Y(n_471) );
NAND3xp33_ASAP7_75t_L g182 ( .A(n_165), .B(n_183), .C(n_186), .Y(n_182) );
INVx2_ASAP7_75t_L g197 ( .A(n_167), .Y(n_197) );
OA21x2_ASAP7_75t_L g200 ( .A1(n_167), .A2(n_201), .B(n_209), .Y(n_200) );
OA21x2_ASAP7_75t_L g210 ( .A1(n_167), .A2(n_211), .B(n_220), .Y(n_210) );
INVx1_ASAP7_75t_L g488 ( .A(n_167), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_167), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_167), .A2(n_520), .B(n_521), .Y(n_519) );
INVx1_ASAP7_75t_L g308 ( .A(n_168), .Y(n_308) );
AND2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_180), .Y(n_168) );
INVx2_ASAP7_75t_L g264 ( .A(n_169), .Y(n_264) );
AND2x2_ASAP7_75t_L g286 ( .A(n_169), .B(n_225), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_169), .B(n_332), .Y(n_337) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_170), .B(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g409 ( .A(n_170), .B(n_373), .Y(n_409) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_179), .Y(n_170) );
INVx4_ASAP7_75t_L g186 ( .A(n_171), .Y(n_186) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_171), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_171), .A2(n_540), .B(n_541), .Y(n_539) );
INVx2_ASAP7_75t_L g223 ( .A(n_180), .Y(n_223) );
INVx3_ASAP7_75t_L g324 ( .A(n_180), .Y(n_324) );
OR2x2_ASAP7_75t_L g354 ( .A(n_180), .B(n_355), .Y(n_354) );
NOR2x1_ASAP7_75t_L g380 ( .A(n_180), .B(n_264), .Y(n_380) );
AND2x4_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
INVx1_ASAP7_75t_L g267 ( .A(n_181), .Y(n_267) );
AO21x1_ASAP7_75t_L g266 ( .A1(n_183), .A2(n_186), .B(n_267), .Y(n_266) );
AO21x2_ASAP7_75t_L g446 ( .A1(n_186), .A2(n_447), .B(n_460), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_186), .B(n_461), .Y(n_460) );
INVx3_ASAP7_75t_L g463 ( .A(n_186), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_186), .B(n_504), .Y(n_503) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_186), .A2(n_509), .B(n_516), .Y(n_508) );
AOI33xp33_ASAP7_75t_L g400 ( .A1(n_187), .A2(n_238), .A3(n_252), .B1(n_324), .B2(n_401), .B3(n_402), .Y(n_400) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
OR2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_198), .Y(n_188) );
OR2x2_ASAP7_75t_L g253 ( .A(n_189), .B(n_254), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_189), .B(n_250), .Y(n_312) );
OR2x2_ASAP7_75t_L g365 ( .A(n_189), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g291 ( .A(n_190), .B(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g316 ( .A(n_190), .B(n_198), .Y(n_316) );
AND2x2_ASAP7_75t_L g383 ( .A(n_190), .B(n_228), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_190), .A2(n_283), .B(n_409), .Y(n_408) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g230 ( .A(n_191), .Y(n_230) );
INVx1_ASAP7_75t_L g243 ( .A(n_191), .Y(n_243) );
AND2x2_ASAP7_75t_L g262 ( .A(n_191), .B(n_232), .Y(n_262) );
AND2x2_ASAP7_75t_L g311 ( .A(n_191), .B(n_231), .Y(n_311) );
INVx2_ASAP7_75t_L g472 ( .A(n_195), .Y(n_472) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_195), .Y(n_502) );
INVx1_ASAP7_75t_L g485 ( .A(n_197), .Y(n_485) );
INVx2_ASAP7_75t_SL g353 ( .A(n_198), .Y(n_353) );
OR2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_210), .Y(n_198) );
INVx2_ASAP7_75t_L g273 ( .A(n_199), .Y(n_273) );
INVx1_ASAP7_75t_L g404 ( .A(n_199), .Y(n_404) );
AND2x2_ASAP7_75t_L g417 ( .A(n_199), .B(n_298), .Y(n_417) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g244 ( .A(n_200), .Y(n_244) );
OR2x2_ASAP7_75t_L g250 ( .A(n_200), .B(n_251), .Y(n_250) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_200), .Y(n_261) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_210), .Y(n_228) );
AND2x2_ASAP7_75t_L g245 ( .A(n_210), .B(n_231), .Y(n_245) );
INVx1_ASAP7_75t_L g251 ( .A(n_210), .Y(n_251) );
INVx1_ASAP7_75t_L g258 ( .A(n_210), .Y(n_258) );
AND2x2_ASAP7_75t_L g283 ( .A(n_210), .B(n_232), .Y(n_283) );
INVx2_ASAP7_75t_L g299 ( .A(n_210), .Y(n_299) );
AND2x2_ASAP7_75t_L g392 ( .A(n_210), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_210), .B(n_273), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_215), .Y(n_212) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_SL g221 ( .A(n_222), .Y(n_221) );
OR2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
INVx2_ASAP7_75t_L g247 ( .A(n_223), .Y(n_247) );
INVx1_ASAP7_75t_L g276 ( .A(n_223), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_223), .B(n_307), .Y(n_373) );
INVx1_ASAP7_75t_SL g333 ( .A(n_224), .Y(n_333) );
INVx2_ASAP7_75t_L g254 ( .A(n_225), .Y(n_254) );
AND2x2_ASAP7_75t_L g323 ( .A(n_225), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g339 ( .A(n_225), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_229), .Y(n_226) );
INVx1_ASAP7_75t_L g401 ( .A(n_227), .Y(n_401) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g256 ( .A(n_229), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g359 ( .A(n_229), .B(n_349), .Y(n_359) );
AOI21xp5_ASAP7_75t_L g411 ( .A1(n_229), .A2(n_370), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
AND2x2_ASAP7_75t_L g272 ( .A(n_230), .B(n_273), .Y(n_272) );
BUFx2_ASAP7_75t_L g297 ( .A(n_230), .Y(n_297) );
INVx1_ASAP7_75t_L g321 ( .A(n_230), .Y(n_321) );
OR2x2_ASAP7_75t_L g385 ( .A(n_231), .B(n_244), .Y(n_385) );
NOR2xp67_ASAP7_75t_L g393 ( .A(n_231), .B(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g298 ( .A(n_232), .B(n_299), .Y(n_298) );
BUFx2_ASAP7_75t_L g305 ( .A(n_232), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_239), .B1(n_246), .B2(n_248), .Y(n_236) );
OR2x2_ASAP7_75t_L g315 ( .A(n_237), .B(n_265), .Y(n_315) );
INVx1_ASAP7_75t_SL g237 ( .A(n_238), .Y(n_237) );
AOI222xp33_ASAP7_75t_L g356 ( .A1(n_238), .A2(n_357), .B1(n_359), .B2(n_360), .C1(n_361), .C2(n_364), .Y(n_356) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_245), .Y(n_240) );
INVx1_ASAP7_75t_SL g241 ( .A(n_242), .Y(n_241) );
OR2x2_ASAP7_75t_L g303 ( .A(n_242), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
AND2x2_ASAP7_75t_SL g257 ( .A(n_244), .B(n_258), .Y(n_257) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_244), .Y(n_328) );
AND2x2_ASAP7_75t_L g376 ( .A(n_244), .B(n_245), .Y(n_376) );
INVx1_ASAP7_75t_L g394 ( .A(n_244), .Y(n_394) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g360 ( .A(n_247), .B(n_286), .Y(n_360) );
AND2x2_ASAP7_75t_L g402 ( .A(n_247), .B(n_278), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_252), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_249), .B(n_297), .Y(n_384) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_250), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g277 ( .A(n_254), .B(n_278), .Y(n_277) );
INVx3_ASAP7_75t_L g345 ( .A(n_254), .Y(n_345) );
O2A1O1Ixp33_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_259), .B(n_263), .C(n_268), .Y(n_255) );
INVxp67_ASAP7_75t_L g269 ( .A(n_256), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_257), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_257), .B(n_304), .Y(n_399) );
BUFx3_ASAP7_75t_L g363 ( .A(n_258), .Y(n_363) );
INVx1_ASAP7_75t_L g270 ( .A(n_259), .Y(n_270) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g289 ( .A(n_261), .B(n_283), .Y(n_289) );
INVx1_ASAP7_75t_SL g329 ( .A(n_262), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx1_ASAP7_75t_L g319 ( .A(n_264), .Y(n_319) );
AND2x2_ASAP7_75t_L g342 ( .A(n_264), .B(n_325), .Y(n_342) );
INVx1_ASAP7_75t_SL g313 ( .A(n_265), .Y(n_313) );
INVx1_ASAP7_75t_L g340 ( .A(n_266), .Y(n_340) );
AOI31xp33_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_270), .A3(n_271), .B(n_274), .Y(n_268) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g361 ( .A(n_272), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g335 ( .A(n_273), .Y(n_335) );
BUFx2_ASAP7_75t_L g349 ( .A(n_273), .Y(n_349) );
AND2x2_ASAP7_75t_L g377 ( .A(n_273), .B(n_298), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_SL g350 ( .A(n_277), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_278), .B(n_345), .Y(n_391) );
AND2x2_ASAP7_75t_L g398 ( .A(n_278), .B(n_324), .Y(n_398) );
AOI211xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_284), .B(n_287), .C(n_302), .Y(n_279) );
INVxp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AOI221xp5_ASAP7_75t_L g310 ( .A1(n_284), .A2(n_311), .B1(n_312), .B2(n_313), .C(n_314), .Y(n_310) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
AND2x2_ASAP7_75t_L g318 ( .A(n_285), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g355 ( .A(n_286), .Y(n_355) );
OAI32xp33_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_290), .A3(n_293), .B1(n_295), .B2(n_300), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
O2A1O1Ixp33_ASAP7_75t_L g341 ( .A1(n_289), .A2(n_342), .B(n_343), .C(n_346), .Y(n_341) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
OAI21xp5_ASAP7_75t_SL g405 ( .A1(n_297), .A2(n_406), .B(n_407), .Y(n_405) );
INVx1_ASAP7_75t_L g366 ( .A(n_298), .Y(n_366) );
INVxp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_303), .B(n_306), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_304), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g352 ( .A(n_304), .B(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g369 ( .A(n_306), .Y(n_369) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
NAND4xp25_ASAP7_75t_SL g309 ( .A(n_310), .B(n_322), .C(n_341), .D(n_356), .Y(n_309) );
AND2x2_ASAP7_75t_L g348 ( .A(n_311), .B(n_349), .Y(n_348) );
AND2x4_ASAP7_75t_L g370 ( .A(n_311), .B(n_363), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_313), .B(n_345), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_316), .B1(n_317), .B2(n_320), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_315), .A2(n_366), .B1(n_397), .B2(n_399), .Y(n_396) );
O2A1O1Ixp33_ASAP7_75t_L g403 ( .A1(n_315), .A2(n_404), .B(n_405), .C(n_408), .Y(n_403) );
INVx2_ASAP7_75t_L g374 ( .A(n_316), .Y(n_374) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AOI222xp33_ASAP7_75t_L g368 ( .A1(n_318), .A2(n_352), .B1(n_369), .B2(n_370), .C1(n_371), .C2(n_374), .Y(n_368) );
O2A1O1Ixp33_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_325), .B(n_326), .C(n_330), .Y(n_322) );
INVx1_ASAP7_75t_L g388 ( .A(n_323), .Y(n_388) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OAI22xp33_ASAP7_75t_L g330 ( .A1(n_327), .A2(n_331), .B1(n_334), .B2(n_336), .Y(n_330) );
OR2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
OR2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g357 ( .A(n_339), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g415 ( .A(n_342), .Y(n_415) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OAI22xp33_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_350), .B1(n_351), .B2(n_354), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_349), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g406 ( .A(n_354), .Y(n_406) );
INVx1_ASAP7_75t_L g387 ( .A(n_358), .Y(n_387) );
CKINVDCx16_ASAP7_75t_R g414 ( .A(n_360), .Y(n_414) );
INVxp67_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND5xp2_ASAP7_75t_L g367 ( .A(n_368), .B(n_375), .C(n_389), .D(n_395), .E(n_400), .Y(n_367) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
O2A1O1Ixp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_377), .B(n_378), .C(n_381), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AOI31xp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .A3(n_385), .B(n_386), .Y(n_381) );
INVx1_ASAP7_75t_L g407 ( .A(n_383), .Y(n_407) );
OR2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI222xp33_ASAP7_75t_L g410 ( .A1(n_397), .A2(n_399), .B1(n_411), .B2(n_414), .C1(n_415), .C2(n_416), .Y(n_410) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx2_ASAP7_75t_L g428 ( .A(n_421), .Y(n_428) );
NOR2x2_ASAP7_75t_L g726 ( .A(n_422), .B(n_440), .Y(n_726) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g439 ( .A(n_423), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
INVx1_ASAP7_75t_L g430 ( .A(n_428), .Y(n_430) );
NAND3xp33_ASAP7_75t_L g431 ( .A(n_429), .B(n_432), .C(n_730), .Y(n_431) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_437), .B1(n_438), .B2(n_441), .Y(n_434) );
INVx2_ASAP7_75t_L g728 ( .A(n_435), .Y(n_728) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI22xp5_ASAP7_75t_SL g727 ( .A1(n_437), .A2(n_441), .B1(n_728), .B2(n_729), .Y(n_727) );
INVx2_ASAP7_75t_L g729 ( .A(n_438), .Y(n_729) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OR3x1_ASAP7_75t_L g441 ( .A(n_442), .B(n_627), .C(n_676), .Y(n_441) );
NAND5xp2_ASAP7_75t_L g442 ( .A(n_443), .B(n_561), .C(n_590), .D(n_598), .E(n_613), .Y(n_442) );
O2A1O1Ixp33_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_489), .B(n_505), .C(n_545), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_445), .B(n_474), .Y(n_444) );
AND2x2_ASAP7_75t_L g556 ( .A(n_445), .B(n_553), .Y(n_556) );
AND2x2_ASAP7_75t_L g589 ( .A(n_445), .B(n_475), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_445), .B(n_493), .Y(n_682) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_462), .Y(n_445) );
INVx2_ASAP7_75t_L g492 ( .A(n_446), .Y(n_492) );
BUFx2_ASAP7_75t_L g656 ( .A(n_446), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_457), .Y(n_447) );
INVx5_ASAP7_75t_L g467 ( .A(n_449), .Y(n_467) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_SL g465 ( .A1(n_456), .A2(n_466), .B(n_467), .C(n_468), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_456), .A2(n_467), .B(n_532), .C(n_533), .Y(n_531) );
BUFx2_ASAP7_75t_L g478 ( .A(n_458), .Y(n_478) );
AND2x2_ASAP7_75t_L g474 ( .A(n_462), .B(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g554 ( .A(n_462), .Y(n_554) );
AND2x2_ASAP7_75t_L g640 ( .A(n_462), .B(n_553), .Y(n_640) );
AND2x2_ASAP7_75t_L g695 ( .A(n_462), .B(n_492), .Y(n_695) );
OA21x2_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_464), .B(n_473), .Y(n_462) );
INVx2_ASAP7_75t_L g498 ( .A(n_467), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVx1_ASAP7_75t_L g612 ( .A(n_474), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_474), .B(n_493), .Y(n_659) );
INVx5_ASAP7_75t_L g553 ( .A(n_475), .Y(n_553) );
AND2x4_ASAP7_75t_L g574 ( .A(n_475), .B(n_554), .Y(n_574) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_475), .Y(n_596) );
AND2x2_ASAP7_75t_L g671 ( .A(n_475), .B(n_656), .Y(n_671) );
AND2x2_ASAP7_75t_L g674 ( .A(n_475), .B(n_494), .Y(n_674) );
OR2x6_ASAP7_75t_L g475 ( .A(n_476), .B(n_486), .Y(n_475) );
AOI21xp5_ASAP7_75t_SL g476 ( .A1(n_477), .A2(n_479), .B(n_485), .Y(n_476) );
INVx2_ASAP7_75t_L g484 ( .A(n_482), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_484), .A2(n_500), .B(n_501), .C(n_502), .Y(n_499) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_484), .A2(n_502), .B(n_523), .C(n_524), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_489), .B(n_554), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_489), .B(n_685), .Y(n_684) );
INVx2_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_493), .Y(n_490) );
AND2x2_ASAP7_75t_L g579 ( .A(n_491), .B(n_554), .Y(n_579) );
AND2x2_ASAP7_75t_L g597 ( .A(n_491), .B(n_494), .Y(n_597) );
INVx1_ASAP7_75t_L g617 ( .A(n_491), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_491), .B(n_553), .Y(n_662) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_491), .Y(n_704) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_492), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_493), .B(n_552), .Y(n_551) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_493), .Y(n_606) );
O2A1O1Ixp33_ASAP7_75t_L g609 ( .A1(n_493), .A2(n_549), .B(n_610), .C(n_612), .Y(n_609) );
AND2x2_ASAP7_75t_L g616 ( .A(n_493), .B(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g625 ( .A(n_493), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g629 ( .A(n_493), .B(n_553), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_493), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g644 ( .A(n_493), .B(n_554), .Y(n_644) );
AND2x2_ASAP7_75t_L g694 ( .A(n_493), .B(n_695), .Y(n_694) );
INVx5_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx2_ASAP7_75t_L g558 ( .A(n_494), .Y(n_558) );
AND2x2_ASAP7_75t_L g599 ( .A(n_494), .B(n_552), .Y(n_599) );
AND2x2_ASAP7_75t_L g611 ( .A(n_494), .B(n_586), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_494), .B(n_640), .Y(n_658) );
OR2x6_ASAP7_75t_L g494 ( .A(n_495), .B(n_503), .Y(n_494) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_526), .Y(n_505) );
INVx1_ASAP7_75t_L g547 ( .A(n_506), .Y(n_547) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_518), .Y(n_506) );
OR2x2_ASAP7_75t_L g549 ( .A(n_507), .B(n_518), .Y(n_549) );
NAND3xp33_ASAP7_75t_L g555 ( .A(n_507), .B(n_556), .C(n_557), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_507), .B(n_528), .Y(n_566) );
OR2x2_ASAP7_75t_L g581 ( .A(n_507), .B(n_569), .Y(n_581) );
AND2x2_ASAP7_75t_L g587 ( .A(n_507), .B(n_537), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_507), .B(n_718), .Y(n_717) );
INVx5_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_508), .B(n_528), .Y(n_584) );
AND2x2_ASAP7_75t_L g623 ( .A(n_508), .B(n_538), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_508), .B(n_537), .Y(n_651) );
OR2x2_ASAP7_75t_L g654 ( .A(n_508), .B(n_537), .Y(n_654) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .B(n_512), .Y(n_509) );
INVx5_ASAP7_75t_SL g569 ( .A(n_518), .Y(n_569) );
OR2x2_ASAP7_75t_L g575 ( .A(n_518), .B(n_527), .Y(n_575) );
AND2x2_ASAP7_75t_L g591 ( .A(n_518), .B(n_592), .Y(n_591) );
AOI321xp33_ASAP7_75t_L g598 ( .A1(n_518), .A2(n_599), .A3(n_600), .B1(n_601), .B2(n_607), .C(n_609), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_518), .B(n_526), .Y(n_608) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_518), .Y(n_621) );
OR2x2_ASAP7_75t_L g668 ( .A(n_518), .B(n_566), .Y(n_668) );
AND2x2_ASAP7_75t_L g690 ( .A(n_518), .B(n_587), .Y(n_690) );
AND2x2_ASAP7_75t_L g709 ( .A(n_518), .B(n_528), .Y(n_709) );
OR2x6_ASAP7_75t_L g518 ( .A(n_519), .B(n_525), .Y(n_518) );
INVx1_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_537), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_528), .B(n_537), .Y(n_550) );
AND2x2_ASAP7_75t_L g559 ( .A(n_528), .B(n_560), .Y(n_559) );
INVx3_ASAP7_75t_L g586 ( .A(n_528), .Y(n_586) );
AND2x2_ASAP7_75t_L g592 ( .A(n_528), .B(n_587), .Y(n_592) );
INVxp67_ASAP7_75t_L g622 ( .A(n_528), .Y(n_622) );
OR2x2_ASAP7_75t_L g664 ( .A(n_528), .B(n_569), .Y(n_664) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_530), .B(n_536), .Y(n_528) );
OR2x2_ASAP7_75t_L g546 ( .A(n_537), .B(n_547), .Y(n_546) );
INVx1_ASAP7_75t_SL g560 ( .A(n_537), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_537), .B(n_549), .Y(n_593) );
AND2x2_ASAP7_75t_L g642 ( .A(n_537), .B(n_586), .Y(n_642) );
AND2x2_ASAP7_75t_L g680 ( .A(n_537), .B(n_569), .Y(n_680) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_538), .B(n_569), .Y(n_568) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_548), .B(n_551), .C(n_555), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_546), .A2(n_548), .B1(n_673), .B2(n_675), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_548), .A2(n_571), .B1(n_626), .B2(n_712), .Y(n_711) );
OR2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
INVx1_ASAP7_75t_SL g700 ( .A(n_549), .Y(n_700) );
INVx1_ASAP7_75t_SL g600 ( .A(n_550), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_552), .B(n_572), .Y(n_602) );
AOI222xp33_ASAP7_75t_L g613 ( .A1(n_552), .A2(n_593), .B1(n_600), .B2(n_614), .C1(n_618), .C2(n_624), .Y(n_613) );
AND2x2_ASAP7_75t_L g703 ( .A(n_552), .B(n_704), .Y(n_703) );
AND2x4_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
INVx2_ASAP7_75t_L g578 ( .A(n_553), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_553), .B(n_573), .Y(n_648) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_553), .Y(n_685) );
AND2x2_ASAP7_75t_L g688 ( .A(n_553), .B(n_597), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_553), .B(n_704), .Y(n_714) );
INVx1_ASAP7_75t_L g605 ( .A(n_554), .Y(n_605) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_554), .Y(n_633) );
O2A1O1Ixp33_ASAP7_75t_L g696 ( .A1(n_556), .A2(n_697), .B(n_698), .C(n_701), .Y(n_696) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
NAND3xp33_ASAP7_75t_L g619 ( .A(n_558), .B(n_620), .C(n_623), .Y(n_619) );
OR2x2_ASAP7_75t_L g647 ( .A(n_558), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_558), .B(n_574), .Y(n_675) );
OR2x2_ASAP7_75t_L g580 ( .A(n_560), .B(n_581), .Y(n_580) );
AOI211xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_564), .B(n_570), .C(n_582), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_563), .B(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g669 ( .A(n_564), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_565), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g583 ( .A(n_568), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_569), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g637 ( .A(n_569), .B(n_587), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_569), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_569), .B(n_586), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_575), .B1(n_576), .B2(n_580), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_572), .B(n_644), .Y(n_643) );
BUFx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_574), .B(n_616), .Y(n_615) );
OAI221xp5_ASAP7_75t_SL g638 ( .A1(n_575), .A2(n_639), .B1(n_641), .B2(n_643), .C(n_645), .Y(n_638) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
AND2x2_ASAP7_75t_L g693 ( .A(n_578), .B(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g706 ( .A(n_578), .B(n_695), .Y(n_706) );
INVx1_ASAP7_75t_L g626 ( .A(n_579), .Y(n_626) );
INVx1_ASAP7_75t_L g697 ( .A(n_580), .Y(n_697) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_581), .A2(n_664), .B(n_687), .Y(n_686) );
AOI21xp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_585), .B(n_588), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OAI21xp5_ASAP7_75t_SL g590 ( .A1(n_591), .A2(n_593), .B(n_594), .Y(n_590) );
INVx1_ASAP7_75t_L g630 ( .A(n_591), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_592), .A2(n_678), .B1(n_681), .B2(n_683), .C(n_686), .Y(n_677) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_600), .A2(n_690), .B1(n_691), .B2(n_693), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx1_ASAP7_75t_L g666 ( .A(n_602), .Y(n_666) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NOR2xp67_ASAP7_75t_SL g604 ( .A(n_605), .B(n_606), .Y(n_604) );
AND2x2_ASAP7_75t_L g670 ( .A(n_606), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g635 ( .A(n_611), .Y(n_635) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_616), .B(n_640), .Y(n_692) );
INVxp67_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_622), .B(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g708 ( .A(n_623), .B(n_709), .Y(n_708) );
AND2x4_ASAP7_75t_L g715 ( .A(n_623), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI211xp5_ASAP7_75t_SL g627 ( .A1(n_628), .A2(n_630), .B(n_631), .C(n_665), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AOI211xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_634), .B(n_638), .C(n_657), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_SL g718 ( .A(n_642), .Y(n_718) );
AND2x2_ASAP7_75t_L g655 ( .A(n_644), .B(n_656), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_649), .B1(n_653), .B2(n_655), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
OR2x2_ASAP7_75t_L g663 ( .A(n_651), .B(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g716 ( .A(n_652), .Y(n_716) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AOI31xp33_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_659), .A3(n_660), .B(n_663), .Y(n_657) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AOI211xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_667), .B(n_669), .C(n_672), .Y(n_665) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
CKINVDCx16_ASAP7_75t_R g673 ( .A(n_674), .Y(n_673) );
NAND5xp2_ASAP7_75t_L g676 ( .A(n_677), .B(n_689), .C(n_696), .D(n_710), .E(n_713), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_688), .A2(n_714), .B1(n_715), .B2(n_717), .Y(n_713) );
INVx1_ASAP7_75t_SL g712 ( .A(n_690), .Y(n_712) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AOI21xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_705), .B(n_707), .Y(n_701) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVxp67_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
CKINVDCx14_ASAP7_75t_R g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
BUFx2_ASAP7_75t_L g741 ( .A(n_734), .Y(n_741) );
OR2x4_ASAP7_75t_L g734 ( .A(n_735), .B(n_737), .Y(n_734) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
endmodule