module fake_netlist_1_78_n_16 (n_3, n_1, n_2, n_0, n_16);
input n_3;
input n_1;
input n_2;
input n_0;
output n_16;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_9;
wire n_5;
wire n_14;
wire n_8;
wire n_15;
wire n_10;
wire n_7;
INVx3_ASAP7_75t_L g4 ( .A(n_1), .Y(n_4) );
NAND2xp5_ASAP7_75t_SL g5 ( .A(n_3), .B(n_1), .Y(n_5) );
INVx1_ASAP7_75t_L g6 ( .A(n_4), .Y(n_6) );
OAI21x1_ASAP7_75t_L g7 ( .A1(n_4), .A2(n_0), .B(n_1), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_6), .B(n_0), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_6), .Y(n_9) );
OR2x2_ASAP7_75t_L g10 ( .A(n_8), .B(n_6), .Y(n_10) );
OAI21xp5_ASAP7_75t_L g11 ( .A1(n_10), .A2(n_7), .B(n_9), .Y(n_11) );
NOR2xp67_ASAP7_75t_L g12 ( .A(n_10), .B(n_0), .Y(n_12) );
AOI211xp5_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_5), .B(n_7), .C(n_2), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_11), .B(n_7), .Y(n_14) );
HB1xp67_ASAP7_75t_L g15 ( .A(n_13), .Y(n_15) );
AOI21xp5_ASAP7_75t_L g16 ( .A1(n_15), .A2(n_14), .B(n_2), .Y(n_16) );
endmodule