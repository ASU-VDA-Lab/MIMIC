module fake_ariane_994_n_3047 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_347, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_349, n_346, n_214, n_348, n_2, n_32, n_379, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_372, n_377, n_15, n_23, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_350, n_291, n_344, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_333, n_376, n_221, n_321, n_86, n_361, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_378, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_118, n_121, n_353, n_22, n_241, n_29, n_357, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_351, n_39, n_359, n_155, n_127, n_3047);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_347;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_379;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_333;
input n_376;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_378;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_118;
input n_121;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_351;
input n_39;
input n_359;
input n_155;
input n_127;

output n_3047;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_2484;
wire n_2866;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_2993;
wire n_1916;
wire n_2879;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_2407;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_524;
wire n_2731;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_462;
wire n_1181;
wire n_1999;
wire n_410;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_737;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_2976;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_520;
wire n_870;
wire n_2547;
wire n_1453;
wire n_945;
wire n_958;
wire n_2554;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_2960;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_625;
wire n_557;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_559;
wire n_2233;
wire n_2370;
wire n_2663;
wire n_495;
wire n_2914;
wire n_1988;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_2782;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_2950;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_2847;
wire n_884;
wire n_1851;
wire n_2162;
wire n_3015;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_432;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_2885;
wire n_2098;
wire n_661;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_3003;
wire n_533;
wire n_2867;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_438;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_3013;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_612;
wire n_2739;
wire n_512;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2956;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1443;
wire n_1021;
wire n_491;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_2909;
wire n_1416;
wire n_1121;
wire n_490;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_2527;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_1716;
wire n_1872;
wire n_380;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_2703;
wire n_2926;
wire n_696;
wire n_1442;
wire n_482;
wire n_2620;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_762;
wire n_1468;
wire n_1661;
wire n_1253;
wire n_2791;
wire n_555;
wire n_2683;
wire n_804;
wire n_1656;
wire n_1382;
wire n_2970;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_514;
wire n_2748;
wire n_418;
wire n_2185;
wire n_3029;
wire n_2398;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_2015;
wire n_1972;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2952;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_2922;
wire n_436;
wire n_3000;
wire n_2871;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_2628;
wire n_619;
wire n_967;
wire n_1083;
wire n_437;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_615;
wire n_1139;
wire n_2836;
wire n_2439;
wire n_2864;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_2224;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_470;
wire n_2668;
wire n_2921;
wire n_1240;
wire n_3046;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_632;
wire n_477;
wire n_650;
wire n_2388;
wire n_425;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2762;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_382;
wire n_3014;
wire n_489;
wire n_2294;
wire n_2274;
wire n_2895;
wire n_2903;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_397;
wire n_2467;
wire n_2768;
wire n_471;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_2924;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_404;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_564;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_522;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_598;
wire n_3031;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_2980;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_2697;
wire n_1387;
wire n_466;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_552;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_2834;
wire n_2483;
wire n_441;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_2996;
wire n_1592;
wire n_637;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_2811;
wire n_3019;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_2983;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_405;
wire n_1611;
wire n_2122;
wire n_2975;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2998;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_481;
wire n_1609;
wire n_1053;
wire n_600;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_529;
wire n_3039;
wire n_2195;
wire n_502;
wire n_2194;
wire n_2937;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_3022;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_727;
wire n_699;
wire n_590;
wire n_1726;
wire n_2075;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_545;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_2853;
wire n_427;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_3035;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_390;
wire n_1156;
wire n_2741;
wire n_501;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_2962;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_735;
wire n_1005;
wire n_527;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_888;
wire n_845;
wire n_2894;
wire n_2300;
wire n_2949;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_551;
wire n_417;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_1844;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_2994;
wire n_534;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_2119;
wire n_1540;
wire n_1719;
wire n_2742;
wire n_1266;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_2946;
wire n_1734;
wire n_1860;
wire n_403;
wire n_3016;
wire n_2785;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_3024;
wire n_2772;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_2893;
wire n_2959;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_1867;
wire n_456;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_704;
wire n_2958;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_2468;
wire n_2171;
wire n_1243;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_2581;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_2992;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_1191;
wire n_618;
wire n_2492;
wire n_2939;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_2900;
wire n_797;
wire n_2026;
wire n_2912;
wire n_1786;
wire n_2627;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_602;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_474;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_2991;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_516;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_1733;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1856;
wire n_2016;
wire n_640;
wire n_2667;
wire n_2723;
wire n_2725;
wire n_2928;
wire n_1118;
wire n_943;
wire n_678;
wire n_2905;
wire n_2884;
wire n_651;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1807;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_2857;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2720;
wire n_2412;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_819;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_586;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_2936;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2986;
wire n_2320;
wire n_3017;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2890;
wire n_2911;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_566;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_2892;
wire n_1201;
wire n_1288;
wire n_2605;
wire n_858;
wire n_2796;
wire n_1185;
wire n_2475;
wire n_2804;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_2947;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_465;
wire n_1103;
wire n_825;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_3043;
wire n_1958;
wire n_2747;
wire n_3027;
wire n_467;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_644;
wire n_1197;
wire n_3011;
wire n_2820;
wire n_2613;
wire n_497;
wire n_1165;
wire n_2934;
wire n_1641;
wire n_538;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_2647;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_2343;
wire n_1048;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1603;
wire n_1370;
wire n_728;
wire n_413;
wire n_2401;
wire n_2935;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_2478;
wire n_685;
wire n_911;
wire n_2658;
wire n_623;
wire n_2608;
wire n_2920;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_3006;
wire n_2767;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_464;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_3008;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_3037;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_2963;
wire n_519;
wire n_384;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_2007;
wire n_1056;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_1653;
wire n_872;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_540;
wire n_692;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_2938;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_2931;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_493;
wire n_2977;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_2828;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_2927;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_2951;
wire n_580;
wire n_1579;
wire n_494;
wire n_2809;
wire n_2181;
wire n_2014;
wire n_434;
wire n_975;
wire n_2974;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2972;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_2858;
wire n_972;
wire n_2251;
wire n_2923;
wire n_2843;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2872;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_2941;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_3034;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_541;
wire n_499;
wire n_2604;
wire n_1775;
wire n_788;
wire n_908;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_2630;
wire n_591;
wire n_2794;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2901;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_1630;
wire n_679;
wire n_1720;
wire n_663;
wire n_2409;
wire n_2966;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_3040;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_2597;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_2787;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_385;
wire n_2395;
wire n_917;
wire n_2868;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_631;
wire n_399;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_898;
wire n_857;
wire n_3042;
wire n_1067;
wire n_968;
wire n_1323;
wire n_1235;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_2967;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_2948;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_2897;
wire n_816;
wire n_1322;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2580;
wire n_2355;
wire n_1390;
wire n_2699;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_2973;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_3038;
wire n_759;
wire n_567;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_614;
wire n_2775;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_550;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_3001;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_671;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2933;
wire n_2856;
wire n_2088;
wire n_1275;
wire n_488;
wire n_3018;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_3028;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_459;
wire n_2515;
wire n_1782;
wire n_458;
wire n_1600;
wire n_1190;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_2846;
wire n_1781;
wire n_709;
wire n_2917;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_3032;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_3020;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_2513;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_2957;
wire n_865;
wire n_1273;
wire n_1983;
wire n_2982;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_860;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_450;
wire n_1923;
wire n_2955;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_902;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_954;
wire n_596;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_2673;
wire n_664;
wire n_1591;
wire n_2585;
wire n_2995;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_537;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_389;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_2875;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_2792;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1368;
wire n_1211;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1722;
wire n_1001;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_3030;
wire n_1339;
wire n_1644;
wire n_1002;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_719;
wire n_2255;
wire n_1252;
wire n_1129;
wire n_2239;
wire n_3045;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2798;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2940;
wire n_548;
wire n_2336;
wire n_523;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_457;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2915;
wire n_431;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_412;
wire n_1251;
wire n_1989;
wire n_3041;
wire n_447;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_3033;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_2953;
wire n_1308;
wire n_796;
wire n_573;
wire n_2851;
wire n_2823;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

BUFx2_ASAP7_75t_L g380 ( 
.A(n_370),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_141),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_337),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_322),
.Y(n_383)
);

CKINVDCx14_ASAP7_75t_R g384 ( 
.A(n_246),
.Y(n_384)
);

BUFx10_ASAP7_75t_L g385 ( 
.A(n_148),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_312),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_147),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_27),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_281),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_351),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_316),
.Y(n_391)
);

BUFx5_ASAP7_75t_L g392 ( 
.A(n_156),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_306),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_8),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_372),
.Y(n_395)
);

BUFx10_ASAP7_75t_L g396 ( 
.A(n_107),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_103),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_65),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_130),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_147),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_36),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_12),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_184),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_374),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_340),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_365),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g407 ( 
.A(n_43),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_240),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_119),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_271),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_164),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_83),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_292),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_280),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_61),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_33),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_36),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_362),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_328),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_106),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_91),
.Y(n_421)
);

INVx4_ASAP7_75t_R g422 ( 
.A(n_284),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_352),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_176),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_20),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_114),
.Y(n_426)
);

BUFx2_ASAP7_75t_SL g427 ( 
.A(n_111),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_378),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_124),
.Y(n_429)
);

BUFx2_ASAP7_75t_SL g430 ( 
.A(n_229),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_57),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_213),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_77),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_205),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_210),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_166),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_222),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_373),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_7),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_218),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_43),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_300),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_180),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_379),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_160),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_196),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_342),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_371),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_131),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_301),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_11),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_375),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_7),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_238),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_54),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_223),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_202),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_94),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_76),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_39),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_49),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_353),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_75),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_349),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_25),
.Y(n_465)
);

INVxp67_ASAP7_75t_SL g466 ( 
.A(n_366),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_168),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_358),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_45),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_188),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_112),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_355),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_338),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_339),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_256),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_203),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_178),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_346),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_211),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_143),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_92),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_89),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_75),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_46),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_264),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_149),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_148),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_121),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_276),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_334),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_152),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_175),
.Y(n_492)
);

BUFx5_ASAP7_75t_L g493 ( 
.A(n_308),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_87),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_164),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_242),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_267),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_132),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_14),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_109),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_93),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_344),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_105),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_61),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_191),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_170),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_98),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_250),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_331),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_27),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_326),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_127),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_18),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_313),
.Y(n_514)
);

BUFx2_ASAP7_75t_SL g515 ( 
.A(n_304),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_368),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_155),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_287),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_324),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_12),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_275),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_22),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_288),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_162),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_197),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_84),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_236),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_51),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_290),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_354),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_62),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_332),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_176),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_343),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_330),
.Y(n_535)
);

CKINVDCx16_ASAP7_75t_R g536 ( 
.A(n_181),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_258),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_347),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_263),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_94),
.Y(n_540)
);

CKINVDCx16_ASAP7_75t_R g541 ( 
.A(n_137),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_244),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_336),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_74),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_185),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_241),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_34),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_30),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_131),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_317),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_348),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_356),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_122),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_6),
.Y(n_554)
);

INVx1_ASAP7_75t_SL g555 ( 
.A(n_10),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_37),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_323),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_189),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_142),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_55),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_227),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_341),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_38),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_207),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_177),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_132),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_128),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_34),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_321),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_291),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_311),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_303),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_41),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_173),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_151),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_329),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_108),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_318),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_268),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_194),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_106),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_216),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_363),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_92),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_136),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_295),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_170),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_297),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_239),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_13),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_163),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_361),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_140),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_100),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_364),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_232),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_335),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_224),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_245),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_156),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_247),
.Y(n_601)
);

CKINVDCx16_ASAP7_75t_R g602 ( 
.A(n_234),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_155),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_157),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_22),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_187),
.Y(n_606)
);

CKINVDCx16_ASAP7_75t_R g607 ( 
.A(n_125),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_367),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_97),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_120),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_357),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_179),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_192),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_278),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_296),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_163),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_255),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_0),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_359),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_41),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_310),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_360),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_108),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_369),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_29),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_23),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_172),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_1),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_376),
.Y(n_629)
);

BUFx10_ASAP7_75t_L g630 ( 
.A(n_26),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_314),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_289),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_233),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_82),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_350),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_138),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_283),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_51),
.Y(n_638)
);

CKINVDCx14_ASAP7_75t_R g639 ( 
.A(n_315),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_333),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_73),
.Y(n_641)
);

CKINVDCx20_ASAP7_75t_R g642 ( 
.A(n_165),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_80),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_119),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_54),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_200),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_173),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_39),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_23),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_46),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_377),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_79),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_95),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_6),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_235),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_138),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_93),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_140),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_169),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_153),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_325),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_294),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_60),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_35),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_327),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_345),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_161),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_110),
.Y(n_668)
);

INVxp33_ASAP7_75t_R g669 ( 
.A(n_195),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_73),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_262),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_162),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_305),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_161),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_105),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_16),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_14),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_137),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_208),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_180),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_154),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_86),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_79),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_78),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_178),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_165),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_487),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_487),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_487),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_380),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_517),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_387),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_380),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_517),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_517),
.Y(n_695)
);

INVxp67_ASAP7_75t_SL g696 ( 
.A(n_649),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_649),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_649),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_402),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_402),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_440),
.Y(n_701)
);

CKINVDCx16_ASAP7_75t_R g702 ( 
.A(n_536),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_461),
.Y(n_703)
);

INVxp33_ASAP7_75t_SL g704 ( 
.A(n_528),
.Y(n_704)
);

CKINVDCx14_ASAP7_75t_R g705 ( 
.A(n_384),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_461),
.Y(n_706)
);

INVxp33_ASAP7_75t_L g707 ( 
.A(n_674),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_392),
.Y(n_708)
);

CKINVDCx16_ASAP7_75t_R g709 ( 
.A(n_541),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_392),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_392),
.Y(n_711)
);

INVxp67_ASAP7_75t_SL g712 ( 
.A(n_463),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_387),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_602),
.Y(n_714)
);

INVxp67_ASAP7_75t_SL g715 ( 
.A(n_463),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_392),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_629),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_494),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_494),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_392),
.Y(n_720)
);

INVxp33_ASAP7_75t_L g721 ( 
.A(n_658),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_392),
.Y(n_722)
);

INVxp33_ASAP7_75t_L g723 ( 
.A(n_658),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_675),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_392),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_629),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_392),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_408),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_382),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_382),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_389),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_629),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_389),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_607),
.Y(n_734)
);

INVxp33_ASAP7_75t_SL g735 ( 
.A(n_464),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_467),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_432),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_467),
.Y(n_738)
);

CKINVDCx16_ASAP7_75t_R g739 ( 
.A(n_385),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_483),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_483),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_675),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_560),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_446),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_560),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_468),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_648),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_648),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_654),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_654),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_478),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_398),
.Y(n_752)
);

INVxp33_ASAP7_75t_L g753 ( 
.A(n_398),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_395),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_420),
.Y(n_755)
);

INVxp33_ASAP7_75t_SL g756 ( 
.A(n_589),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_588),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_427),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_420),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_615),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_424),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_424),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_426),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_426),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_433),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_433),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_449),
.Y(n_767)
);

BUFx2_ASAP7_75t_SL g768 ( 
.A(n_632),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_666),
.Y(n_769)
);

CKINVDCx14_ASAP7_75t_R g770 ( 
.A(n_639),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_397),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_449),
.Y(n_772)
);

NOR2xp67_ASAP7_75t_L g773 ( 
.A(n_407),
.B(n_0),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_471),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_471),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_381),
.Y(n_776)
);

INVxp33_ASAP7_75t_SL g777 ( 
.A(n_388),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_477),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_477),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_480),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_480),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_481),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_431),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_481),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_482),
.Y(n_785)
);

INVxp33_ASAP7_75t_L g786 ( 
.A(n_482),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_429),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_394),
.Y(n_788)
);

INVxp67_ASAP7_75t_SL g789 ( 
.A(n_488),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_488),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_399),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_520),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_520),
.Y(n_793)
);

INVxp33_ASAP7_75t_SL g794 ( 
.A(n_400),
.Y(n_794)
);

BUFx3_ASAP7_75t_L g795 ( 
.A(n_393),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_385),
.B(n_1),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_395),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_441),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_427),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_544),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_544),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_547),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_547),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_548),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_401),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_548),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_553),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_553),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_554),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_412),
.Y(n_810)
);

INVxp67_ASAP7_75t_SL g811 ( 
.A(n_554),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_556),
.Y(n_812)
);

INVx1_ASAP7_75t_SL g813 ( 
.A(n_453),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_404),
.Y(n_814)
);

BUFx2_ASAP7_75t_L g815 ( 
.A(n_407),
.Y(n_815)
);

INVxp33_ASAP7_75t_L g816 ( 
.A(n_556),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_404),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_418),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_418),
.Y(n_819)
);

INVxp33_ASAP7_75t_SL g820 ( 
.A(n_415),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_416),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_428),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_417),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_559),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_559),
.Y(n_825)
);

INVxp67_ASAP7_75t_SL g826 ( 
.A(n_566),
.Y(n_826)
);

INVxp67_ASAP7_75t_SL g827 ( 
.A(n_566),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_393),
.Y(n_828)
);

INVx4_ASAP7_75t_L g829 ( 
.A(n_754),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_708),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_708),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_795),
.B(n_451),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_696),
.B(n_428),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_710),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_753),
.B(n_786),
.Y(n_835)
);

BUFx2_ASAP7_75t_L g836 ( 
.A(n_734),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_710),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_795),
.Y(n_838)
);

INVx5_ASAP7_75t_L g839 ( 
.A(n_754),
.Y(n_839)
);

AOI22x1_ASAP7_75t_SL g840 ( 
.A1(n_771),
.A2(n_522),
.B1(n_540),
.B2(n_486),
.Y(n_840)
);

AND2x6_ASAP7_75t_L g841 ( 
.A(n_729),
.B(n_447),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_816),
.B(n_385),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_711),
.Y(n_843)
);

NAND2x1p5_ASAP7_75t_L g844 ( 
.A(n_729),
.B(n_534),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_711),
.Y(n_845)
);

CKINVDCx6p67_ASAP7_75t_R g846 ( 
.A(n_768),
.Y(n_846)
);

INVx4_ASAP7_75t_L g847 ( 
.A(n_828),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_716),
.Y(n_848)
);

OAI21x1_ASAP7_75t_L g849 ( 
.A1(n_716),
.A2(n_444),
.B(n_435),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_720),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_712),
.B(n_715),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_828),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_720),
.Y(n_853)
);

OA21x2_ASAP7_75t_L g854 ( 
.A1(n_722),
.A2(n_727),
.B(n_725),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_722),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_725),
.Y(n_856)
);

CKINVDCx6p67_ASAP7_75t_R g857 ( 
.A(n_768),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_705),
.B(n_770),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_727),
.Y(n_859)
);

INVx5_ASAP7_75t_L g860 ( 
.A(n_783),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_687),
.Y(n_861)
);

AND2x6_ASAP7_75t_L g862 ( 
.A(n_730),
.B(n_447),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_737),
.Y(n_863)
);

BUFx8_ASAP7_75t_SL g864 ( 
.A(n_787),
.Y(n_864)
);

INVx4_ASAP7_75t_L g865 ( 
.A(n_730),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_731),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_688),
.Y(n_867)
);

BUFx8_ASAP7_75t_L g868 ( 
.A(n_713),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_689),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_691),
.Y(n_870)
);

INVx5_ASAP7_75t_L g871 ( 
.A(n_783),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_694),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_731),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_695),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_733),
.Y(n_875)
);

INVx6_ASAP7_75t_L g876 ( 
.A(n_796),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_697),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_733),
.Y(n_878)
);

AND2x6_ASAP7_75t_L g879 ( 
.A(n_797),
.B(n_454),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_797),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_814),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_698),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_814),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_815),
.B(n_396),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_817),
.Y(n_885)
);

BUFx2_ASAP7_75t_L g886 ( 
.A(n_734),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_817),
.Y(n_887)
);

HB1xp67_ASAP7_75t_L g888 ( 
.A(n_702),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_699),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_704),
.A2(n_623),
.B1(n_642),
.B2(n_563),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_709),
.Y(n_891)
);

AND2x6_ASAP7_75t_L g892 ( 
.A(n_818),
.B(n_454),
.Y(n_892)
);

INVx5_ASAP7_75t_L g893 ( 
.A(n_783),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_818),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_819),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_819),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_776),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_822),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_822),
.Y(n_899)
);

AOI22x1_ASAP7_75t_SL g900 ( 
.A1(n_798),
.A2(n_682),
.B1(n_744),
.B2(n_728),
.Y(n_900)
);

NOR2x1_ASAP7_75t_L g901 ( 
.A(n_752),
.B(n_534),
.Y(n_901)
);

BUFx8_ASAP7_75t_SL g902 ( 
.A(n_757),
.Y(n_902)
);

INVxp33_ASAP7_75t_SL g903 ( 
.A(n_701),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_755),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_759),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_761),
.Y(n_906)
);

OA21x2_ASAP7_75t_L g907 ( 
.A1(n_762),
.A2(n_444),
.B(n_435),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_704),
.A2(n_409),
.B1(n_575),
.B2(n_555),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_763),
.Y(n_909)
);

BUFx12f_ASAP7_75t_L g910 ( 
.A(n_701),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_815),
.B(n_396),
.Y(n_911)
);

OA21x2_ASAP7_75t_L g912 ( 
.A1(n_764),
.A2(n_473),
.B(n_472),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_765),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_766),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_767),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_772),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_717),
.B(n_622),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_747),
.B(n_396),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_747),
.B(n_472),
.Y(n_919)
);

CKINVDCx16_ASAP7_75t_R g920 ( 
.A(n_739),
.Y(n_920)
);

BUFx12f_ASAP7_75t_L g921 ( 
.A(n_714),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_774),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_737),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_775),
.Y(n_924)
);

AOI22xp5_ASAP7_75t_L g925 ( 
.A1(n_735),
.A2(n_451),
.B1(n_425),
.B2(n_436),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_796),
.B(n_789),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_778),
.Y(n_927)
);

BUFx12f_ASAP7_75t_L g928 ( 
.A(n_714),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_779),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_780),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_781),
.Y(n_931)
);

OA21x2_ASAP7_75t_L g932 ( 
.A1(n_782),
.A2(n_475),
.B(n_473),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_784),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_811),
.B(n_431),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_785),
.Y(n_935)
);

OAI22x1_ASAP7_75t_SL g936 ( 
.A1(n_735),
.A2(n_421),
.B1(n_443),
.B2(n_439),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_790),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_792),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_793),
.Y(n_939)
);

INVxp67_ASAP7_75t_L g940 ( 
.A(n_813),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_776),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_800),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_700),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_801),
.Y(n_944)
);

INVx5_ASAP7_75t_L g945 ( 
.A(n_713),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_802),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_803),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_703),
.B(n_630),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_706),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_788),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_717),
.B(n_726),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_804),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_806),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_925),
.A2(n_756),
.B1(n_693),
.B2(n_690),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_855),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_830),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_830),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_926),
.B(n_726),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_830),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_830),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_855),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_835),
.B(n_826),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_855),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_926),
.B(n_827),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_859),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_926),
.B(n_732),
.Y(n_966)
);

AND2x2_ASAP7_75t_SL g967 ( 
.A(n_926),
.B(n_465),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_859),
.Y(n_968)
);

NAND3xp33_ASAP7_75t_L g969 ( 
.A(n_925),
.B(n_693),
.C(n_690),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_835),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_859),
.Y(n_971)
);

OAI21x1_ASAP7_75t_L g972 ( 
.A1(n_849),
.A2(n_508),
.B(n_475),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_847),
.B(n_777),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_866),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_848),
.Y(n_975)
);

INVxp67_ASAP7_75t_L g976 ( 
.A(n_940),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_866),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_848),
.Y(n_978)
);

NAND2xp33_ASAP7_75t_SL g979 ( 
.A(n_951),
.B(n_732),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_842),
.B(n_721),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_838),
.B(n_758),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_854),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_866),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_866),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_854),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_847),
.B(n_777),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_854),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_854),
.Y(n_988)
);

OR2x6_ASAP7_75t_L g989 ( 
.A(n_876),
.B(n_669),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_842),
.B(n_723),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_866),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_866),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_902),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_830),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_878),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_909),
.B(n_707),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_878),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_878),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_878),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_831),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_878),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_847),
.B(n_756),
.Y(n_1002)
);

AND2x6_ASAP7_75t_L g1003 ( 
.A(n_948),
.B(n_508),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_838),
.B(n_799),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_836),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_888),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_831),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_838),
.B(n_852),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_878),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_891),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_847),
.B(n_788),
.Y(n_1011)
);

OA21x2_ASAP7_75t_L g1012 ( 
.A1(n_849),
.A2(n_511),
.B(n_509),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_881),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_909),
.B(n_736),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_881),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_881),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_831),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_SL g1018 ( 
.A1(n_890),
.A2(n_751),
.B1(n_760),
.B2(n_746),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_831),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_945),
.B(n_794),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_853),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_851),
.B(n_794),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_881),
.Y(n_1023)
);

AND2x6_ASAP7_75t_L g1024 ( 
.A(n_948),
.B(n_509),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_881),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_853),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_853),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_852),
.B(n_773),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_881),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_883),
.Y(n_1030)
);

OR2x2_ASAP7_75t_L g1031 ( 
.A(n_920),
.B(n_724),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_853),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_883),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_945),
.B(n_820),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_853),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_843),
.A2(n_519),
.B(n_511),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_863),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_853),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_856),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_927),
.B(n_738),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_852),
.B(n_820),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_923),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_883),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_856),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_927),
.B(n_740),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_883),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_856),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_856),
.Y(n_1048)
);

CKINVDCx20_ASAP7_75t_R g1049 ( 
.A(n_864),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_856),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_836),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_856),
.Y(n_1052)
);

OA21x2_ASAP7_75t_L g1053 ( 
.A1(n_834),
.A2(n_521),
.B(n_519),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_883),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_843),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_883),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_886),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_843),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_843),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_885),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_845),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_845),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_885),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_885),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_885),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_845),
.Y(n_1066)
);

INVxp67_ASAP7_75t_L g1067 ( 
.A(n_886),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_845),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_885),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_885),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_918),
.A2(n_805),
.B1(n_810),
.B2(n_791),
.Y(n_1071)
);

NAND2xp33_ASAP7_75t_SL g1072 ( 
.A(n_897),
.B(n_791),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_945),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_896),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_834),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_837),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_896),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_896),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_865),
.B(n_805),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_896),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_945),
.B(n_810),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_837),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_850),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_896),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_896),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_898),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_850),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_898),
.Y(n_1088)
);

INVxp67_ASAP7_75t_L g1089 ( 
.A(n_868),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_898),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_898),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_899),
.Y(n_1092)
);

INVx1_ASAP7_75t_SL g1093 ( 
.A(n_846),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_904),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_930),
.B(n_741),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_899),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_899),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_910),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_899),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_930),
.B(n_743),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_873),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_894),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_904),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_894),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_873),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_875),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_875),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_846),
.Y(n_1108)
);

XNOR2x2_ASAP7_75t_L g1109 ( 
.A(n_908),
.B(n_577),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_880),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_910),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_880),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_865),
.B(n_821),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_904),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_887),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_895),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_904),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_865),
.B(n_821),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_895),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_887),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_904),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1101),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_967),
.A2(n_912),
.B1(n_932),
.B2(n_907),
.Y(n_1123)
);

INVx4_ASAP7_75t_L g1124 ( 
.A(n_1008),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1101),
.B(n_865),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_1005),
.B(n_920),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_1022),
.B(n_917),
.Y(n_1127)
);

INVx8_ASAP7_75t_L g1128 ( 
.A(n_1003),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1075),
.Y(n_1129)
);

NAND2xp33_ASAP7_75t_L g1130 ( 
.A(n_956),
.B(n_941),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_964),
.B(n_945),
.Y(n_1131)
);

INVxp67_ASAP7_75t_SL g1132 ( 
.A(n_982),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_1008),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1105),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1105),
.B(n_953),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1075),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1106),
.B(n_953),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1106),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1107),
.B(n_953),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1076),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_967),
.A2(n_912),
.B1(n_932),
.B2(n_907),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1076),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_980),
.B(n_990),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1082),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_993),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1107),
.B(n_953),
.Y(n_1146)
);

NAND2xp33_ASAP7_75t_L g1147 ( 
.A(n_956),
.B(n_950),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_980),
.B(n_884),
.Y(n_1148)
);

AND2x2_ASAP7_75t_SL g1149 ( 
.A(n_1053),
.B(n_907),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1110),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1082),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_1008),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_1094),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_964),
.Y(n_1154)
);

OA22x2_ASAP7_75t_L g1155 ( 
.A1(n_964),
.A2(n_890),
.B1(n_908),
.B2(n_742),
.Y(n_1155)
);

INVx2_ASAP7_75t_SL g1156 ( 
.A(n_1006),
.Y(n_1156)
);

BUFx10_ASAP7_75t_L g1157 ( 
.A(n_993),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1083),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1110),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1109),
.A2(n_912),
.B1(n_932),
.B2(n_907),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1083),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_SL g1162 ( 
.A(n_989),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1093),
.B(n_934),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1071),
.B(n_945),
.Y(n_1164)
);

INVx4_ASAP7_75t_L g1165 ( 
.A(n_981),
.Y(n_1165)
);

INVx1_ASAP7_75t_SL g1166 ( 
.A(n_1051),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1112),
.Y(n_1167)
);

NAND3xp33_ASAP7_75t_L g1168 ( 
.A(n_954),
.B(n_1041),
.C(n_1067),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_1108),
.B(n_934),
.Y(n_1169)
);

INVx4_ASAP7_75t_SL g1170 ( 
.A(n_1003),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_1049),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_958),
.B(n_903),
.Y(n_1172)
);

INVx5_ASAP7_75t_L g1173 ( 
.A(n_956),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1112),
.B(n_844),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1087),
.Y(n_1175)
);

INVx5_ASAP7_75t_L g1176 ( 
.A(n_956),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_976),
.B(n_857),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1115),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1115),
.B(n_844),
.Y(n_1179)
);

INVx4_ASAP7_75t_L g1180 ( 
.A(n_981),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_990),
.B(n_884),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1120),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1120),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1086),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_966),
.B(n_911),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_970),
.B(n_911),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1109),
.A2(n_932),
.B1(n_912),
.B2(n_934),
.Y(n_1187)
);

NAND2xp33_ASAP7_75t_L g1188 ( 
.A(n_956),
.B(n_844),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1094),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_981),
.B(n_934),
.Y(n_1190)
);

AND2x2_ASAP7_75t_SL g1191 ( 
.A(n_1053),
.B(n_521),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1086),
.B(n_876),
.Y(n_1192)
);

INVx6_ASAP7_75t_L g1193 ( 
.A(n_1004),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1087),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1097),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_1055),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1097),
.B(n_876),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1014),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1014),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_955),
.Y(n_1200)
);

OR2x6_ASAP7_75t_L g1201 ( 
.A(n_989),
.B(n_921),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_969),
.A2(n_833),
.B1(n_581),
.B2(n_584),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1040),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_955),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_1079),
.B(n_857),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1004),
.B(n_918),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1088),
.B(n_876),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1004),
.B(n_921),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1055),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_973),
.B(n_928),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1058),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1098),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1113),
.B(n_746),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_986),
.B(n_928),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1040),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1045),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1045),
.Y(n_1217)
);

OR2x6_ASAP7_75t_L g1218 ( 
.A(n_989),
.B(n_858),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1095),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_962),
.A2(n_841),
.B1(n_879),
.B2(n_862),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1118),
.B(n_889),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_962),
.A2(n_841),
.B1(n_879),
.B2(n_862),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_982),
.A2(n_841),
.B1(n_879),
.B2(n_862),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1088),
.B(n_829),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_970),
.A2(n_581),
.B1(n_584),
.B2(n_577),
.Y(n_1225)
);

INVx5_ASAP7_75t_L g1226 ( 
.A(n_959),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1002),
.B(n_889),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_996),
.B(n_751),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1095),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_1028),
.B(n_823),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1100),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1100),
.Y(n_1232)
);

NAND2xp33_ASAP7_75t_SL g1233 ( 
.A(n_1020),
.B(n_823),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_985),
.A2(n_841),
.B1(n_879),
.B2(n_862),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_1094),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_985),
.A2(n_988),
.B1(n_987),
.B2(n_1003),
.Y(n_1236)
);

OR2x6_ASAP7_75t_L g1237 ( 
.A(n_989),
.B(n_832),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1090),
.B(n_829),
.Y(n_1238)
);

INVx2_ASAP7_75t_SL g1239 ( 
.A(n_1006),
.Y(n_1239)
);

INVx4_ASAP7_75t_L g1240 ( 
.A(n_959),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_1098),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1028),
.B(n_832),
.Y(n_1242)
);

INVx4_ASAP7_75t_L g1243 ( 
.A(n_959),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_1111),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1111),
.Y(n_1245)
);

AND2x2_ASAP7_75t_SL g1246 ( 
.A(n_1053),
.B(n_527),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1094),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_1094),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1003),
.A2(n_829),
.B1(n_913),
.B2(n_906),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1090),
.B(n_829),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1011),
.B(n_889),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1091),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_987),
.A2(n_862),
.B1(n_879),
.B2(n_841),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_968),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1091),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1092),
.Y(n_1256)
);

NAND2xp33_ASAP7_75t_L g1257 ( 
.A(n_959),
.B(n_1019),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1031),
.B(n_760),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1010),
.Y(n_1259)
);

CKINVDCx11_ASAP7_75t_R g1260 ( 
.A(n_1037),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1092),
.B(n_1096),
.Y(n_1261)
);

INVx4_ASAP7_75t_L g1262 ( 
.A(n_959),
.Y(n_1262)
);

BUFx10_ASAP7_75t_L g1263 ( 
.A(n_1042),
.Y(n_1263)
);

INVx5_ASAP7_75t_L g1264 ( 
.A(n_960),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1096),
.Y(n_1265)
);

INVx4_ASAP7_75t_L g1266 ( 
.A(n_960),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1099),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1028),
.B(n_979),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_996),
.B(n_769),
.Y(n_1269)
);

OR2x6_ASAP7_75t_L g1270 ( 
.A(n_1089),
.B(n_832),
.Y(n_1270)
);

INVx6_ASAP7_75t_L g1271 ( 
.A(n_1103),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1034),
.B(n_943),
.Y(n_1272)
);

OR2x6_ASAP7_75t_L g1273 ( 
.A(n_1018),
.B(n_1031),
.Y(n_1273)
);

INVx2_ASAP7_75t_SL g1274 ( 
.A(n_1057),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1099),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1102),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1072),
.B(n_769),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_1103),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1102),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1003),
.B(n_719),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1104),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1103),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_988),
.A2(n_1024),
.B1(n_1003),
.B2(n_1104),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1003),
.B(n_724),
.Y(n_1284)
);

INVx3_ASAP7_75t_L g1285 ( 
.A(n_1058),
.Y(n_1285)
);

BUFx10_ASAP7_75t_L g1286 ( 
.A(n_1024),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_961),
.B(n_904),
.Y(n_1287)
);

INVxp67_ASAP7_75t_SL g1288 ( 
.A(n_1053),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1024),
.A2(n_862),
.B1(n_879),
.B2(n_841),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_968),
.Y(n_1290)
);

INVx4_ASAP7_75t_L g1291 ( 
.A(n_960),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_975),
.Y(n_1292)
);

INVx4_ASAP7_75t_L g1293 ( 
.A(n_960),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1081),
.B(n_943),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1024),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1024),
.B(n_692),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_975),
.Y(n_1297)
);

INVx1_ASAP7_75t_SL g1298 ( 
.A(n_1024),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_961),
.B(n_963),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_978),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1073),
.B(n_868),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_963),
.B(n_905),
.Y(n_1302)
);

AND2x6_ASAP7_75t_L g1303 ( 
.A(n_1059),
.B(n_1061),
.Y(n_1303)
);

AND2x6_ASAP7_75t_L g1304 ( 
.A(n_1059),
.B(n_832),
.Y(n_1304)
);

AND2x6_ASAP7_75t_L g1305 ( 
.A(n_1061),
.B(n_901),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1116),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1116),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_965),
.B(n_905),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_978),
.Y(n_1309)
);

BUFx6f_ASAP7_75t_L g1310 ( 
.A(n_1103),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_965),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1119),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1119),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_971),
.B(n_718),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_971),
.B(n_905),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1062),
.B(n_905),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1062),
.B(n_943),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1154),
.B(n_1024),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1122),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1155),
.A2(n_862),
.B1(n_879),
.B2(n_841),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_1153),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1154),
.B(n_1066),
.Y(n_1322)
);

INVxp67_ASAP7_75t_L g1323 ( 
.A(n_1166),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1200),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1127),
.B(n_861),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1193),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1127),
.A2(n_1069),
.B1(n_1070),
.B2(n_1063),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1168),
.B(n_1066),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1134),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1186),
.B(n_949),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1138),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1205),
.B(n_861),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1204),
.Y(n_1333)
);

BUFx12f_ASAP7_75t_L g1334 ( 
.A(n_1260),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1165),
.B(n_1180),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1150),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1213),
.B(n_1190),
.Y(n_1337)
);

NAND2xp33_ASAP7_75t_L g1338 ( 
.A(n_1128),
.B(n_1068),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_1153),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1159),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1148),
.B(n_949),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1193),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1190),
.B(n_861),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1165),
.B(n_1068),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1280),
.B(n_949),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1167),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1181),
.B(n_906),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1227),
.B(n_1284),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1143),
.B(n_913),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1227),
.B(n_914),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1170),
.B(n_1295),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1178),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1182),
.Y(n_1353)
);

INVx2_ASAP7_75t_SL g1354 ( 
.A(n_1245),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1254),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1261),
.A2(n_1299),
.B(n_1137),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1290),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1198),
.B(n_914),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1292),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1170),
.B(n_960),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1183),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1199),
.B(n_915),
.Y(n_1362)
);

INVx2_ASAP7_75t_SL g1363 ( 
.A(n_1156),
.Y(n_1363)
);

AOI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1193),
.A2(n_1069),
.B1(n_1070),
.B2(n_1063),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1228),
.B(n_915),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1203),
.B(n_924),
.Y(n_1366)
);

A2O1A1Ixp33_ASAP7_75t_L g1367 ( 
.A1(n_1174),
.A2(n_1036),
.B(n_1065),
.C(n_1064),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1215),
.B(n_924),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1216),
.B(n_935),
.Y(n_1369)
);

A2O1A1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1174),
.A2(n_1036),
.B(n_1065),
.C(n_1064),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1184),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_SL g1372 ( 
.A(n_1180),
.B(n_994),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1171),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1217),
.B(n_935),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1195),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_SL g1376 ( 
.A(n_1124),
.B(n_994),
.Y(n_1376)
);

INVx2_ASAP7_75t_SL g1377 ( 
.A(n_1239),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1219),
.B(n_944),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1317),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1229),
.B(n_944),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_1124),
.B(n_994),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1297),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1259),
.B(n_994),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_SL g1384 ( 
.A(n_1133),
.B(n_994),
.Y(n_1384)
);

INVx1_ASAP7_75t_SL g1385 ( 
.A(n_1126),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1252),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1300),
.Y(n_1387)
);

INVxp33_ASAP7_75t_L g1388 ( 
.A(n_1258),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_SL g1389 ( 
.A(n_1133),
.B(n_1017),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1231),
.B(n_946),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1309),
.Y(n_1391)
);

AOI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1296),
.A2(n_1069),
.B1(n_1070),
.B2(n_1063),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1311),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1145),
.Y(n_1394)
);

INVx4_ASAP7_75t_L g1395 ( 
.A(n_1128),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1232),
.B(n_946),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_SL g1397 ( 
.A(n_1152),
.B(n_1017),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1255),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1256),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1265),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1274),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1206),
.B(n_905),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_SL g1403 ( 
.A(n_1170),
.B(n_1017),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1163),
.B(n_905),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1163),
.B(n_916),
.Y(n_1405)
);

NOR3xp33_ASAP7_75t_L g1406 ( 
.A(n_1172),
.B(n_411),
.C(n_458),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1169),
.B(n_916),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1169),
.B(n_916),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1185),
.B(n_957),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1152),
.B(n_957),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1267),
.Y(n_1411)
);

OAI21xp33_ASAP7_75t_L g1412 ( 
.A1(n_1179),
.A2(n_460),
.B(n_445),
.Y(n_1412)
);

INVx8_ASAP7_75t_L g1413 ( 
.A(n_1128),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1275),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1132),
.B(n_916),
.Y(n_1415)
);

AO22x2_ASAP7_75t_L g1416 ( 
.A1(n_1202),
.A2(n_900),
.B1(n_840),
.B2(n_868),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1276),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_SL g1418 ( 
.A(n_1283),
.B(n_1017),
.Y(n_1418)
);

NAND3xp33_ASAP7_75t_L g1419 ( 
.A(n_1177),
.B(n_868),
.C(n_974),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_SL g1420 ( 
.A(n_1212),
.B(n_1241),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1132),
.B(n_916),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1207),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1279),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1155),
.A2(n_892),
.B1(n_952),
.B2(n_937),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1187),
.A2(n_892),
.B1(n_952),
.B2(n_937),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_SL g1426 ( 
.A(n_1283),
.B(n_1017),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1242),
.B(n_957),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1221),
.B(n_916),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1286),
.B(n_1298),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_SL g1430 ( 
.A(n_1286),
.B(n_1019),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_SL g1431 ( 
.A(n_1236),
.B(n_1019),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1269),
.B(n_931),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1314),
.B(n_931),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1301),
.B(n_1263),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1281),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1221),
.B(n_1304),
.Y(n_1436)
);

NOR2xp67_ASAP7_75t_L g1437 ( 
.A(n_1244),
.B(n_919),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1201),
.B(n_939),
.Y(n_1438)
);

BUFx3_ASAP7_75t_L g1439 ( 
.A(n_1157),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1304),
.B(n_922),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1304),
.B(n_922),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1179),
.A2(n_1044),
.B1(n_1027),
.B2(n_977),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1230),
.B(n_1027),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1307),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1263),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1131),
.B(n_1027),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1304),
.B(n_922),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1313),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1129),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1207),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1210),
.B(n_1044),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1153),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1214),
.B(n_1044),
.Y(n_1453)
);

NOR2x1p5_ASAP7_75t_L g1454 ( 
.A(n_1277),
.B(n_1157),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1304),
.B(n_922),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1251),
.B(n_922),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1237),
.B(n_939),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1251),
.B(n_922),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1187),
.B(n_929),
.Y(n_1459)
);

INVx3_ASAP7_75t_L g1460 ( 
.A(n_1271),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1224),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1273),
.B(n_947),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1224),
.Y(n_1463)
);

INVxp67_ASAP7_75t_L g1464 ( 
.A(n_1225),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1238),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1238),
.Y(n_1466)
);

AND3x1_ASAP7_75t_L g1467 ( 
.A(n_1249),
.B(n_936),
.C(n_616),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1135),
.B(n_929),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1135),
.B(n_929),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1319),
.Y(n_1470)
);

AND2x6_ASAP7_75t_L g1471 ( 
.A(n_1318),
.B(n_1413),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1324),
.Y(n_1472)
);

NOR2x1p5_ASAP7_75t_L g1473 ( 
.A(n_1394),
.B(n_1201),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1464),
.B(n_1202),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1337),
.B(n_1225),
.Y(n_1475)
);

BUFx3_ASAP7_75t_L g1476 ( 
.A(n_1373),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1324),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1333),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1349),
.B(n_1137),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1329),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1393),
.Y(n_1481)
);

NAND2xp33_ASAP7_75t_SL g1482 ( 
.A(n_1395),
.B(n_1236),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1413),
.Y(n_1483)
);

AOI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1388),
.A2(n_1273),
.B1(n_1208),
.B2(n_1237),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1331),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_1334),
.Y(n_1486)
);

INVxp67_ASAP7_75t_SL g1487 ( 
.A(n_1415),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1365),
.B(n_1139),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1432),
.B(n_1139),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1336),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1373),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1340),
.Y(n_1492)
);

BUFx2_ASAP7_75t_L g1493 ( 
.A(n_1323),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1385),
.B(n_1273),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1348),
.B(n_1191),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1350),
.A2(n_1146),
.B1(n_1125),
.B2(n_1192),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1333),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1346),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1413),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1330),
.B(n_1146),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1352),
.Y(n_1501)
);

INVx3_ASAP7_75t_L g1502 ( 
.A(n_1395),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1433),
.B(n_1237),
.Y(n_1503)
);

BUFx12f_ASAP7_75t_L g1504 ( 
.A(n_1354),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1353),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1321),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_1321),
.Y(n_1507)
);

NAND2xp33_ASAP7_75t_L g1508 ( 
.A(n_1321),
.B(n_1303),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1341),
.B(n_1125),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_SL g1510 ( 
.A(n_1436),
.B(n_1328),
.Y(n_1510)
);

NOR2x2_ASAP7_75t_L g1511 ( 
.A(n_1420),
.B(n_1201),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1325),
.B(n_1218),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1361),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1401),
.B(n_1218),
.Y(n_1514)
);

NOR2x1_ASAP7_75t_L g1515 ( 
.A(n_1454),
.B(n_1218),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1379),
.B(n_1272),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1371),
.Y(n_1517)
);

BUFx8_ASAP7_75t_L g1518 ( 
.A(n_1439),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1326),
.B(n_1270),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1375),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1386),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1355),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1398),
.Y(n_1523)
);

OR2x6_ASAP7_75t_L g1524 ( 
.A(n_1438),
.B(n_1270),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1347),
.B(n_1272),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1400),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1462),
.B(n_1270),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1461),
.B(n_1164),
.Y(n_1528)
);

NAND3xp33_ASAP7_75t_L g1529 ( 
.A(n_1328),
.B(n_1147),
.C(n_1130),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1326),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1355),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1414),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1393),
.Y(n_1533)
);

NOR2xp67_ASAP7_75t_L g1534 ( 
.A(n_1445),
.B(n_1268),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1417),
.Y(n_1535)
);

BUFx3_ASAP7_75t_L g1536 ( 
.A(n_1342),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1417),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1321),
.B(n_1191),
.Y(n_1538)
);

AND2x6_ASAP7_75t_SL g1539 ( 
.A(n_1443),
.B(n_900),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1363),
.A2(n_1233),
.B1(n_936),
.B2(n_1188),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1342),
.B(n_1173),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1423),
.Y(n_1542)
);

NOR2xp67_ASAP7_75t_L g1543 ( 
.A(n_1377),
.B(n_1294),
.Y(n_1543)
);

NOR2x1p5_ASAP7_75t_L g1544 ( 
.A(n_1439),
.B(n_947),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1423),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1345),
.B(n_1192),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1438),
.B(n_1173),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1435),
.Y(n_1548)
);

AND2x6_ASAP7_75t_L g1549 ( 
.A(n_1318),
.B(n_1136),
.Y(n_1549)
);

AOI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1467),
.A2(n_1437),
.B1(n_1434),
.B2(n_1451),
.Y(n_1550)
);

NAND2x1p5_ASAP7_75t_L g1551 ( 
.A(n_1351),
.B(n_1360),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_L g1552 ( 
.A(n_1343),
.B(n_1197),
.Y(n_1552)
);

NOR2x2_ASAP7_75t_L g1553 ( 
.A(n_1416),
.B(n_840),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1435),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1444),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1416),
.A2(n_1142),
.B1(n_1144),
.B2(n_1140),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1357),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_SL g1558 ( 
.A(n_1475),
.B(n_1419),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1547),
.B(n_1457),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1525),
.B(n_1332),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1474),
.B(n_1424),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_SL g1562 ( 
.A(n_1550),
.B(n_1339),
.Y(n_1562)
);

NAND2xp33_ASAP7_75t_SL g1563 ( 
.A(n_1488),
.B(n_1335),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_1479),
.B(n_1339),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1516),
.B(n_1424),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1493),
.B(n_1358),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1484),
.B(n_1339),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1512),
.B(n_1339),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_SL g1569 ( 
.A(n_1512),
.B(n_1452),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1489),
.B(n_1362),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_SL g1571 ( 
.A(n_1543),
.B(n_1452),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1500),
.B(n_1452),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1503),
.B(n_1366),
.Y(n_1573)
);

NAND2xp33_ASAP7_75t_SL g1574 ( 
.A(n_1544),
.B(n_1162),
.Y(n_1574)
);

NAND2xp33_ASAP7_75t_SL g1575 ( 
.A(n_1483),
.B(n_1162),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1519),
.B(n_1452),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1547),
.B(n_1460),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_SL g1578 ( 
.A(n_1519),
.B(n_1451),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1494),
.B(n_1527),
.Y(n_1579)
);

NAND2xp33_ASAP7_75t_SL g1580 ( 
.A(n_1483),
.B(n_1368),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1527),
.B(n_1369),
.Y(n_1581)
);

NAND2xp33_ASAP7_75t_SL g1582 ( 
.A(n_1499),
.B(n_1374),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1536),
.B(n_1460),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_SL g1584 ( 
.A(n_1491),
.B(n_1453),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1509),
.B(n_1453),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1470),
.B(n_1378),
.Y(n_1586)
);

NAND2xp33_ASAP7_75t_L g1587 ( 
.A(n_1471),
.B(n_1463),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_1514),
.B(n_1344),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1480),
.B(n_1485),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1514),
.B(n_1344),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1476),
.B(n_1322),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1476),
.B(n_1322),
.Y(n_1592)
);

NAND2xp33_ASAP7_75t_SL g1593 ( 
.A(n_1499),
.B(n_1380),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1536),
.B(n_1351),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1540),
.B(n_1392),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1524),
.B(n_1360),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_SL g1597 ( 
.A(n_1529),
.B(n_1465),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_SL g1598 ( 
.A(n_1552),
.B(n_1466),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1490),
.B(n_1492),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1552),
.B(n_1410),
.Y(n_1600)
);

NAND2xp33_ASAP7_75t_SL g1601 ( 
.A(n_1473),
.B(n_1390),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1498),
.B(n_1396),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1524),
.B(n_1416),
.Y(n_1603)
);

NAND2xp33_ASAP7_75t_SL g1604 ( 
.A(n_1502),
.B(n_1197),
.Y(n_1604)
);

NAND2xp33_ASAP7_75t_SL g1605 ( 
.A(n_1502),
.B(n_1422),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1546),
.B(n_1356),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_SL g1607 ( 
.A(n_1546),
.B(n_1442),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1501),
.B(n_1320),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1496),
.B(n_1428),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_SL g1610 ( 
.A(n_1510),
.B(n_1456),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1596),
.B(n_1506),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1581),
.B(n_1505),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1566),
.B(n_1513),
.Y(n_1613)
);

BUFx6f_ASAP7_75t_L g1614 ( 
.A(n_1596),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1573),
.B(n_1517),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1610),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1610),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1595),
.A2(n_1556),
.B1(n_1443),
.B2(n_1524),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1570),
.B(n_1520),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1589),
.Y(n_1620)
);

NAND2x1_ASAP7_75t_L g1621 ( 
.A(n_1594),
.B(n_1549),
.Y(n_1621)
);

BUFx6f_ASAP7_75t_L g1622 ( 
.A(n_1594),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1583),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1606),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1586),
.B(n_1521),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1559),
.B(n_1506),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1599),
.B(n_1510),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1606),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1579),
.B(n_1523),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1602),
.B(n_1526),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1598),
.B(n_1532),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1561),
.B(n_1538),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1559),
.B(n_1530),
.Y(n_1633)
);

INVx5_ASAP7_75t_L g1634 ( 
.A(n_1583),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1597),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1608),
.B(n_1538),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1568),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1564),
.Y(n_1638)
);

NAND3xp33_ASAP7_75t_SL g1639 ( 
.A(n_1601),
.B(n_1406),
.C(n_1556),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1609),
.Y(n_1640)
);

CKINVDCx20_ASAP7_75t_R g1641 ( 
.A(n_1584),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1572),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1609),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1607),
.B(n_1495),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_SL g1645 ( 
.A1(n_1577),
.A2(n_1486),
.B1(n_1553),
.B2(n_1504),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1607),
.B(n_1495),
.Y(n_1646)
);

AOI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1578),
.A2(n_1482),
.B1(n_1534),
.B2(n_1549),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1558),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1565),
.B(n_1530),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1588),
.A2(n_1482),
.B1(n_1549),
.B2(n_1515),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1577),
.B(n_1518),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1569),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1574),
.Y(n_1653)
);

INVx11_ASAP7_75t_L g1654 ( 
.A(n_1575),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1603),
.B(n_1535),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1600),
.B(n_1537),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1587),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1590),
.B(n_1542),
.Y(n_1658)
);

INVx5_ASAP7_75t_L g1659 ( 
.A(n_1605),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1560),
.Y(n_1660)
);

BUFx3_ASAP7_75t_L g1661 ( 
.A(n_1621),
.Y(n_1661)
);

AO21x2_ASAP7_75t_L g1662 ( 
.A1(n_1648),
.A2(n_1567),
.B(n_1562),
.Y(n_1662)
);

AND2x2_ASAP7_75t_SL g1663 ( 
.A(n_1657),
.B(n_1508),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1624),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1659),
.B(n_1507),
.Y(n_1665)
);

OAI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1648),
.A2(n_1585),
.B(n_1563),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1624),
.Y(n_1667)
);

INVxp67_ASAP7_75t_SL g1668 ( 
.A(n_1640),
.Y(n_1668)
);

AO21x2_ASAP7_75t_L g1669 ( 
.A1(n_1628),
.A2(n_1459),
.B(n_1370),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1628),
.Y(n_1670)
);

BUFx4f_ASAP7_75t_L g1671 ( 
.A(n_1657),
.Y(n_1671)
);

BUFx2_ASAP7_75t_R g1672 ( 
.A(n_1653),
.Y(n_1672)
);

INVx2_ASAP7_75t_SL g1673 ( 
.A(n_1659),
.Y(n_1673)
);

OAI21x1_ASAP7_75t_L g1674 ( 
.A1(n_1621),
.A2(n_1551),
.B(n_1458),
.Y(n_1674)
);

NAND2x1p5_ASAP7_75t_L g1675 ( 
.A(n_1659),
.B(n_1640),
.Y(n_1675)
);

OAI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1639),
.A2(n_1582),
.B(n_1580),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1627),
.B(n_1487),
.Y(n_1677)
);

INVx4_ASAP7_75t_L g1678 ( 
.A(n_1659),
.Y(n_1678)
);

INVx2_ASAP7_75t_SL g1679 ( 
.A(n_1659),
.Y(n_1679)
);

OAI21x1_ASAP7_75t_L g1680 ( 
.A1(n_1643),
.A2(n_1551),
.B(n_1528),
.Y(n_1680)
);

BUFx3_ASAP7_75t_L g1681 ( 
.A(n_1622),
.Y(n_1681)
);

BUFx2_ASAP7_75t_L g1682 ( 
.A(n_1643),
.Y(n_1682)
);

BUFx2_ASAP7_75t_SL g1683 ( 
.A(n_1659),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1616),
.Y(n_1684)
);

OAI21x1_ASAP7_75t_L g1685 ( 
.A1(n_1616),
.A2(n_1487),
.B(n_1469),
.Y(n_1685)
);

OAI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1617),
.A2(n_1468),
.B(n_1431),
.Y(n_1686)
);

AO21x2_ASAP7_75t_L g1687 ( 
.A1(n_1649),
.A2(n_1367),
.B(n_1288),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1627),
.B(n_1591),
.Y(n_1688)
);

CKINVDCx20_ASAP7_75t_R g1689 ( 
.A(n_1641),
.Y(n_1689)
);

CKINVDCx20_ASAP7_75t_R g1690 ( 
.A(n_1645),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1617),
.Y(n_1691)
);

OAI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1635),
.A2(n_1593),
.B(n_1592),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1644),
.Y(n_1693)
);

BUFx3_ASAP7_75t_L g1694 ( 
.A(n_1622),
.Y(n_1694)
);

BUFx8_ASAP7_75t_SL g1695 ( 
.A(n_1623),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1635),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1644),
.Y(n_1697)
);

OAI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1660),
.A2(n_1549),
.B(n_1246),
.Y(n_1698)
);

BUFx2_ASAP7_75t_R g1699 ( 
.A(n_1653),
.Y(n_1699)
);

AO21x2_ASAP7_75t_L g1700 ( 
.A1(n_1618),
.A2(n_1288),
.B(n_1431),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1622),
.Y(n_1701)
);

OAI21x1_ASAP7_75t_L g1702 ( 
.A1(n_1646),
.A2(n_972),
.B(n_1418),
.Y(n_1702)
);

INVx3_ASAP7_75t_L g1703 ( 
.A(n_1646),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1660),
.Y(n_1704)
);

INVx4_ASAP7_75t_L g1705 ( 
.A(n_1654),
.Y(n_1705)
);

INVx4_ASAP7_75t_L g1706 ( 
.A(n_1654),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1636),
.Y(n_1707)
);

AO21x2_ASAP7_75t_L g1708 ( 
.A1(n_1652),
.A2(n_1426),
.B(n_1418),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1636),
.Y(n_1709)
);

OAI21x1_ASAP7_75t_L g1710 ( 
.A1(n_1638),
.A2(n_972),
.B(n_1426),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1638),
.Y(n_1711)
);

OA21x2_ASAP7_75t_L g1712 ( 
.A1(n_1642),
.A2(n_1160),
.B(n_532),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1642),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1656),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1656),
.Y(n_1715)
);

NAND2x1p5_ASAP7_75t_L g1716 ( 
.A(n_1647),
.B(n_1507),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1652),
.Y(n_1717)
);

OAI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1612),
.A2(n_1549),
.B(n_1246),
.Y(n_1718)
);

BUFx3_ASAP7_75t_L g1719 ( 
.A(n_1622),
.Y(n_1719)
);

OAI21x1_ASAP7_75t_L g1720 ( 
.A1(n_1650),
.A2(n_1421),
.B(n_1430),
.Y(n_1720)
);

INVx3_ASAP7_75t_L g1721 ( 
.A(n_1622),
.Y(n_1721)
);

BUFx3_ASAP7_75t_L g1722 ( 
.A(n_1634),
.Y(n_1722)
);

INVx3_ASAP7_75t_L g1723 ( 
.A(n_1623),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1632),
.Y(n_1724)
);

AOI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1632),
.A2(n_1320),
.B1(n_1412),
.B2(n_616),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1655),
.Y(n_1726)
);

BUFx6f_ASAP7_75t_L g1727 ( 
.A(n_1634),
.Y(n_1727)
);

HB1xp67_ASAP7_75t_L g1728 ( 
.A(n_1620),
.Y(n_1728)
);

INVx3_ASAP7_75t_L g1729 ( 
.A(n_1623),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1655),
.B(n_1629),
.Y(n_1730)
);

OAI21x1_ASAP7_75t_L g1731 ( 
.A1(n_1658),
.A2(n_1430),
.B(n_1440),
.Y(n_1731)
);

OAI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1619),
.A2(n_1409),
.B(n_1427),
.Y(n_1732)
);

BUFx3_ASAP7_75t_L g1733 ( 
.A(n_1634),
.Y(n_1733)
);

AO21x2_ASAP7_75t_L g1734 ( 
.A1(n_1631),
.A2(n_1447),
.B(n_1441),
.Y(n_1734)
);

OA21x2_ASAP7_75t_L g1735 ( 
.A1(n_1625),
.A2(n_1160),
.B(n_532),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1634),
.B(n_1507),
.Y(n_1736)
);

BUFx4f_ASAP7_75t_SL g1737 ( 
.A(n_1626),
.Y(n_1737)
);

BUFx3_ASAP7_75t_L g1738 ( 
.A(n_1634),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1637),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1611),
.B(n_1507),
.Y(n_1740)
);

BUFx3_ASAP7_75t_L g1741 ( 
.A(n_1614),
.Y(n_1741)
);

INVx3_ASAP7_75t_L g1742 ( 
.A(n_1611),
.Y(n_1742)
);

OAI21xp5_ASAP7_75t_L g1743 ( 
.A1(n_1615),
.A2(n_1409),
.B(n_1427),
.Y(n_1743)
);

INVx3_ASAP7_75t_L g1744 ( 
.A(n_1611),
.Y(n_1744)
);

AOI21x1_ASAP7_75t_L g1745 ( 
.A1(n_1630),
.A2(n_1571),
.B(n_1576),
.Y(n_1745)
);

OAI21x1_ASAP7_75t_SL g1746 ( 
.A1(n_1637),
.A2(n_1450),
.B(n_1299),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1728),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1728),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1704),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1704),
.Y(n_1750)
);

BUFx8_ASAP7_75t_L g1751 ( 
.A(n_1689),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1696),
.Y(n_1752)
);

CKINVDCx6p67_ASAP7_75t_R g1753 ( 
.A(n_1690),
.Y(n_1753)
);

AO22x1_ASAP7_75t_L g1754 ( 
.A1(n_1676),
.A2(n_1629),
.B1(n_1651),
.B2(n_1613),
.Y(n_1754)
);

AOI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1725),
.A2(n_1633),
.B1(n_1614),
.B2(n_1626),
.Y(n_1755)
);

CKINVDCx11_ASAP7_75t_R g1756 ( 
.A(n_1705),
.Y(n_1756)
);

CKINVDCx20_ASAP7_75t_R g1757 ( 
.A(n_1695),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1696),
.Y(n_1758)
);

AOI22xp33_ASAP7_75t_L g1759 ( 
.A1(n_1735),
.A2(n_1614),
.B1(n_1481),
.B2(n_1472),
.Y(n_1759)
);

OAI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1725),
.A2(n_1614),
.B1(n_1626),
.B2(n_628),
.Y(n_1760)
);

OAI21xp5_ASAP7_75t_SL g1761 ( 
.A1(n_1676),
.A2(n_628),
.B(n_600),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_SL g1762 ( 
.A1(n_1735),
.A2(n_1614),
.B1(n_1539),
.B2(n_1511),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1730),
.B(n_600),
.Y(n_1763)
);

OAI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1671),
.A2(n_660),
.B1(n_664),
.B2(n_653),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_SL g1765 ( 
.A1(n_1735),
.A2(n_1545),
.B1(n_1554),
.B2(n_1548),
.Y(n_1765)
);

CKINVDCx6p67_ASAP7_75t_R g1766 ( 
.A(n_1705),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1714),
.Y(n_1767)
);

BUFx12f_ASAP7_75t_L g1768 ( 
.A(n_1705),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_L g1769 ( 
.A1(n_1735),
.A2(n_1472),
.B1(n_1478),
.B2(n_1477),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1713),
.Y(n_1770)
);

OAI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1718),
.A2(n_660),
.B1(n_664),
.B2(n_653),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1713),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1682),
.Y(n_1773)
);

OAI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1671),
.A2(n_676),
.B1(n_683),
.B2(n_672),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1713),
.Y(n_1775)
);

AND2x4_ASAP7_75t_SL g1776 ( 
.A(n_1705),
.B(n_1706),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1735),
.A2(n_1477),
.B1(n_1497),
.B2(n_1478),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1717),
.Y(n_1778)
);

OAI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1718),
.A2(n_676),
.B1(n_683),
.B2(n_672),
.Y(n_1779)
);

BUFx6f_ASAP7_75t_SL g1780 ( 
.A(n_1706),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1714),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1698),
.A2(n_1497),
.B1(n_1531),
.B2(n_1522),
.Y(n_1782)
);

CKINVDCx11_ASAP7_75t_R g1783 ( 
.A(n_1706),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1715),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1715),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1698),
.A2(n_1522),
.B1(n_1557),
.B2(n_1531),
.Y(n_1786)
);

AOI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1700),
.A2(n_503),
.B1(n_524),
.B2(n_465),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1700),
.A2(n_524),
.B1(n_647),
.B2(n_503),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1730),
.B(n_603),
.Y(n_1789)
);

AOI22xp33_ASAP7_75t_L g1790 ( 
.A1(n_1700),
.A2(n_1662),
.B1(n_1724),
.B2(n_1726),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1700),
.A2(n_1557),
.B1(n_1533),
.B2(n_1449),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1717),
.Y(n_1792)
);

INVx6_ASAP7_75t_L g1793 ( 
.A(n_1706),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1730),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1726),
.Y(n_1795)
);

INVx6_ASAP7_75t_L g1796 ( 
.A(n_1740),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1726),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1688),
.B(n_527),
.Y(n_1798)
);

OAI22x1_ASAP7_75t_SL g1799 ( 
.A1(n_1672),
.A2(n_459),
.B1(n_469),
.B2(n_455),
.Y(n_1799)
);

INVx6_ASAP7_75t_L g1800 ( 
.A(n_1740),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1717),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1739),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1684),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1684),
.Y(n_1804)
);

INVx6_ASAP7_75t_L g1805 ( 
.A(n_1740),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1684),
.Y(n_1806)
);

INVx8_ASAP7_75t_L g1807 ( 
.A(n_1740),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1703),
.B(n_605),
.Y(n_1808)
);

AOI22xp33_ASAP7_75t_L g1809 ( 
.A1(n_1662),
.A2(n_1449),
.B1(n_1158),
.B2(n_1161),
.Y(n_1809)
);

BUFx3_ASAP7_75t_L g1810 ( 
.A(n_1737),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1691),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1711),
.Y(n_1812)
);

OAI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1671),
.A2(n_1737),
.B1(n_1688),
.B2(n_1666),
.Y(n_1813)
);

INVx1_ASAP7_75t_SL g1814 ( 
.A(n_1682),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1691),
.Y(n_1815)
);

AOI22xp33_ASAP7_75t_SL g1816 ( 
.A1(n_1712),
.A2(n_1555),
.B1(n_630),
.B2(n_430),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1711),
.Y(n_1817)
);

INVx6_ASAP7_75t_L g1818 ( 
.A(n_1681),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1691),
.Y(n_1819)
);

CKINVDCx11_ASAP7_75t_R g1820 ( 
.A(n_1681),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1671),
.A2(n_1425),
.B1(n_647),
.B2(n_1327),
.Y(n_1821)
);

AOI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1662),
.A2(n_1175),
.B1(n_1194),
.B2(n_1151),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1707),
.Y(n_1823)
);

BUFx6f_ASAP7_75t_L g1824 ( 
.A(n_1727),
.Y(n_1824)
);

BUFx3_ASAP7_75t_L g1825 ( 
.A(n_1681),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_SL g1826 ( 
.A1(n_1712),
.A2(n_630),
.B1(n_430),
.B2(n_515),
.Y(n_1826)
);

CKINVDCx11_ASAP7_75t_R g1827 ( 
.A(n_1694),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1724),
.B(n_535),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1707),
.B(n_1709),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_L g1830 ( 
.A1(n_1662),
.A2(n_1359),
.B1(n_1387),
.B2(n_1382),
.Y(n_1830)
);

INVx1_ASAP7_75t_SL g1831 ( 
.A(n_1683),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1709),
.Y(n_1832)
);

INVx3_ASAP7_75t_L g1833 ( 
.A(n_1678),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1677),
.B(n_535),
.Y(n_1834)
);

CKINVDCx11_ASAP7_75t_R g1835 ( 
.A(n_1694),
.Y(n_1835)
);

BUFx4f_ASAP7_75t_L g1836 ( 
.A(n_1727),
.Y(n_1836)
);

INVx2_ASAP7_75t_SL g1837 ( 
.A(n_1694),
.Y(n_1837)
);

BUFx2_ASAP7_75t_L g1838 ( 
.A(n_1703),
.Y(n_1838)
);

INVx3_ASAP7_75t_L g1839 ( 
.A(n_1678),
.Y(n_1839)
);

CKINVDCx20_ASAP7_75t_R g1840 ( 
.A(n_1701),
.Y(n_1840)
);

OAI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1677),
.A2(n_538),
.B1(n_546),
.B2(n_537),
.Y(n_1841)
);

BUFx6f_ASAP7_75t_L g1842 ( 
.A(n_1727),
.Y(n_1842)
);

OAI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1666),
.A2(n_538),
.B1(n_546),
.B2(n_537),
.Y(n_1843)
);

INVx3_ASAP7_75t_L g1844 ( 
.A(n_1678),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1739),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1697),
.A2(n_1359),
.B1(n_1387),
.B2(n_1382),
.Y(n_1846)
);

OAI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1716),
.A2(n_569),
.B1(n_570),
.B2(n_551),
.Y(n_1847)
);

CKINVDCx11_ASAP7_75t_R g1848 ( 
.A(n_1701),
.Y(n_1848)
);

AOI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1732),
.A2(n_1425),
.B1(n_1604),
.B2(n_569),
.Y(n_1849)
);

AOI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1732),
.A2(n_633),
.B1(n_570),
.B2(n_571),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1693),
.Y(n_1851)
);

BUFx10_ASAP7_75t_L g1852 ( 
.A(n_1736),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_SL g1853 ( 
.A1(n_1712),
.A2(n_515),
.B1(n_582),
.B2(n_622),
.Y(n_1853)
);

OAI22x1_ASAP7_75t_L g1854 ( 
.A1(n_1675),
.A2(n_491),
.B1(n_492),
.B2(n_484),
.Y(n_1854)
);

INVx3_ASAP7_75t_L g1855 ( 
.A(n_1678),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1697),
.A2(n_1391),
.B1(n_1448),
.B2(n_1444),
.Y(n_1856)
);

BUFx2_ASAP7_75t_L g1857 ( 
.A(n_1703),
.Y(n_1857)
);

BUFx2_ASAP7_75t_L g1858 ( 
.A(n_1703),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1693),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1693),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1670),
.Y(n_1861)
);

INVx4_ASAP7_75t_L g1862 ( 
.A(n_1723),
.Y(n_1862)
);

AOI22xp33_ASAP7_75t_SL g1863 ( 
.A1(n_1712),
.A2(n_582),
.B1(n_571),
.B2(n_551),
.Y(n_1863)
);

AOI22xp33_ASAP7_75t_L g1864 ( 
.A1(n_1712),
.A2(n_1708),
.B1(n_1391),
.B2(n_1448),
.Y(n_1864)
);

OAI22xp33_ASAP7_75t_L g1865 ( 
.A1(n_1716),
.A2(n_595),
.B1(n_599),
.B2(n_592),
.Y(n_1865)
);

BUFx2_ASAP7_75t_SL g1866 ( 
.A(n_1673),
.Y(n_1866)
);

INVx6_ASAP7_75t_L g1867 ( 
.A(n_1701),
.Y(n_1867)
);

INVx6_ASAP7_75t_L g1868 ( 
.A(n_1719),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1670),
.Y(n_1869)
);

CKINVDCx11_ASAP7_75t_R g1870 ( 
.A(n_1719),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1742),
.B(n_807),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1719),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1664),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1708),
.A2(n_1663),
.B1(n_1746),
.B2(n_1357),
.Y(n_1874)
);

AOI22xp33_ASAP7_75t_SL g1875 ( 
.A1(n_1663),
.A2(n_595),
.B1(n_599),
.B2(n_592),
.Y(n_1875)
);

AOI22xp33_ASAP7_75t_SL g1876 ( 
.A1(n_1663),
.A2(n_611),
.B1(n_613),
.B2(n_606),
.Y(n_1876)
);

BUFx12f_ASAP7_75t_L g1877 ( 
.A(n_1736),
.Y(n_1877)
);

AOI22xp5_ASAP7_75t_SL g1878 ( 
.A1(n_1683),
.A2(n_1471),
.B1(n_498),
.B2(n_499),
.Y(n_1878)
);

BUFx2_ASAP7_75t_L g1879 ( 
.A(n_1742),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1742),
.B(n_808),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1741),
.Y(n_1881)
);

INVx3_ASAP7_75t_L g1882 ( 
.A(n_1661),
.Y(n_1882)
);

OAI21xp5_ASAP7_75t_SL g1883 ( 
.A1(n_1692),
.A2(n_617),
.B(n_606),
.Y(n_1883)
);

INVx6_ASAP7_75t_L g1884 ( 
.A(n_1741),
.Y(n_1884)
);

CKINVDCx11_ASAP7_75t_R g1885 ( 
.A(n_1741),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1664),
.Y(n_1886)
);

AOI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1743),
.A2(n_613),
.B1(n_617),
.B2(n_611),
.Y(n_1887)
);

BUFx12f_ASAP7_75t_L g1888 ( 
.A(n_1736),
.Y(n_1888)
);

OAI22xp33_ASAP7_75t_L g1889 ( 
.A1(n_1716),
.A2(n_633),
.B1(n_635),
.B2(n_624),
.Y(n_1889)
);

INVx3_ASAP7_75t_L g1890 ( 
.A(n_1661),
.Y(n_1890)
);

INVx3_ASAP7_75t_L g1891 ( 
.A(n_1661),
.Y(n_1891)
);

AOI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1708),
.A2(n_1746),
.B1(n_1305),
.B2(n_1743),
.Y(n_1892)
);

AOI22xp33_ASAP7_75t_L g1893 ( 
.A1(n_1708),
.A2(n_1305),
.B1(n_1411),
.B2(n_1399),
.Y(n_1893)
);

BUFx6f_ASAP7_75t_L g1894 ( 
.A(n_1727),
.Y(n_1894)
);

OAI21xp5_ASAP7_75t_SL g1895 ( 
.A1(n_1692),
.A2(n_635),
.B(n_624),
.Y(n_1895)
);

AOI22xp5_ASAP7_75t_SL g1896 ( 
.A1(n_1673),
.A2(n_1471),
.B1(n_500),
.B2(n_501),
.Y(n_1896)
);

CKINVDCx11_ASAP7_75t_R g1897 ( 
.A(n_1727),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1668),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1748),
.Y(n_1899)
);

OAI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1761),
.A2(n_1672),
.B1(n_1699),
.B2(n_1668),
.Y(n_1900)
);

CKINVDCx20_ASAP7_75t_R g1901 ( 
.A(n_1751),
.Y(n_1901)
);

AOI22xp33_ASAP7_75t_L g1902 ( 
.A1(n_1762),
.A2(n_1734),
.B1(n_1305),
.B2(n_1669),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1747),
.B(n_1667),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1794),
.B(n_1742),
.Y(n_1904)
);

OAI21x1_ASAP7_75t_L g1905 ( 
.A1(n_1787),
.A2(n_1685),
.B(n_1788),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_1751),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1770),
.Y(n_1907)
);

OAI21x1_ASAP7_75t_L g1908 ( 
.A1(n_1787),
.A2(n_1685),
.B(n_1731),
.Y(n_1908)
);

AOI22xp33_ASAP7_75t_L g1909 ( 
.A1(n_1771),
.A2(n_1734),
.B1(n_1305),
.B2(n_1669),
.Y(n_1909)
);

AOI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1883),
.A2(n_1716),
.B1(n_1679),
.B2(n_1673),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1808),
.B(n_1667),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1823),
.Y(n_1912)
);

AOI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1883),
.A2(n_1679),
.B(n_1675),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1832),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1869),
.Y(n_1915)
);

AOI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1895),
.A2(n_1679),
.B(n_1675),
.Y(n_1916)
);

OAI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1761),
.A2(n_1699),
.B1(n_1675),
.B2(n_1667),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1772),
.Y(n_1918)
);

AOI221xp5_ASAP7_75t_L g1919 ( 
.A1(n_1843),
.A2(n_506),
.B1(n_507),
.B2(n_504),
.C(n_495),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1775),
.Y(n_1920)
);

OAI21x1_ASAP7_75t_L g1921 ( 
.A1(n_1788),
.A2(n_1685),
.B(n_1731),
.Y(n_1921)
);

OAI22xp5_ASAP7_75t_SL g1922 ( 
.A1(n_1757),
.A2(n_1727),
.B1(n_1733),
.B2(n_1722),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_1753),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1778),
.Y(n_1924)
);

AO31x2_ASAP7_75t_L g1925 ( 
.A1(n_1813),
.A2(n_679),
.A3(n_1734),
.B(n_812),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1789),
.B(n_1667),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1749),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1750),
.Y(n_1928)
);

OAI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1895),
.A2(n_1680),
.B(n_1731),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1829),
.Y(n_1930)
);

OAI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1850),
.A2(n_1680),
.B(n_1745),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_SL g1932 ( 
.A(n_1813),
.B(n_1722),
.Y(n_1932)
);

OA21x2_ASAP7_75t_L g1933 ( 
.A1(n_1790),
.A2(n_1686),
.B(n_1680),
.Y(n_1933)
);

BUFx2_ASAP7_75t_L g1934 ( 
.A(n_1840),
.Y(n_1934)
);

AOI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1764),
.A2(n_1665),
.B(n_1674),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1767),
.Y(n_1936)
);

AOI22xp33_ASAP7_75t_L g1937 ( 
.A1(n_1779),
.A2(n_1734),
.B1(n_1305),
.B2(n_1669),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1802),
.B(n_1723),
.Y(n_1938)
);

OAI22xp5_ASAP7_75t_L g1939 ( 
.A1(n_1764),
.A2(n_1774),
.B1(n_1876),
.B2(n_1875),
.Y(n_1939)
);

AOI22xp33_ASAP7_75t_L g1940 ( 
.A1(n_1826),
.A2(n_1669),
.B1(n_1411),
.B2(n_1399),
.Y(n_1940)
);

O2A1O1Ixp33_ASAP7_75t_L g1941 ( 
.A1(n_1774),
.A2(n_679),
.B(n_490),
.C(n_809),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1781),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1792),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1784),
.Y(n_1944)
);

AOI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1816),
.A2(n_1744),
.B1(n_1405),
.B2(n_1407),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1801),
.Y(n_1946)
);

OA21x2_ASAP7_75t_L g1947 ( 
.A1(n_1898),
.A2(n_1686),
.B(n_1710),
.Y(n_1947)
);

OA21x2_ASAP7_75t_L g1948 ( 
.A1(n_1873),
.A2(n_1686),
.B(n_1710),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1754),
.A2(n_1665),
.B(n_1674),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1785),
.Y(n_1950)
);

AO21x2_ASAP7_75t_L g1951 ( 
.A1(n_1834),
.A2(n_1828),
.B(n_1798),
.Y(n_1951)
);

AOI21x1_ASAP7_75t_L g1952 ( 
.A1(n_1763),
.A2(n_1745),
.B(n_1665),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1752),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1758),
.Y(n_1954)
);

AO21x2_ASAP7_75t_L g1955 ( 
.A1(n_1847),
.A2(n_1687),
.B(n_1710),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1814),
.B(n_1723),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1861),
.Y(n_1957)
);

HB1xp67_ASAP7_75t_L g1958 ( 
.A(n_1773),
.Y(n_1958)
);

OAI21x1_ASAP7_75t_L g1959 ( 
.A1(n_1892),
.A2(n_1702),
.B(n_1674),
.Y(n_1959)
);

AOI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1821),
.A2(n_1665),
.B(n_1687),
.Y(n_1960)
);

AO31x2_ASAP7_75t_L g1961 ( 
.A1(n_1803),
.A2(n_825),
.A3(n_824),
.B(n_952),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1812),
.Y(n_1962)
);

OR2x2_ASAP7_75t_L g1963 ( 
.A(n_1814),
.B(n_1744),
.Y(n_1963)
);

A2O1A1Ixp33_ASAP7_75t_L g1964 ( 
.A1(n_1878),
.A2(n_1733),
.B(n_1738),
.C(n_1722),
.Y(n_1964)
);

OR2x2_ASAP7_75t_L g1965 ( 
.A(n_1886),
.B(n_1744),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1795),
.B(n_1744),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1817),
.Y(n_1967)
);

OAI22xp5_ASAP7_75t_L g1968 ( 
.A1(n_1850),
.A2(n_1723),
.B1(n_1729),
.B2(n_1727),
.Y(n_1968)
);

AOI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1821),
.A2(n_1687),
.B(n_1720),
.Y(n_1969)
);

AOI21xp5_ASAP7_75t_L g1970 ( 
.A1(n_1836),
.A2(n_1831),
.B(n_1849),
.Y(n_1970)
);

OAI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1887),
.A2(n_1729),
.B1(n_1738),
.B2(n_1733),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_SL g1972 ( 
.A(n_1810),
.B(n_1729),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1879),
.B(n_1729),
.Y(n_1973)
);

INVx2_ASAP7_75t_SL g1974 ( 
.A(n_1818),
.Y(n_1974)
);

OA21x2_ASAP7_75t_L g1975 ( 
.A1(n_1804),
.A2(n_1702),
.B(n_1720),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1838),
.B(n_1721),
.Y(n_1976)
);

INVx3_ASAP7_75t_L g1977 ( 
.A(n_1818),
.Y(n_1977)
);

INVx3_ASAP7_75t_L g1978 ( 
.A(n_1867),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1845),
.B(n_1721),
.Y(n_1979)
);

AOI22xp33_ASAP7_75t_SL g1980 ( 
.A1(n_1896),
.A2(n_1738),
.B1(n_1687),
.B2(n_1721),
.Y(n_1980)
);

OAI21x1_ASAP7_75t_L g1981 ( 
.A1(n_1874),
.A2(n_1702),
.B(n_1720),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1851),
.Y(n_1982)
);

OAI22xp5_ASAP7_75t_L g1983 ( 
.A1(n_1887),
.A2(n_1721),
.B1(n_1736),
.B2(n_510),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1797),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1859),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1860),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1806),
.Y(n_1987)
);

OR2x2_ASAP7_75t_L g1988 ( 
.A(n_1857),
.B(n_745),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1811),
.Y(n_1989)
);

INVx1_ASAP7_75t_SL g1990 ( 
.A(n_1820),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1858),
.B(n_1518),
.Y(n_1991)
);

AO31x2_ASAP7_75t_L g1992 ( 
.A1(n_1815),
.A2(n_1446),
.A3(n_749),
.B(n_750),
.Y(n_1992)
);

OAI21xp33_ASAP7_75t_L g1993 ( 
.A1(n_1849),
.A2(n_513),
.B(n_512),
.Y(n_1993)
);

AOI21xp5_ASAP7_75t_L g1994 ( 
.A1(n_1836),
.A2(n_1338),
.B(n_1403),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1819),
.Y(n_1995)
);

OAI21xp5_ASAP7_75t_L g1996 ( 
.A1(n_1878),
.A2(n_673),
.B(n_405),
.Y(n_1996)
);

OAI221xp5_ASAP7_75t_L g1997 ( 
.A1(n_1896),
.A2(n_531),
.B1(n_549),
.B2(n_533),
.C(n_526),
.Y(n_1997)
);

INVxp67_ASAP7_75t_L g1998 ( 
.A(n_1872),
.Y(n_1998)
);

A2O1A1Ixp33_ASAP7_75t_L g1999 ( 
.A1(n_1755),
.A2(n_466),
.B(n_567),
.C(n_565),
.Y(n_1999)
);

HB1xp67_ASAP7_75t_L g2000 ( 
.A(n_1881),
.Y(n_2000)
);

AO21x2_ASAP7_75t_L g2001 ( 
.A1(n_1865),
.A2(n_1889),
.B(n_1841),
.Y(n_2001)
);

AO31x2_ASAP7_75t_L g2002 ( 
.A1(n_1854),
.A2(n_1446),
.A3(n_748),
.B(n_1294),
.Y(n_2002)
);

INVx8_ASAP7_75t_L g2003 ( 
.A(n_1780),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_1756),
.Y(n_2004)
);

A2O1A1Ixp33_ASAP7_75t_L g2005 ( 
.A1(n_1755),
.A2(n_573),
.B(n_574),
.C(n_568),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1871),
.B(n_585),
.Y(n_2006)
);

AO31x2_ASAP7_75t_L g2007 ( 
.A1(n_1862),
.A2(n_867),
.A3(n_870),
.B(n_869),
.Y(n_2007)
);

OAI221xp5_ASAP7_75t_L g2008 ( 
.A1(n_1853),
.A2(n_591),
.B1(n_593),
.B2(n_590),
.C(n_587),
.Y(n_2008)
);

OA21x2_ASAP7_75t_L g2009 ( 
.A1(n_1791),
.A2(n_604),
.B(n_594),
.Y(n_2009)
);

AOI21xp5_ASAP7_75t_SL g2010 ( 
.A1(n_1780),
.A2(n_1541),
.B(n_1383),
.Y(n_2010)
);

NAND2x1p5_ASAP7_75t_L g2011 ( 
.A(n_1831),
.B(n_1541),
.Y(n_2011)
);

OAI21x1_ASAP7_75t_L g2012 ( 
.A1(n_1833),
.A2(n_1455),
.B(n_1402),
.Y(n_2012)
);

AOI21xp33_ASAP7_75t_L g2013 ( 
.A1(n_1880),
.A2(n_610),
.B(n_609),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1867),
.Y(n_2014)
);

HB1xp67_ASAP7_75t_L g2015 ( 
.A(n_1837),
.Y(n_2015)
);

BUFx3_ASAP7_75t_L g2016 ( 
.A(n_1783),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1825),
.Y(n_2017)
);

OA21x2_ASAP7_75t_L g2018 ( 
.A1(n_1759),
.A2(n_618),
.B(n_612),
.Y(n_2018)
);

OAI21xp33_ASAP7_75t_L g2019 ( 
.A1(n_1863),
.A2(n_1765),
.B(n_625),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1868),
.Y(n_2020)
);

AOI21xp33_ASAP7_75t_L g2021 ( 
.A1(n_1760),
.A2(n_626),
.B(n_620),
.Y(n_2021)
);

AND2x4_ASAP7_75t_L g2022 ( 
.A(n_1882),
.B(n_1890),
.Y(n_2022)
);

OR2x6_ASAP7_75t_L g2023 ( 
.A(n_1807),
.B(n_1403),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1868),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1882),
.B(n_627),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1890),
.B(n_634),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1827),
.B(n_2),
.Y(n_2027)
);

OAI21x1_ASAP7_75t_L g2028 ( 
.A1(n_1833),
.A2(n_1302),
.B(n_1287),
.Y(n_2028)
);

BUFx2_ASAP7_75t_L g2029 ( 
.A(n_1884),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1884),
.Y(n_2030)
);

AO21x2_ASAP7_75t_L g2031 ( 
.A1(n_1830),
.A2(n_1302),
.B(n_1287),
.Y(n_2031)
);

OA21x2_ASAP7_75t_L g2032 ( 
.A1(n_1864),
.A2(n_638),
.B(n_636),
.Y(n_2032)
);

BUFx4f_ASAP7_75t_SL g2033 ( 
.A(n_1768),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1891),
.B(n_641),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1796),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1835),
.B(n_2),
.Y(n_2036)
);

A2O1A1Ixp33_ASAP7_75t_L g2037 ( 
.A1(n_1799),
.A2(n_643),
.B(n_645),
.C(n_644),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1796),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1891),
.Y(n_2039)
);

BUFx2_ASAP7_75t_L g2040 ( 
.A(n_1824),
.Y(n_2040)
);

OR2x6_ASAP7_75t_L g2041 ( 
.A(n_1807),
.B(n_1404),
.Y(n_2041)
);

HB1xp67_ASAP7_75t_L g2042 ( 
.A(n_1862),
.Y(n_2042)
);

AND2x4_ASAP7_75t_L g2043 ( 
.A(n_1839),
.B(n_1471),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1800),
.Y(n_2044)
);

OAI22xp5_ASAP7_75t_L g2045 ( 
.A1(n_1766),
.A2(n_650),
.B1(n_656),
.B2(n_652),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1866),
.B(n_657),
.Y(n_2046)
);

OA21x2_ASAP7_75t_L g2047 ( 
.A1(n_1893),
.A2(n_663),
.B(n_659),
.Y(n_2047)
);

AOI21x1_ASAP7_75t_L g2048 ( 
.A1(n_1793),
.A2(n_901),
.B(n_869),
.Y(n_2048)
);

CKINVDCx5p33_ASAP7_75t_R g2049 ( 
.A(n_1906),
.Y(n_2049)
);

AND2x4_ASAP7_75t_L g2050 ( 
.A(n_1977),
.B(n_1839),
.Y(n_2050)
);

AOI22xp33_ASAP7_75t_L g2051 ( 
.A1(n_2001),
.A2(n_1786),
.B1(n_1782),
.B2(n_1809),
.Y(n_2051)
);

AOI22xp33_ASAP7_75t_L g2052 ( 
.A1(n_2001),
.A2(n_1822),
.B1(n_1846),
.B2(n_1856),
.Y(n_2052)
);

BUFx4f_ASAP7_75t_SL g2053 ( 
.A(n_1901),
.Y(n_2053)
);

AOI22xp33_ASAP7_75t_L g2054 ( 
.A1(n_2009),
.A2(n_1769),
.B1(n_1777),
.B2(n_1800),
.Y(n_2054)
);

OAI221xp5_ASAP7_75t_L g2055 ( 
.A1(n_1996),
.A2(n_667),
.B1(n_677),
.B2(n_670),
.C(n_668),
.Y(n_2055)
);

INVx3_ASAP7_75t_L g2056 ( 
.A(n_2022),
.Y(n_2056)
);

OAI22xp5_ASAP7_75t_L g2057 ( 
.A1(n_1900),
.A2(n_1793),
.B1(n_1776),
.B2(n_1844),
.Y(n_2057)
);

AOI22xp33_ASAP7_75t_SL g2058 ( 
.A1(n_1900),
.A2(n_1807),
.B1(n_1805),
.B2(n_1877),
.Y(n_2058)
);

OAI22xp33_ASAP7_75t_L g2059 ( 
.A1(n_1910),
.A2(n_1805),
.B1(n_1842),
.B2(n_1824),
.Y(n_2059)
);

AOI211xp5_ASAP7_75t_L g2060 ( 
.A1(n_1917),
.A2(n_680),
.B(n_681),
.C(n_678),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1953),
.Y(n_2061)
);

OAI221xp5_ASAP7_75t_L g2062 ( 
.A1(n_1996),
.A2(n_684),
.B1(n_686),
.B2(n_685),
.C(n_1824),
.Y(n_2062)
);

OAI211xp5_ASAP7_75t_SL g2063 ( 
.A1(n_2046),
.A2(n_1848),
.B(n_1885),
.C(n_1870),
.Y(n_2063)
);

BUFx4f_ASAP7_75t_SL g2064 ( 
.A(n_2016),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1930),
.B(n_1844),
.Y(n_2065)
);

OR2x2_ASAP7_75t_L g2066 ( 
.A(n_1958),
.B(n_1855),
.Y(n_2066)
);

AOI22xp33_ASAP7_75t_L g2067 ( 
.A1(n_2009),
.A2(n_1888),
.B1(n_1894),
.B2(n_1842),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1954),
.Y(n_2068)
);

BUFx3_ASAP7_75t_L g2069 ( 
.A(n_2004),
.Y(n_2069)
);

AOI22xp5_ASAP7_75t_L g2070 ( 
.A1(n_1939),
.A2(n_1842),
.B1(n_1894),
.B2(n_1897),
.Y(n_2070)
);

AOI22xp33_ASAP7_75t_L g2071 ( 
.A1(n_2032),
.A2(n_1894),
.B1(n_1852),
.B2(n_1408),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_2029),
.B(n_1855),
.Y(n_2072)
);

AOI221xp5_ASAP7_75t_L g2073 ( 
.A1(n_1997),
.A2(n_651),
.B1(n_601),
.B2(n_933),
.C(n_929),
.Y(n_2073)
);

AOI22xp33_ASAP7_75t_L g2074 ( 
.A1(n_2032),
.A2(n_1852),
.B1(n_1306),
.B2(n_1312),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1899),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_2014),
.B(n_3),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1987),
.Y(n_2077)
);

BUFx6f_ASAP7_75t_L g2078 ( 
.A(n_2003),
.Y(n_2078)
);

OAI22xp5_ASAP7_75t_L g2079 ( 
.A1(n_1917),
.A2(n_1364),
.B1(n_1222),
.B2(n_1220),
.Y(n_2079)
);

AOI221xp5_ASAP7_75t_L g2080 ( 
.A1(n_1939),
.A2(n_651),
.B1(n_601),
.B2(n_933),
.C(n_929),
.Y(n_2080)
);

HB1xp67_ASAP7_75t_L g2081 ( 
.A(n_1988),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1989),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_2020),
.B(n_3),
.Y(n_2083)
);

CKINVDCx5p33_ASAP7_75t_R g2084 ( 
.A(n_1923),
.Y(n_2084)
);

AO21x1_ASAP7_75t_SL g2085 ( 
.A1(n_1938),
.A2(n_1316),
.B(n_1315),
.Y(n_2085)
);

AOI22xp33_ASAP7_75t_L g2086 ( 
.A1(n_2047),
.A2(n_1429),
.B1(n_493),
.B2(n_892),
.Y(n_2086)
);

AOI22xp33_ASAP7_75t_L g2087 ( 
.A1(n_2047),
.A2(n_1429),
.B1(n_493),
.B2(n_892),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1903),
.B(n_4),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1995),
.Y(n_2089)
);

AOI221xp5_ASAP7_75t_L g2090 ( 
.A1(n_1993),
.A2(n_651),
.B1(n_601),
.B2(n_933),
.C(n_929),
.Y(n_2090)
);

OAI21xp5_ASAP7_75t_L g2091 ( 
.A1(n_1980),
.A2(n_1471),
.B(n_870),
.Y(n_2091)
);

BUFx3_ASAP7_75t_L g2092 ( 
.A(n_1934),
.Y(n_2092)
);

AOI21xp33_ASAP7_75t_L g2093 ( 
.A1(n_1951),
.A2(n_4),
.B(n_5),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1915),
.Y(n_2094)
);

AO31x2_ASAP7_75t_L g2095 ( 
.A1(n_1949),
.A2(n_872),
.A3(n_874),
.B(n_867),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_2024),
.B(n_5),
.Y(n_2096)
);

AOI222xp33_ASAP7_75t_L g2097 ( 
.A1(n_1993),
.A2(n_892),
.B1(n_651),
.B2(n_601),
.C1(n_874),
.C2(n_877),
.Y(n_2097)
);

OAI22xp33_ASAP7_75t_L g2098 ( 
.A1(n_1910),
.A2(n_651),
.B1(n_601),
.B2(n_386),
.Y(n_2098)
);

INVx1_ASAP7_75t_SL g2099 ( 
.A(n_1963),
.Y(n_2099)
);

OAI21xp5_ASAP7_75t_L g2100 ( 
.A1(n_1983),
.A2(n_877),
.B(n_872),
.Y(n_2100)
);

AOI33xp33_ASAP7_75t_L g2101 ( 
.A1(n_2027),
.A2(n_10),
.A3(n_13),
.B1(n_8),
.B2(n_9),
.B3(n_11),
.Y(n_2101)
);

AOI21x1_ASAP7_75t_L g2102 ( 
.A1(n_2025),
.A2(n_882),
.B(n_1308),
.Y(n_2102)
);

AOI22xp33_ASAP7_75t_L g2103 ( 
.A1(n_2018),
.A2(n_493),
.B1(n_892),
.B2(n_1308),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1907),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1926),
.B(n_9),
.Y(n_2105)
);

AOI22xp33_ASAP7_75t_L g2106 ( 
.A1(n_2018),
.A2(n_493),
.B1(n_892),
.B2(n_1315),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1951),
.B(n_15),
.Y(n_2107)
);

AOI22xp33_ASAP7_75t_SL g2108 ( 
.A1(n_1932),
.A2(n_1983),
.B1(n_1955),
.B2(n_2036),
.Y(n_2108)
);

AOI21xp5_ASAP7_75t_L g2109 ( 
.A1(n_1969),
.A2(n_1257),
.B(n_1372),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_2030),
.B(n_15),
.Y(n_2110)
);

AOI22xp33_ASAP7_75t_L g2111 ( 
.A1(n_2019),
.A2(n_493),
.B1(n_938),
.B2(n_933),
.Y(n_2111)
);

INVx4_ASAP7_75t_L g2112 ( 
.A(n_2003),
.Y(n_2112)
);

INVx4_ASAP7_75t_L g2113 ( 
.A(n_2003),
.Y(n_2113)
);

AOI21xp33_ASAP7_75t_L g2114 ( 
.A1(n_2026),
.A2(n_16),
.B(n_17),
.Y(n_2114)
);

AOI22xp33_ASAP7_75t_L g2115 ( 
.A1(n_2019),
.A2(n_493),
.B1(n_938),
.B2(n_933),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1927),
.Y(n_2116)
);

AOI221xp5_ASAP7_75t_L g2117 ( 
.A1(n_2021),
.A2(n_938),
.B1(n_942),
.B2(n_933),
.C(n_882),
.Y(n_2117)
);

OAI22xp5_ASAP7_75t_L g2118 ( 
.A1(n_1970),
.A2(n_1971),
.B1(n_1964),
.B2(n_1913),
.Y(n_2118)
);

INVx8_ASAP7_75t_L g2119 ( 
.A(n_2041),
.Y(n_2119)
);

NAND4xp25_ASAP7_75t_L g2120 ( 
.A(n_2045),
.B(n_19),
.C(n_17),
.D(n_18),
.Y(n_2120)
);

AOI22xp33_ASAP7_75t_L g2121 ( 
.A1(n_1902),
.A2(n_493),
.B1(n_942),
.B2(n_938),
.Y(n_2121)
);

AOI22xp33_ASAP7_75t_L g2122 ( 
.A1(n_1909),
.A2(n_1937),
.B1(n_1940),
.B2(n_1955),
.Y(n_2122)
);

AOI21xp5_ASAP7_75t_L g2123 ( 
.A1(n_1929),
.A2(n_1389),
.B(n_1384),
.Y(n_2123)
);

AOI22xp33_ASAP7_75t_L g2124 ( 
.A1(n_2031),
.A2(n_493),
.B1(n_942),
.B2(n_938),
.Y(n_2124)
);

NOR2xp33_ASAP7_75t_L g2125 ( 
.A(n_1990),
.B(n_19),
.Y(n_2125)
);

AOI21xp33_ASAP7_75t_L g2126 ( 
.A1(n_2034),
.A2(n_20),
.B(n_21),
.Y(n_2126)
);

A2O1A1Ixp33_ASAP7_75t_L g2127 ( 
.A1(n_1999),
.A2(n_2005),
.B(n_2037),
.C(n_1960),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1918),
.Y(n_2128)
);

AOI211xp5_ASAP7_75t_L g2129 ( 
.A1(n_2045),
.A2(n_25),
.B(n_21),
.C(n_24),
.Y(n_2129)
);

OAI221xp5_ASAP7_75t_L g2130 ( 
.A1(n_2006),
.A2(n_1222),
.B1(n_1220),
.B2(n_391),
.C(n_403),
.Y(n_2130)
);

AOI22xp33_ASAP7_75t_L g2131 ( 
.A1(n_2031),
.A2(n_938),
.B1(n_942),
.B2(n_974),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_1977),
.B(n_24),
.Y(n_2132)
);

HB1xp67_ASAP7_75t_SL g2133 ( 
.A(n_1974),
.Y(n_2133)
);

AOI22xp5_ASAP7_75t_L g2134 ( 
.A1(n_1932),
.A2(n_1381),
.B1(n_1376),
.B2(n_1397),
.Y(n_2134)
);

CKINVDCx5p33_ASAP7_75t_R g2135 ( 
.A(n_1990),
.Y(n_2135)
);

AND2x4_ASAP7_75t_L g2136 ( 
.A(n_1978),
.B(n_26),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1928),
.Y(n_2137)
);

OAI22xp5_ASAP7_75t_L g2138 ( 
.A1(n_1971),
.A2(n_1916),
.B1(n_2041),
.B2(n_1968),
.Y(n_2138)
);

AND2x4_ASAP7_75t_L g2139 ( 
.A(n_1978),
.B(n_28),
.Y(n_2139)
);

OAI22xp5_ASAP7_75t_L g2140 ( 
.A1(n_2041),
.A2(n_1410),
.B1(n_1289),
.B2(n_1261),
.Y(n_2140)
);

OAI22xp33_ASAP7_75t_L g2141 ( 
.A1(n_1968),
.A2(n_390),
.B1(n_406),
.B2(n_383),
.Y(n_2141)
);

OR2x2_ASAP7_75t_L g2142 ( 
.A(n_1965),
.B(n_28),
.Y(n_2142)
);

AOI221xp5_ASAP7_75t_L g2143 ( 
.A1(n_2021),
.A2(n_942),
.B1(n_414),
.B2(n_419),
.C(n_413),
.Y(n_2143)
);

AOI22xp33_ASAP7_75t_L g2144 ( 
.A1(n_1931),
.A2(n_942),
.B1(n_983),
.B2(n_977),
.Y(n_2144)
);

AOI22xp33_ASAP7_75t_L g2145 ( 
.A1(n_1931),
.A2(n_983),
.B1(n_991),
.B2(n_984),
.Y(n_2145)
);

AOI22xp33_ASAP7_75t_SL g2146 ( 
.A1(n_1929),
.A2(n_1933),
.B1(n_1905),
.B2(n_1922),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1912),
.B(n_29),
.Y(n_2147)
);

OAI22xp5_ASAP7_75t_L g2148 ( 
.A1(n_2011),
.A2(n_1289),
.B1(n_1209),
.B2(n_1211),
.Y(n_2148)
);

AOI22xp5_ASAP7_75t_L g2149 ( 
.A1(n_2044),
.A2(n_1149),
.B1(n_1303),
.B2(n_423),
.Y(n_2149)
);

AOI21xp33_ASAP7_75t_L g2150 ( 
.A1(n_1933),
.A2(n_30),
.B(n_31),
.Y(n_2150)
);

OR2x2_ASAP7_75t_L g2151 ( 
.A(n_1966),
.B(n_31),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_1914),
.B(n_32),
.Y(n_2152)
);

AOI221x1_ASAP7_75t_SL g2153 ( 
.A1(n_1991),
.A2(n_35),
.B1(n_32),
.B2(n_33),
.C(n_37),
.Y(n_2153)
);

NOR2xp67_ASAP7_75t_L g2154 ( 
.A(n_2042),
.B(n_38),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1957),
.Y(n_2155)
);

BUFx6f_ASAP7_75t_L g2156 ( 
.A(n_2048),
.Y(n_2156)
);

OAI22xp5_ASAP7_75t_L g2157 ( 
.A1(n_2011),
.A2(n_1209),
.B1(n_1211),
.B2(n_1196),
.Y(n_2157)
);

BUFx6f_ASAP7_75t_L g2158 ( 
.A(n_2028),
.Y(n_2158)
);

OAI22xp5_ASAP7_75t_L g2159 ( 
.A1(n_1922),
.A2(n_1285),
.B1(n_1196),
.B2(n_1141),
.Y(n_2159)
);

BUFx3_ASAP7_75t_L g2160 ( 
.A(n_2033),
.Y(n_2160)
);

AOI22xp33_ASAP7_75t_L g2161 ( 
.A1(n_2013),
.A2(n_984),
.B1(n_992),
.B2(n_991),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1920),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_2022),
.B(n_40),
.Y(n_2163)
);

NAND3xp33_ASAP7_75t_L g2164 ( 
.A(n_1941),
.B(n_434),
.C(n_410),
.Y(n_2164)
);

NOR2xp33_ASAP7_75t_L g2165 ( 
.A(n_2017),
.B(n_40),
.Y(n_2165)
);

OA21x2_ASAP7_75t_L g2166 ( 
.A1(n_2039),
.A2(n_1316),
.B(n_1141),
.Y(n_2166)
);

OAI221xp5_ASAP7_75t_L g2167 ( 
.A1(n_1919),
.A2(n_442),
.B1(n_448),
.B2(n_438),
.C(n_437),
.Y(n_2167)
);

INVx1_ASAP7_75t_SL g2168 ( 
.A(n_2015),
.Y(n_2168)
);

OA21x2_ASAP7_75t_L g2169 ( 
.A1(n_1956),
.A2(n_1123),
.B(n_995),
.Y(n_2169)
);

AND2x4_ASAP7_75t_L g2170 ( 
.A(n_2043),
.B(n_42),
.Y(n_2170)
);

AOI22xp33_ASAP7_75t_SL g2171 ( 
.A1(n_1981),
.A2(n_1149),
.B1(n_452),
.B2(n_456),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_1904),
.B(n_42),
.Y(n_2172)
);

AOI221xp5_ASAP7_75t_L g2173 ( 
.A1(n_2008),
.A2(n_462),
.B1(n_470),
.B2(n_457),
.C(n_450),
.Y(n_2173)
);

OAI22xp33_ASAP7_75t_L g2174 ( 
.A1(n_1935),
.A2(n_476),
.B1(n_479),
.B2(n_474),
.Y(n_2174)
);

INVxp67_ASAP7_75t_SL g2175 ( 
.A(n_2000),
.Y(n_2175)
);

AOI22xp33_ASAP7_75t_L g2176 ( 
.A1(n_1945),
.A2(n_992),
.B1(n_997),
.B2(n_995),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_1924),
.Y(n_2177)
);

AOI21xp5_ASAP7_75t_L g2178 ( 
.A1(n_2010),
.A2(n_1123),
.B(n_1250),
.Y(n_2178)
);

AOI221x1_ASAP7_75t_L g2179 ( 
.A1(n_2035),
.A2(n_998),
.B1(n_1001),
.B2(n_999),
.C(n_997),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1936),
.Y(n_2180)
);

AOI222xp33_ASAP7_75t_L g2181 ( 
.A1(n_1984),
.A2(n_871),
.B1(n_893),
.B2(n_860),
.C1(n_497),
.C2(n_489),
.Y(n_2181)
);

AOI22xp33_ASAP7_75t_L g2182 ( 
.A1(n_2038),
.A2(n_998),
.B1(n_1001),
.B2(n_999),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1942),
.Y(n_2183)
);

AOI22xp33_ASAP7_75t_L g2184 ( 
.A1(n_1943),
.A2(n_1009),
.B1(n_1015),
.B2(n_1013),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1944),
.Y(n_2185)
);

AO31x2_ASAP7_75t_L g2186 ( 
.A1(n_1985),
.A2(n_1013),
.A3(n_1015),
.B(n_1009),
.Y(n_2186)
);

OAI22xp33_ASAP7_75t_L g2187 ( 
.A1(n_2023),
.A2(n_496),
.B1(n_502),
.B2(n_485),
.Y(n_2187)
);

AOI21xp5_ASAP7_75t_L g2188 ( 
.A1(n_1972),
.A2(n_1250),
.B(n_1234),
.Y(n_2188)
);

AOI21xp5_ASAP7_75t_L g2189 ( 
.A1(n_1911),
.A2(n_1234),
.B(n_1223),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_1950),
.B(n_44),
.Y(n_2190)
);

OAI22xp5_ASAP7_75t_L g2191 ( 
.A1(n_2043),
.A2(n_1285),
.B1(n_514),
.B2(n_516),
.Y(n_2191)
);

HB1xp67_ASAP7_75t_L g2192 ( 
.A(n_1986),
.Y(n_2192)
);

AOI22xp33_ASAP7_75t_L g2193 ( 
.A1(n_1946),
.A2(n_1982),
.B1(n_1962),
.B2(n_1967),
.Y(n_2193)
);

OAI33xp33_ASAP7_75t_L g2194 ( 
.A1(n_1998),
.A2(n_505),
.A3(n_518),
.B1(n_523),
.B2(n_525),
.B3(n_529),
.Y(n_2194)
);

AOI21xp33_ASAP7_75t_L g2195 ( 
.A1(n_1948),
.A2(n_44),
.B(n_45),
.Y(n_2195)
);

AOI22xp33_ASAP7_75t_L g2196 ( 
.A1(n_1959),
.A2(n_1016),
.B1(n_1025),
.B2(n_1023),
.Y(n_2196)
);

OAI22xp33_ASAP7_75t_L g2197 ( 
.A1(n_2023),
.A2(n_539),
.B1(n_542),
.B2(n_530),
.Y(n_2197)
);

AOI22xp33_ASAP7_75t_L g2198 ( 
.A1(n_2023),
.A2(n_1016),
.B1(n_1025),
.B2(n_1023),
.Y(n_2198)
);

AOI221xp5_ASAP7_75t_L g2199 ( 
.A1(n_1979),
.A2(n_1925),
.B1(n_550),
.B2(n_552),
.C(n_545),
.Y(n_2199)
);

BUFx2_ASAP7_75t_L g2200 ( 
.A(n_1973),
.Y(n_2200)
);

OAI22xp33_ASAP7_75t_L g2201 ( 
.A1(n_1952),
.A2(n_557),
.B1(n_558),
.B2(n_543),
.Y(n_2201)
);

HB1xp67_ASAP7_75t_L g2202 ( 
.A(n_2081),
.Y(n_2202)
);

HB1xp67_ASAP7_75t_L g2203 ( 
.A(n_2192),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_2056),
.B(n_1976),
.Y(n_2204)
);

BUFx2_ASAP7_75t_L g2205 ( 
.A(n_2056),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_2200),
.B(n_2040),
.Y(n_2206)
);

INVx3_ASAP7_75t_L g2207 ( 
.A(n_2158),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2077),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2082),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2104),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2128),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2089),
.Y(n_2212)
);

AOI21x1_ASAP7_75t_L g2213 ( 
.A1(n_2107),
.A2(n_2154),
.B(n_2088),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2094),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2099),
.B(n_1948),
.Y(n_2215)
);

BUFx2_ASAP7_75t_L g2216 ( 
.A(n_2112),
.Y(n_2216)
);

INVx3_ASAP7_75t_L g2217 ( 
.A(n_2158),
.Y(n_2217)
);

BUFx2_ASAP7_75t_L g2218 ( 
.A(n_2112),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2116),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_2162),
.Y(n_2220)
);

BUFx2_ASAP7_75t_L g2221 ( 
.A(n_2113),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_2177),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2137),
.Y(n_2223)
);

OR2x2_ASAP7_75t_L g2224 ( 
.A(n_2099),
.B(n_1925),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2180),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_2158),
.Y(n_2226)
);

INVx1_ASAP7_75t_SL g2227 ( 
.A(n_2053),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2072),
.B(n_2050),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2183),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_2075),
.B(n_1925),
.Y(n_2230)
);

HB1xp67_ASAP7_75t_L g2231 ( 
.A(n_2175),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_2050),
.B(n_1947),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_2168),
.B(n_1947),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2061),
.B(n_1975),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2185),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_2066),
.B(n_1975),
.Y(n_2236)
);

BUFx3_ASAP7_75t_L g2237 ( 
.A(n_2064),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2146),
.B(n_2007),
.Y(n_2238)
);

INVx1_ASAP7_75t_SL g2239 ( 
.A(n_2135),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2068),
.B(n_1961),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2108),
.B(n_1961),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_2155),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2147),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_2138),
.B(n_2007),
.Y(n_2244)
);

OAI22xp5_ASAP7_75t_L g2245 ( 
.A1(n_2070),
.A2(n_1994),
.B1(n_2002),
.B2(n_2012),
.Y(n_2245)
);

AND2x4_ASAP7_75t_L g2246 ( 
.A(n_2113),
.B(n_2007),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_2151),
.Y(n_2247)
);

INVx2_ASAP7_75t_SL g2248 ( 
.A(n_2078),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_2142),
.B(n_1908),
.Y(n_2249)
);

HB1xp67_ASAP7_75t_L g2250 ( 
.A(n_2065),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2172),
.B(n_1921),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_2186),
.Y(n_2252)
);

HB1xp67_ASAP7_75t_L g2253 ( 
.A(n_2152),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2190),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2092),
.B(n_1961),
.Y(n_2255)
);

OAI22xp5_ASAP7_75t_L g2256 ( 
.A1(n_2060),
.A2(n_2002),
.B1(n_1992),
.B2(n_1253),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2105),
.B(n_1992),
.Y(n_2257)
);

INVxp67_ASAP7_75t_SL g2258 ( 
.A(n_2133),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2186),
.Y(n_2259)
);

HB1xp67_ASAP7_75t_L g2260 ( 
.A(n_2118),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2186),
.Y(n_2261)
);

AND2x4_ASAP7_75t_L g2262 ( 
.A(n_2170),
.B(n_1992),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2193),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_2156),
.Y(n_2264)
);

AND2x4_ASAP7_75t_L g2265 ( 
.A(n_2170),
.B(n_2002),
.Y(n_2265)
);

HB1xp67_ASAP7_75t_L g2266 ( 
.A(n_2163),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_2058),
.B(n_47),
.Y(n_2267)
);

AND2x2_ASAP7_75t_L g2268 ( 
.A(n_2057),
.B(n_47),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2153),
.B(n_48),
.Y(n_2269)
);

BUFx3_ASAP7_75t_L g2270 ( 
.A(n_2160),
.Y(n_2270)
);

AND2x4_ASAP7_75t_L g2271 ( 
.A(n_2078),
.B(n_48),
.Y(n_2271)
);

BUFx2_ASAP7_75t_L g2272 ( 
.A(n_2078),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_2085),
.B(n_49),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_2083),
.B(n_50),
.Y(n_2274)
);

OAI22xp5_ASAP7_75t_L g2275 ( 
.A1(n_2060),
.A2(n_1253),
.B1(n_1223),
.B2(n_1271),
.Y(n_2275)
);

AND2x2_ASAP7_75t_L g2276 ( 
.A(n_2096),
.B(n_50),
.Y(n_2276)
);

INVx3_ASAP7_75t_L g2277 ( 
.A(n_2119),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2119),
.Y(n_2278)
);

OR2x2_ASAP7_75t_L g2279 ( 
.A(n_2166),
.B(n_52),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2110),
.B(n_52),
.Y(n_2280)
);

OR2x6_ASAP7_75t_L g2281 ( 
.A(n_2119),
.B(n_1271),
.Y(n_2281)
);

INVx5_ASAP7_75t_L g2282 ( 
.A(n_2156),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2076),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2136),
.B(n_2139),
.Y(n_2284)
);

INVx5_ASAP7_75t_L g2285 ( 
.A(n_2156),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2169),
.Y(n_2286)
);

AND2x4_ASAP7_75t_L g2287 ( 
.A(n_2136),
.B(n_53),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2132),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2102),
.Y(n_2289)
);

NAND2x1_ASAP7_75t_L g2290 ( 
.A(n_2139),
.B(n_1303),
.Y(n_2290)
);

NAND4xp75_ASAP7_75t_L g2291 ( 
.A(n_2080),
.B(n_56),
.C(n_53),
.D(n_55),
.Y(n_2291)
);

OR2x2_ASAP7_75t_L g2292 ( 
.A(n_2166),
.B(n_56),
.Y(n_2292)
);

INVxp67_ASAP7_75t_L g2293 ( 
.A(n_2125),
.Y(n_2293)
);

AND2x4_ASAP7_75t_L g2294 ( 
.A(n_2069),
.B(n_57),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2169),
.Y(n_2295)
);

HB1xp67_ASAP7_75t_L g2296 ( 
.A(n_2195),
.Y(n_2296)
);

NOR2xp33_ASAP7_75t_L g2297 ( 
.A(n_2049),
.B(n_58),
.Y(n_2297)
);

INVxp67_ASAP7_75t_L g2298 ( 
.A(n_2165),
.Y(n_2298)
);

BUFx3_ASAP7_75t_L g2299 ( 
.A(n_2084),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2059),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_2095),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2095),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2095),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2122),
.B(n_58),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_2157),
.Y(n_2305)
);

OAI22xp5_ASAP7_75t_L g2306 ( 
.A1(n_2171),
.A2(n_562),
.B1(n_564),
.B2(n_561),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2150),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_2196),
.B(n_59),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2159),
.Y(n_2309)
);

OR2x2_ASAP7_75t_L g2310 ( 
.A(n_2131),
.B(n_59),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2153),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2148),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2091),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2093),
.Y(n_2314)
);

AND2x2_ASAP7_75t_L g2315 ( 
.A(n_2067),
.B(n_60),
.Y(n_2315)
);

AND2x2_ASAP7_75t_L g2316 ( 
.A(n_2145),
.B(n_62),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2174),
.B(n_2199),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_2101),
.B(n_63),
.Y(n_2318)
);

INVxp67_ASAP7_75t_SL g2319 ( 
.A(n_2201),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_2062),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_2134),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2149),
.Y(n_2322)
);

NAND2xp33_ASAP7_75t_R g2323 ( 
.A(n_2063),
.B(n_63),
.Y(n_2323)
);

OR2x2_ASAP7_75t_L g2324 ( 
.A(n_2144),
.B(n_2120),
.Y(n_2324)
);

NOR2xp33_ASAP7_75t_L g2325 ( 
.A(n_2120),
.B(n_64),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2228),
.B(n_2123),
.Y(n_2326)
);

NOR2xp33_ASAP7_75t_L g2327 ( 
.A(n_2260),
.B(n_2258),
.Y(n_2327)
);

BUFx2_ASAP7_75t_L g2328 ( 
.A(n_2272),
.Y(n_2328)
);

INVxp67_ASAP7_75t_L g2329 ( 
.A(n_2319),
.Y(n_2329)
);

INVx3_ASAP7_75t_L g2330 ( 
.A(n_2270),
.Y(n_2330)
);

AOI21xp5_ASAP7_75t_L g2331 ( 
.A1(n_2269),
.A2(n_2127),
.B(n_2129),
.Y(n_2331)
);

BUFx6f_ASAP7_75t_L g2332 ( 
.A(n_2237),
.Y(n_2332)
);

INVxp67_ASAP7_75t_SL g2333 ( 
.A(n_2311),
.Y(n_2333)
);

AOI21xp5_ASAP7_75t_L g2334 ( 
.A1(n_2324),
.A2(n_2129),
.B(n_2098),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2265),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2265),
.Y(n_2336)
);

BUFx2_ASAP7_75t_L g2337 ( 
.A(n_2272),
.Y(n_2337)
);

INVxp33_ASAP7_75t_L g2338 ( 
.A(n_2231),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2208),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2209),
.Y(n_2340)
);

OR2x2_ASAP7_75t_L g2341 ( 
.A(n_2202),
.B(n_2051),
.Y(n_2341)
);

AOI22xp33_ASAP7_75t_SL g2342 ( 
.A1(n_2318),
.A2(n_2238),
.B1(n_2324),
.B2(n_2304),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_2265),
.Y(n_2343)
);

AOI21xp5_ASAP7_75t_L g2344 ( 
.A1(n_2325),
.A2(n_2126),
.B(n_2114),
.Y(n_2344)
);

AOI22xp33_ASAP7_75t_L g2345 ( 
.A1(n_2304),
.A2(n_2052),
.B1(n_2073),
.B2(n_2055),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2264),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_2264),
.Y(n_2347)
);

INVx1_ASAP7_75t_SL g2348 ( 
.A(n_2239),
.Y(n_2348)
);

O2A1O1Ixp33_ASAP7_75t_L g2349 ( 
.A1(n_2318),
.A2(n_2164),
.B(n_2141),
.C(n_2187),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2212),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2228),
.B(n_2071),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2214),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2226),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2226),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2262),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2262),
.Y(n_2356)
);

A2O1A1Ixp33_ASAP7_75t_L g2357 ( 
.A1(n_2317),
.A2(n_2090),
.B(n_2164),
.C(n_2115),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_2262),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2219),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2242),
.B(n_2124),
.Y(n_2360)
);

OAI22xp33_ASAP7_75t_L g2361 ( 
.A1(n_2309),
.A2(n_2197),
.B1(n_2109),
.B2(n_2179),
.Y(n_2361)
);

O2A1O1Ixp5_ASAP7_75t_L g2362 ( 
.A1(n_2213),
.A2(n_2194),
.B(n_2191),
.C(n_2079),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2223),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2225),
.Y(n_2364)
);

OAI21xp5_ASAP7_75t_L g2365 ( 
.A1(n_2213),
.A2(n_2106),
.B(n_2103),
.Y(n_2365)
);

AOI21xp5_ASAP7_75t_L g2366 ( 
.A1(n_2241),
.A2(n_2117),
.B(n_2097),
.Y(n_2366)
);

AND2x4_ASAP7_75t_L g2367 ( 
.A(n_2277),
.B(n_2198),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2229),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2235),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2203),
.Y(n_2370)
);

AOI22xp5_ASAP7_75t_L g2371 ( 
.A1(n_2313),
.A2(n_2307),
.B1(n_2314),
.B2(n_2296),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2242),
.Y(n_2372)
);

BUFx3_ASAP7_75t_L g2373 ( 
.A(n_2237),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2247),
.Y(n_2374)
);

OAI22xp5_ASAP7_75t_L g2375 ( 
.A1(n_2309),
.A2(n_2298),
.B1(n_2313),
.B2(n_2293),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_2247),
.Y(n_2376)
);

AND2x2_ASAP7_75t_L g2377 ( 
.A(n_2206),
.B(n_2054),
.Y(n_2377)
);

OAI22xp5_ASAP7_75t_L g2378 ( 
.A1(n_2277),
.A2(n_2074),
.B1(n_2176),
.B2(n_2087),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2240),
.Y(n_2379)
);

AND2x2_ASAP7_75t_L g2380 ( 
.A(n_2206),
.B(n_2182),
.Y(n_2380)
);

HB1xp67_ASAP7_75t_L g2381 ( 
.A(n_2230),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2255),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2255),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2243),
.B(n_2181),
.Y(n_2384)
);

AOI22xp33_ASAP7_75t_L g2385 ( 
.A1(n_2314),
.A2(n_2111),
.B1(n_2143),
.B2(n_2086),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_2207),
.Y(n_2386)
);

AND2x4_ASAP7_75t_L g2387 ( 
.A(n_2277),
.B(n_2100),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2243),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2207),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_2207),
.Y(n_2390)
);

AND2x2_ASAP7_75t_L g2391 ( 
.A(n_2266),
.B(n_2184),
.Y(n_2391)
);

AOI22xp5_ASAP7_75t_L g2392 ( 
.A1(n_2307),
.A2(n_2121),
.B1(n_2161),
.B2(n_2130),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2253),
.B(n_2189),
.Y(n_2393)
);

AOI22xp33_ASAP7_75t_L g2394 ( 
.A1(n_2322),
.A2(n_2173),
.B1(n_2167),
.B2(n_2178),
.Y(n_2394)
);

AND2x2_ASAP7_75t_L g2395 ( 
.A(n_2204),
.B(n_2188),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2254),
.Y(n_2396)
);

AND2x2_ASAP7_75t_L g2397 ( 
.A(n_2204),
.B(n_2140),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2216),
.B(n_64),
.Y(n_2398)
);

OAI21xp5_ASAP7_75t_L g2399 ( 
.A1(n_2238),
.A2(n_576),
.B(n_572),
.Y(n_2399)
);

INVx4_ASAP7_75t_L g2400 ( 
.A(n_2270),
.Y(n_2400)
);

CKINVDCx5p33_ASAP7_75t_R g2401 ( 
.A(n_2299),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2250),
.B(n_65),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_2217),
.Y(n_2403)
);

INVxp67_ASAP7_75t_L g2404 ( 
.A(n_2257),
.Y(n_2404)
);

AOI22xp33_ASAP7_75t_L g2405 ( 
.A1(n_2322),
.A2(n_579),
.B1(n_580),
.B2(n_578),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2224),
.Y(n_2406)
);

BUFx6f_ASAP7_75t_L g2407 ( 
.A(n_2271),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2224),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_2217),
.Y(n_2409)
);

AOI21xp5_ASAP7_75t_L g2410 ( 
.A1(n_2245),
.A2(n_66),
.B(n_67),
.Y(n_2410)
);

INVx2_ASAP7_75t_L g2411 ( 
.A(n_2217),
.Y(n_2411)
);

AOI22xp33_ASAP7_75t_L g2412 ( 
.A1(n_2320),
.A2(n_586),
.B1(n_596),
.B2(n_583),
.Y(n_2412)
);

AND2x4_ASAP7_75t_L g2413 ( 
.A(n_2216),
.B(n_66),
.Y(n_2413)
);

HB1xp67_ASAP7_75t_L g2414 ( 
.A(n_2233),
.Y(n_2414)
);

INVx3_ASAP7_75t_L g2415 ( 
.A(n_2282),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2249),
.B(n_67),
.Y(n_2416)
);

OR2x2_ASAP7_75t_L g2417 ( 
.A(n_2321),
.B(n_68),
.Y(n_2417)
);

AND2x2_ASAP7_75t_L g2418 ( 
.A(n_2218),
.B(n_2221),
.Y(n_2418)
);

OAI22xp33_ASAP7_75t_L g2419 ( 
.A1(n_2323),
.A2(n_598),
.B1(n_608),
.B2(n_597),
.Y(n_2419)
);

OAI21xp5_ASAP7_75t_L g2420 ( 
.A1(n_2267),
.A2(n_619),
.B(n_614),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2210),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2321),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2259),
.Y(n_2423)
);

OR2x2_ASAP7_75t_L g2424 ( 
.A(n_2312),
.B(n_68),
.Y(n_2424)
);

BUFx6f_ASAP7_75t_SL g2425 ( 
.A(n_2271),
.Y(n_2425)
);

BUFx12f_ASAP7_75t_L g2426 ( 
.A(n_2294),
.Y(n_2426)
);

OA21x2_ASAP7_75t_L g2427 ( 
.A1(n_2234),
.A2(n_1030),
.B(n_1029),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2261),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2305),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_2210),
.Y(n_2430)
);

AND2x2_ASAP7_75t_L g2431 ( 
.A(n_2218),
.B(n_69),
.Y(n_2431)
);

BUFx5_ASAP7_75t_L g2432 ( 
.A(n_2271),
.Y(n_2432)
);

AND2x2_ASAP7_75t_L g2433 ( 
.A(n_2221),
.B(n_69),
.Y(n_2433)
);

AOI22xp5_ASAP7_75t_L g2434 ( 
.A1(n_2320),
.A2(n_631),
.B1(n_637),
.B2(n_621),
.Y(n_2434)
);

NAND3xp33_ASAP7_75t_L g2435 ( 
.A(n_2244),
.B(n_1030),
.C(n_1029),
.Y(n_2435)
);

AOI221xp5_ASAP7_75t_L g2436 ( 
.A1(n_2244),
.A2(n_640),
.B1(n_646),
.B2(n_655),
.C(n_661),
.Y(n_2436)
);

O2A1O1Ixp5_ASAP7_75t_L g2437 ( 
.A1(n_2267),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_2437)
);

OAI21xp5_ASAP7_75t_L g2438 ( 
.A1(n_2273),
.A2(n_665),
.B(n_662),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2339),
.Y(n_2439)
);

OAI33xp33_ASAP7_75t_L g2440 ( 
.A1(n_2329),
.A2(n_2283),
.A3(n_2300),
.B1(n_2263),
.B2(n_2295),
.B3(n_2288),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_2432),
.Y(n_2441)
);

NAND3xp33_ASAP7_75t_SL g2442 ( 
.A(n_2342),
.B(n_2268),
.C(n_2273),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2432),
.Y(n_2443)
);

AND2x2_ASAP7_75t_L g2444 ( 
.A(n_2330),
.B(n_2248),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2340),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2350),
.Y(n_2446)
);

BUFx2_ASAP7_75t_L g2447 ( 
.A(n_2426),
.Y(n_2447)
);

CKINVDCx5p33_ASAP7_75t_R g2448 ( 
.A(n_2401),
.Y(n_2448)
);

INVx1_ASAP7_75t_SL g2449 ( 
.A(n_2373),
.Y(n_2449)
);

AOI221xp5_ASAP7_75t_L g2450 ( 
.A1(n_2331),
.A2(n_2342),
.B1(n_2329),
.B2(n_2334),
.C(n_2361),
.Y(n_2450)
);

AND2x2_ASAP7_75t_L g2451 ( 
.A(n_2330),
.B(n_2248),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2352),
.Y(n_2452)
);

AND2x2_ASAP7_75t_L g2453 ( 
.A(n_2326),
.B(n_2205),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2359),
.Y(n_2454)
);

HB1xp67_ASAP7_75t_L g2455 ( 
.A(n_2388),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_2400),
.B(n_2227),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_2418),
.B(n_2205),
.Y(n_2457)
);

OR2x2_ASAP7_75t_L g2458 ( 
.A(n_2341),
.B(n_2305),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_2400),
.B(n_2284),
.Y(n_2459)
);

AND2x4_ASAP7_75t_L g2460 ( 
.A(n_2328),
.B(n_2282),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2327),
.B(n_2284),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2331),
.B(n_2274),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_2432),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2432),
.Y(n_2464)
);

AND2x4_ASAP7_75t_L g2465 ( 
.A(n_2337),
.B(n_2282),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_2432),
.Y(n_2466)
);

AND2x4_ASAP7_75t_L g2467 ( 
.A(n_2335),
.B(n_2282),
.Y(n_2467)
);

OR2x2_ASAP7_75t_L g2468 ( 
.A(n_2416),
.B(n_2312),
.Y(n_2468)
);

OR2x2_ASAP7_75t_L g2469 ( 
.A(n_2416),
.B(n_2249),
.Y(n_2469)
);

AND2x2_ASAP7_75t_L g2470 ( 
.A(n_2327),
.B(n_2268),
.Y(n_2470)
);

AND2x4_ASAP7_75t_L g2471 ( 
.A(n_2336),
.B(n_2282),
.Y(n_2471)
);

INVx4_ASAP7_75t_L g2472 ( 
.A(n_2332),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2363),
.Y(n_2473)
);

AND2x2_ASAP7_75t_L g2474 ( 
.A(n_2333),
.B(n_2395),
.Y(n_2474)
);

OAI21x1_ASAP7_75t_L g2475 ( 
.A1(n_2386),
.A2(n_2300),
.B(n_2233),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2364),
.Y(n_2476)
);

HB1xp67_ASAP7_75t_L g2477 ( 
.A(n_2370),
.Y(n_2477)
);

OAI222xp33_ASAP7_75t_L g2478 ( 
.A1(n_2371),
.A2(n_2279),
.B1(n_2292),
.B2(n_2286),
.C1(n_2215),
.C2(n_2251),
.Y(n_2478)
);

INVx4_ASAP7_75t_L g2479 ( 
.A(n_2332),
.Y(n_2479)
);

AOI22xp33_ASAP7_75t_L g2480 ( 
.A1(n_2334),
.A2(n_2279),
.B1(n_2292),
.B2(n_2286),
.Y(n_2480)
);

AND2x4_ASAP7_75t_L g2481 ( 
.A(n_2343),
.B(n_2285),
.Y(n_2481)
);

HB1xp67_ASAP7_75t_L g2482 ( 
.A(n_2396),
.Y(n_2482)
);

INVx5_ASAP7_75t_L g2483 ( 
.A(n_2332),
.Y(n_2483)
);

AOI22xp33_ASAP7_75t_L g2484 ( 
.A1(n_2384),
.A2(n_2256),
.B1(n_2308),
.B2(n_2276),
.Y(n_2484)
);

AND2x2_ASAP7_75t_L g2485 ( 
.A(n_2380),
.B(n_2251),
.Y(n_2485)
);

OA21x2_ASAP7_75t_L g2486 ( 
.A1(n_2333),
.A2(n_2215),
.B(n_2252),
.Y(n_2486)
);

BUFx2_ASAP7_75t_L g2487 ( 
.A(n_2332),
.Y(n_2487)
);

HB1xp67_ASAP7_75t_L g2488 ( 
.A(n_2346),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2432),
.Y(n_2489)
);

INVxp67_ASAP7_75t_L g2490 ( 
.A(n_2425),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2436),
.B(n_2274),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2368),
.Y(n_2492)
);

AND2x4_ASAP7_75t_L g2493 ( 
.A(n_2407),
.B(n_2285),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2436),
.B(n_2276),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2410),
.B(n_2280),
.Y(n_2495)
);

INVx3_ASAP7_75t_L g2496 ( 
.A(n_2407),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2369),
.Y(n_2497)
);

NOR2xp67_ASAP7_75t_SL g2498 ( 
.A(n_2407),
.B(n_2299),
.Y(n_2498)
);

AO21x2_ASAP7_75t_L g2499 ( 
.A1(n_2384),
.A2(n_2297),
.B(n_2280),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_2397),
.B(n_2294),
.Y(n_2500)
);

OR2x2_ASAP7_75t_L g2501 ( 
.A(n_2393),
.B(n_2278),
.Y(n_2501)
);

INVx5_ASAP7_75t_L g2502 ( 
.A(n_2415),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2407),
.Y(n_2503)
);

AOI221xp5_ASAP7_75t_L g2504 ( 
.A1(n_2361),
.A2(n_2236),
.B1(n_2289),
.B2(n_2232),
.C(n_2315),
.Y(n_2504)
);

OR2x2_ASAP7_75t_L g2505 ( 
.A(n_2393),
.B(n_2246),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2374),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2410),
.B(n_2294),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2402),
.B(n_2429),
.Y(n_2508)
);

NAND2x1p5_ASAP7_75t_SL g2509 ( 
.A(n_2398),
.B(n_2315),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2424),
.Y(n_2510)
);

OR2x6_ASAP7_75t_L g2511 ( 
.A(n_2399),
.B(n_2287),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2417),
.Y(n_2512)
);

INVxp67_ASAP7_75t_L g2513 ( 
.A(n_2425),
.Y(n_2513)
);

AND2x4_ASAP7_75t_L g2514 ( 
.A(n_2415),
.B(n_2285),
.Y(n_2514)
);

HB1xp67_ASAP7_75t_L g2515 ( 
.A(n_2347),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2355),
.Y(n_2516)
);

AND2x2_ASAP7_75t_L g2517 ( 
.A(n_2338),
.B(n_2414),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_2356),
.Y(n_2518)
);

HB1xp67_ASAP7_75t_L g2519 ( 
.A(n_2414),
.Y(n_2519)
);

OR2x2_ASAP7_75t_L g2520 ( 
.A(n_2402),
.B(n_2246),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2423),
.Y(n_2521)
);

INVx3_ASAP7_75t_L g2522 ( 
.A(n_2413),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2428),
.Y(n_2523)
);

OAI21xp5_ASAP7_75t_L g2524 ( 
.A1(n_2362),
.A2(n_2287),
.B(n_2291),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2351),
.B(n_2232),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2358),
.Y(n_2526)
);

HB1xp67_ASAP7_75t_L g2527 ( 
.A(n_2519),
.Y(n_2527)
);

BUFx3_ASAP7_75t_L g2528 ( 
.A(n_2448),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2519),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2462),
.B(n_2375),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2474),
.B(n_2391),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2486),
.Y(n_2532)
);

HB1xp67_ASAP7_75t_L g2533 ( 
.A(n_2517),
.Y(n_2533)
);

INVxp67_ASAP7_75t_L g2534 ( 
.A(n_2456),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2486),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2474),
.B(n_2377),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_2499),
.B(n_2431),
.Y(n_2537)
);

INVx2_ASAP7_75t_SL g2538 ( 
.A(n_2483),
.Y(n_2538)
);

NOR2xp67_ASAP7_75t_L g2539 ( 
.A(n_2483),
.B(n_2285),
.Y(n_2539)
);

NAND2xp33_ASAP7_75t_SL g2540 ( 
.A(n_2498),
.B(n_2338),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2470),
.B(n_2389),
.Y(n_2541)
);

AND2x2_ASAP7_75t_L g2542 ( 
.A(n_2461),
.B(n_2390),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2455),
.Y(n_2543)
);

INVxp67_ASAP7_75t_L g2544 ( 
.A(n_2456),
.Y(n_2544)
);

OR2x2_ASAP7_75t_L g2545 ( 
.A(n_2442),
.B(n_2372),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2455),
.Y(n_2546)
);

INVx3_ASAP7_75t_L g2547 ( 
.A(n_2486),
.Y(n_2547)
);

OR2x2_ASAP7_75t_L g2548 ( 
.A(n_2477),
.B(n_2379),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_2522),
.B(n_2403),
.Y(n_2549)
);

AND2x2_ASAP7_75t_L g2550 ( 
.A(n_2522),
.B(n_2409),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2509),
.Y(n_2551)
);

OAI21xp5_ASAP7_75t_L g2552 ( 
.A1(n_2450),
.A2(n_2362),
.B(n_2437),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2499),
.B(n_2433),
.Y(n_2553)
);

OR2x2_ASAP7_75t_L g2554 ( 
.A(n_2477),
.B(n_2381),
.Y(n_2554)
);

BUFx2_ASAP7_75t_L g2555 ( 
.A(n_2447),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2482),
.Y(n_2556)
);

AND2x2_ASAP7_75t_L g2557 ( 
.A(n_2522),
.B(n_2453),
.Y(n_2557)
);

AND2x4_ASAP7_75t_L g2558 ( 
.A(n_2483),
.B(n_2411),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2482),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2509),
.Y(n_2560)
);

INVx3_ASAP7_75t_L g2561 ( 
.A(n_2472),
.Y(n_2561)
);

OR2x2_ASAP7_75t_L g2562 ( 
.A(n_2508),
.B(n_2381),
.Y(n_2562)
);

AND2x2_ASAP7_75t_L g2563 ( 
.A(n_2487),
.B(n_2413),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2521),
.Y(n_2564)
);

OR2x2_ASAP7_75t_L g2565 ( 
.A(n_2469),
.B(n_2360),
.Y(n_2565)
);

AND2x4_ASAP7_75t_L g2566 ( 
.A(n_2483),
.B(n_2353),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2496),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2523),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2496),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2496),
.Y(n_2570)
);

INVx3_ASAP7_75t_L g2571 ( 
.A(n_2472),
.Y(n_2571)
);

CKINVDCx16_ASAP7_75t_R g2572 ( 
.A(n_2524),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2439),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2445),
.Y(n_2574)
);

AND3x1_ASAP7_75t_L g2575 ( 
.A(n_2504),
.B(n_2438),
.C(n_2349),
.Y(n_2575)
);

AND2x2_ASAP7_75t_L g2576 ( 
.A(n_2500),
.B(n_2459),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2457),
.B(n_2348),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2446),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2457),
.B(n_2493),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_L g2580 ( 
.A(n_2495),
.B(n_2344),
.Y(n_2580)
);

AND2x2_ASAP7_75t_L g2581 ( 
.A(n_2493),
.B(n_2236),
.Y(n_2581)
);

NOR2xp33_ASAP7_75t_L g2582 ( 
.A(n_2448),
.B(n_2419),
.Y(n_2582)
);

HB1xp67_ASAP7_75t_L g2583 ( 
.A(n_2517),
.Y(n_2583)
);

NAND2x1p5_ASAP7_75t_L g2584 ( 
.A(n_2472),
.B(n_2287),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2503),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2468),
.B(n_2344),
.Y(n_2586)
);

BUFx3_ASAP7_75t_L g2587 ( 
.A(n_2479),
.Y(n_2587)
);

AND2x2_ASAP7_75t_L g2588 ( 
.A(n_2493),
.B(n_2444),
.Y(n_2588)
);

INVx2_ASAP7_75t_L g2589 ( 
.A(n_2503),
.Y(n_2589)
);

NOR2xp33_ASAP7_75t_L g2590 ( 
.A(n_2449),
.B(n_2419),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2491),
.B(n_2367),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2452),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2510),
.Y(n_2593)
);

HB1xp67_ASAP7_75t_L g2594 ( 
.A(n_2501),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_2510),
.Y(n_2595)
);

INVx2_ASAP7_75t_L g2596 ( 
.A(n_2475),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2454),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_2475),
.Y(n_2598)
);

AND2x2_ASAP7_75t_L g2599 ( 
.A(n_2451),
.B(n_2367),
.Y(n_2599)
);

OR2x2_ASAP7_75t_L g2600 ( 
.A(n_2506),
.B(n_2360),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2512),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2473),
.Y(n_2602)
);

BUFx2_ASAP7_75t_L g2603 ( 
.A(n_2479),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2512),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2525),
.B(n_2354),
.Y(n_2605)
);

BUFx2_ASAP7_75t_L g2606 ( 
.A(n_2479),
.Y(n_2606)
);

HB1xp67_ASAP7_75t_L g2607 ( 
.A(n_2490),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2476),
.Y(n_2608)
);

XOR2x2_ASAP7_75t_L g2609 ( 
.A(n_2575),
.B(n_2494),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2527),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2547),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2533),
.Y(n_2612)
);

NOR3xp33_ASAP7_75t_SL g2613 ( 
.A(n_2572),
.B(n_2540),
.C(n_2552),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2583),
.Y(n_2614)
);

INVx2_ASAP7_75t_SL g2615 ( 
.A(n_2528),
.Y(n_2615)
);

XOR2x2_ASAP7_75t_L g2616 ( 
.A(n_2575),
.B(n_2507),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2547),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_2572),
.B(n_2492),
.Y(n_2618)
);

NAND3xp33_ASAP7_75t_L g2619 ( 
.A(n_2580),
.B(n_2437),
.C(n_2513),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2529),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2577),
.B(n_2485),
.Y(n_2621)
);

AND2x2_ASAP7_75t_L g2622 ( 
.A(n_2577),
.B(n_2460),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2547),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2551),
.B(n_2497),
.Y(n_2624)
);

AOI22xp5_ASAP7_75t_L g2625 ( 
.A1(n_2551),
.A2(n_2440),
.B1(n_2480),
.B2(n_2484),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2529),
.Y(n_2626)
);

NAND4xp75_ASAP7_75t_SL g2627 ( 
.A(n_2539),
.B(n_2427),
.C(n_2502),
.D(n_2465),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2543),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2532),
.Y(n_2629)
);

AND2x2_ASAP7_75t_L g2630 ( 
.A(n_2579),
.B(n_2460),
.Y(n_2630)
);

AND2x2_ASAP7_75t_L g2631 ( 
.A(n_2579),
.B(n_2460),
.Y(n_2631)
);

OAI21xp5_ASAP7_75t_SL g2632 ( 
.A1(n_2560),
.A2(n_2478),
.B(n_2349),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2543),
.Y(n_2633)
);

XOR2x2_ASAP7_75t_L g2634 ( 
.A(n_2530),
.B(n_2484),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2546),
.Y(n_2635)
);

NAND4xp75_ASAP7_75t_L g2636 ( 
.A(n_2560),
.B(n_2366),
.C(n_2443),
.D(n_2441),
.Y(n_2636)
);

XNOR2xp5_ASAP7_75t_L g2637 ( 
.A(n_2528),
.B(n_2345),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2532),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_L g2639 ( 
.A(n_2594),
.B(n_2480),
.Y(n_2639)
);

INVxp67_ASAP7_75t_SL g2640 ( 
.A(n_2535),
.Y(n_2640)
);

OR2x2_ASAP7_75t_L g2641 ( 
.A(n_2536),
.B(n_2520),
.Y(n_2641)
);

AND2x2_ASAP7_75t_L g2642 ( 
.A(n_2555),
.B(n_2465),
.Y(n_2642)
);

AND2x2_ASAP7_75t_L g2643 ( 
.A(n_2555),
.B(n_2465),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2586),
.B(n_2488),
.Y(n_2644)
);

OAI22xp5_ASAP7_75t_L g2645 ( 
.A1(n_2545),
.A2(n_2511),
.B1(n_2345),
.B2(n_2394),
.Y(n_2645)
);

XNOR2xp5_ASAP7_75t_L g2646 ( 
.A(n_2528),
.B(n_2599),
.Y(n_2646)
);

XNOR2xp5_ASAP7_75t_L g2647 ( 
.A(n_2599),
.B(n_2392),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2546),
.Y(n_2648)
);

AND2x2_ASAP7_75t_L g2649 ( 
.A(n_2576),
.B(n_2514),
.Y(n_2649)
);

NOR4xp25_ASAP7_75t_L g2650 ( 
.A(n_2534),
.B(n_2544),
.C(n_2553),
.D(n_2537),
.Y(n_2650)
);

AND2x2_ASAP7_75t_L g2651 ( 
.A(n_2576),
.B(n_2514),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2556),
.Y(n_2652)
);

NAND3xp33_ASAP7_75t_SL g2653 ( 
.A(n_2545),
.B(n_2420),
.C(n_2405),
.Y(n_2653)
);

XOR2x2_ASAP7_75t_L g2654 ( 
.A(n_2591),
.B(n_2582),
.Y(n_2654)
);

INVx2_ASAP7_75t_SL g2655 ( 
.A(n_2563),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_L g2656 ( 
.A(n_2565),
.B(n_2488),
.Y(n_2656)
);

NAND4xp75_ASAP7_75t_L g2657 ( 
.A(n_2539),
.B(n_2366),
.C(n_2443),
.D(n_2441),
.Y(n_2657)
);

NAND4xp75_ASAP7_75t_L g2658 ( 
.A(n_2535),
.B(n_2464),
.C(n_2466),
.D(n_2463),
.Y(n_2658)
);

NOR4xp25_ASAP7_75t_L g2659 ( 
.A(n_2556),
.B(n_2463),
.C(n_2466),
.D(n_2464),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2559),
.Y(n_2660)
);

AND2x2_ASAP7_75t_L g2661 ( 
.A(n_2563),
.B(n_2514),
.Y(n_2661)
);

NOR2x1_ASAP7_75t_L g2662 ( 
.A(n_2587),
.B(n_2489),
.Y(n_2662)
);

INVx2_ASAP7_75t_SL g2663 ( 
.A(n_2588),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2559),
.Y(n_2664)
);

NAND4xp75_ASAP7_75t_L g2665 ( 
.A(n_2557),
.B(n_2489),
.C(n_2365),
.D(n_2516),
.Y(n_2665)
);

BUFx3_ASAP7_75t_L g2666 ( 
.A(n_2587),
.Y(n_2666)
);

BUFx2_ASAP7_75t_L g2667 ( 
.A(n_2584),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2565),
.B(n_2515),
.Y(n_2668)
);

INVxp67_ASAP7_75t_SL g2669 ( 
.A(n_2590),
.Y(n_2669)
);

XNOR2x1_ASAP7_75t_L g2670 ( 
.A(n_2584),
.B(n_2511),
.Y(n_2670)
);

AOI22xp5_ASAP7_75t_L g2671 ( 
.A1(n_2616),
.A2(n_2598),
.B1(n_2596),
.B2(n_2511),
.Y(n_2671)
);

INVx2_ASAP7_75t_SL g2672 ( 
.A(n_2642),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2637),
.B(n_2557),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2640),
.Y(n_2674)
);

AND2x2_ASAP7_75t_L g2675 ( 
.A(n_2621),
.B(n_2588),
.Y(n_2675)
);

INVx2_ASAP7_75t_SL g2676 ( 
.A(n_2643),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2655),
.B(n_2607),
.Y(n_2677)
);

AND2x2_ASAP7_75t_L g2678 ( 
.A(n_2622),
.B(n_2584),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2609),
.Y(n_2679)
);

AND2x2_ASAP7_75t_L g2680 ( 
.A(n_2649),
.B(n_2541),
.Y(n_2680)
);

AND2x2_ASAP7_75t_L g2681 ( 
.A(n_2651),
.B(n_2541),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2640),
.Y(n_2682)
);

NAND2x1p5_ASAP7_75t_L g2683 ( 
.A(n_2666),
.B(n_2587),
.Y(n_2683)
);

AND2x2_ASAP7_75t_L g2684 ( 
.A(n_2613),
.B(n_2542),
.Y(n_2684)
);

AND2x4_ASAP7_75t_L g2685 ( 
.A(n_2661),
.B(n_2603),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2634),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2639),
.Y(n_2687)
);

AND2x2_ASAP7_75t_L g2688 ( 
.A(n_2613),
.B(n_2542),
.Y(n_2688)
);

AND2x2_ASAP7_75t_L g2689 ( 
.A(n_2630),
.B(n_2631),
.Y(n_2689)
);

OAI211xp5_ASAP7_75t_L g2690 ( 
.A1(n_2650),
.A2(n_2554),
.B(n_2606),
.C(n_2603),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2611),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2615),
.B(n_2531),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2611),
.Y(n_2693)
);

AOI22xp5_ASAP7_75t_L g2694 ( 
.A1(n_2625),
.A2(n_2598),
.B1(n_2596),
.B2(n_2511),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2663),
.B(n_2549),
.Y(n_2695)
);

INVx2_ASAP7_75t_L g2696 ( 
.A(n_2617),
.Y(n_2696)
);

AND2x2_ASAP7_75t_L g2697 ( 
.A(n_2646),
.B(n_2549),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2667),
.B(n_2550),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2617),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2623),
.Y(n_2700)
);

INVx2_ASAP7_75t_SL g2701 ( 
.A(n_2670),
.Y(n_2701)
);

NOR2x1_ASAP7_75t_L g2702 ( 
.A(n_2666),
.B(n_2606),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2623),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2656),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2656),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2668),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2647),
.B(n_2605),
.Y(n_2707)
);

OAI21xp5_ASAP7_75t_L g2708 ( 
.A1(n_2632),
.A2(n_2554),
.B(n_2600),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2668),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2639),
.Y(n_2710)
);

AND2x2_ASAP7_75t_L g2711 ( 
.A(n_2612),
.B(n_2550),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2629),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2629),
.Y(n_2713)
);

AND2x2_ASAP7_75t_L g2714 ( 
.A(n_2614),
.B(n_2538),
.Y(n_2714)
);

NOR2xp33_ASAP7_75t_L g2715 ( 
.A(n_2653),
.B(n_2600),
.Y(n_2715)
);

NOR3xp33_ASAP7_75t_L g2716 ( 
.A(n_2653),
.B(n_2538),
.C(n_2561),
.Y(n_2716)
);

AND2x2_ASAP7_75t_L g2717 ( 
.A(n_2641),
.B(n_2605),
.Y(n_2717)
);

OAI22xp5_ASAP7_75t_L g2718 ( 
.A1(n_2673),
.A2(n_2636),
.B1(n_2665),
.B2(n_2619),
.Y(n_2718)
);

O2A1O1Ixp33_ASAP7_75t_L g2719 ( 
.A1(n_2715),
.A2(n_2645),
.B(n_2669),
.C(n_2644),
.Y(n_2719)
);

AOI22xp5_ASAP7_75t_L g2720 ( 
.A1(n_2679),
.A2(n_2645),
.B1(n_2669),
.B2(n_2654),
.Y(n_2720)
);

NAND4xp25_ASAP7_75t_L g2721 ( 
.A(n_2684),
.B(n_2610),
.C(n_2618),
.D(n_2620),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2717),
.Y(n_2722)
);

INVx2_ASAP7_75t_L g2723 ( 
.A(n_2675),
.Y(n_2723)
);

OAI22xp33_ASAP7_75t_L g2724 ( 
.A1(n_2687),
.A2(n_2710),
.B1(n_2708),
.B2(n_2694),
.Y(n_2724)
);

OAI221xp5_ASAP7_75t_L g2725 ( 
.A1(n_2687),
.A2(n_2618),
.B1(n_2644),
.B2(n_2659),
.C(n_2624),
.Y(n_2725)
);

OAI21xp33_ASAP7_75t_L g2726 ( 
.A1(n_2675),
.A2(n_2624),
.B(n_2581),
.Y(n_2726)
);

NOR2xp67_ASAP7_75t_L g2727 ( 
.A(n_2672),
.B(n_2561),
.Y(n_2727)
);

OAI21xp5_ASAP7_75t_L g2728 ( 
.A1(n_2684),
.A2(n_2657),
.B(n_2658),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2717),
.Y(n_2729)
);

OAI221xp5_ASAP7_75t_L g2730 ( 
.A1(n_2710),
.A2(n_2638),
.B1(n_2562),
.B2(n_2458),
.C(n_2589),
.Y(n_2730)
);

AOI22xp33_ASAP7_75t_L g2731 ( 
.A1(n_2679),
.A2(n_2638),
.B1(n_2593),
.B2(n_2601),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2674),
.Y(n_2732)
);

OAI21xp5_ASAP7_75t_L g2733 ( 
.A1(n_2690),
.A2(n_2626),
.B(n_2664),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2682),
.Y(n_2734)
);

XNOR2x2_ASAP7_75t_L g2735 ( 
.A(n_2702),
.B(n_2628),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2696),
.Y(n_2736)
);

AOI22xp33_ASAP7_75t_L g2737 ( 
.A1(n_2686),
.A2(n_2593),
.B1(n_2601),
.B2(n_2595),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2696),
.Y(n_2738)
);

NOR2xp33_ASAP7_75t_L g2739 ( 
.A(n_2685),
.B(n_2562),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2711),
.Y(n_2740)
);

OAI22xp5_ASAP7_75t_L g2741 ( 
.A1(n_2688),
.A2(n_2672),
.B1(n_2676),
.B2(n_2697),
.Y(n_2741)
);

AO22x1_ASAP7_75t_L g2742 ( 
.A1(n_2688),
.A2(n_2697),
.B1(n_2685),
.B2(n_2676),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2711),
.Y(n_2743)
);

AOI22xp5_ASAP7_75t_L g2744 ( 
.A1(n_2686),
.A2(n_2604),
.B1(n_2595),
.B2(n_2434),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2712),
.Y(n_2745)
);

AOI21xp33_ASAP7_75t_L g2746 ( 
.A1(n_2707),
.A2(n_2604),
.B(n_2589),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2713),
.Y(n_2747)
);

OAI21xp33_ASAP7_75t_L g2748 ( 
.A1(n_2680),
.A2(n_2581),
.B(n_2585),
.Y(n_2748)
);

OAI21xp33_ASAP7_75t_SL g2749 ( 
.A1(n_2680),
.A2(n_2627),
.B(n_2548),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2681),
.B(n_2564),
.Y(n_2750)
);

AOI21xp5_ASAP7_75t_L g2751 ( 
.A1(n_2677),
.A2(n_2548),
.B(n_2566),
.Y(n_2751)
);

OAI21xp5_ASAP7_75t_L g2752 ( 
.A1(n_2698),
.A2(n_2566),
.B(n_2662),
.Y(n_2752)
);

AOI221xp5_ASAP7_75t_L g2753 ( 
.A1(n_2671),
.A2(n_2648),
.B1(n_2652),
.B2(n_2635),
.C(n_2633),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2681),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2695),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2723),
.Y(n_2756)
);

NOR2xp33_ASAP7_75t_L g2757 ( 
.A(n_2726),
.B(n_2685),
.Y(n_2757)
);

OAI21xp33_ASAP7_75t_L g2758 ( 
.A1(n_2754),
.A2(n_2689),
.B(n_2678),
.Y(n_2758)
);

NOR2xp33_ASAP7_75t_L g2759 ( 
.A(n_2748),
.B(n_2689),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2722),
.Y(n_2760)
);

OAI22xp33_ASAP7_75t_L g2761 ( 
.A1(n_2720),
.A2(n_2701),
.B1(n_2505),
.B2(n_2693),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2739),
.B(n_2695),
.Y(n_2762)
);

INVx1_ASAP7_75t_SL g2763 ( 
.A(n_2729),
.Y(n_2763)
);

AOI332xp33_ASAP7_75t_L g2764 ( 
.A1(n_2740),
.A2(n_2704),
.A3(n_2705),
.B1(n_2709),
.B2(n_2706),
.B3(n_2691),
.C1(n_2703),
.C2(n_2699),
.Y(n_2764)
);

INVxp67_ASAP7_75t_SL g2765 ( 
.A(n_2735),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2742),
.B(n_2698),
.Y(n_2766)
);

AOI222xp33_ASAP7_75t_L g2767 ( 
.A1(n_2725),
.A2(n_2700),
.B1(n_2660),
.B2(n_2701),
.C1(n_2564),
.C2(n_2578),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2743),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2750),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2755),
.Y(n_2770)
);

AOI221xp5_ASAP7_75t_L g2771 ( 
.A1(n_2724),
.A2(n_2716),
.B1(n_2574),
.B2(n_2578),
.C(n_2573),
.Y(n_2771)
);

OR2x2_ASAP7_75t_L g2772 ( 
.A(n_2721),
.B(n_2692),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2736),
.Y(n_2773)
);

AOI211xp5_ASAP7_75t_SL g2774 ( 
.A1(n_2741),
.A2(n_2714),
.B(n_2561),
.C(n_2571),
.Y(n_2774)
);

AOI22xp33_ASAP7_75t_L g2775 ( 
.A1(n_2718),
.A2(n_2516),
.B1(n_2526),
.B2(n_2518),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2738),
.Y(n_2776)
);

AOI311xp33_ASAP7_75t_L g2777 ( 
.A1(n_2733),
.A2(n_2568),
.A3(n_2592),
.B(n_2574),
.C(n_2573),
.Y(n_2777)
);

NOR2xp33_ASAP7_75t_SL g2778 ( 
.A(n_2719),
.B(n_2683),
.Y(n_2778)
);

AOI322xp5_ASAP7_75t_L g2779 ( 
.A1(n_2731),
.A2(n_2714),
.A3(n_2678),
.B1(n_2597),
.B2(n_2592),
.C1(n_2608),
.C2(n_2602),
.Y(n_2779)
);

OAI21xp5_ASAP7_75t_L g2780 ( 
.A1(n_2749),
.A2(n_2683),
.B(n_2566),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_SL g2781 ( 
.A(n_2727),
.B(n_2502),
.Y(n_2781)
);

O2A1O1Ixp33_ASAP7_75t_L g2782 ( 
.A1(n_2733),
.A2(n_2683),
.B(n_2568),
.C(n_2602),
.Y(n_2782)
);

OA21x2_ASAP7_75t_L g2783 ( 
.A1(n_2728),
.A2(n_2585),
.B(n_2569),
.Y(n_2783)
);

AOI221xp5_ASAP7_75t_SL g2784 ( 
.A1(n_2721),
.A2(n_2608),
.B1(n_2597),
.B2(n_2569),
.C(n_2570),
.Y(n_2784)
);

AND2x2_ASAP7_75t_L g2785 ( 
.A(n_2752),
.B(n_2571),
.Y(n_2785)
);

OR2x2_ASAP7_75t_L g2786 ( 
.A(n_2745),
.B(n_2571),
.Y(n_2786)
);

OR2x2_ASAP7_75t_L g2787 ( 
.A(n_2747),
.B(n_2567),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2765),
.B(n_2751),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2762),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2763),
.B(n_2759),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2782),
.Y(n_2791)
);

A2O1A1Ixp33_ASAP7_75t_L g2792 ( 
.A1(n_2778),
.A2(n_2730),
.B(n_2746),
.C(n_2753),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2758),
.B(n_2732),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2756),
.Y(n_2794)
);

OR2x2_ASAP7_75t_L g2795 ( 
.A(n_2772),
.B(n_2734),
.Y(n_2795)
);

OAI221xp5_ASAP7_75t_L g2796 ( 
.A1(n_2767),
.A2(n_2737),
.B1(n_2744),
.B2(n_2570),
.C(n_2567),
.Y(n_2796)
);

OAI21xp5_ASAP7_75t_SL g2797 ( 
.A1(n_2774),
.A2(n_2566),
.B(n_2558),
.Y(n_2797)
);

OAI21xp33_ASAP7_75t_SL g2798 ( 
.A1(n_2779),
.A2(n_2627),
.B(n_2515),
.Y(n_2798)
);

NOR2xp33_ASAP7_75t_L g2799 ( 
.A(n_2778),
.B(n_2558),
.Y(n_2799)
);

INVx2_ASAP7_75t_L g2800 ( 
.A(n_2783),
.Y(n_2800)
);

NAND3xp33_ASAP7_75t_L g2801 ( 
.A(n_2777),
.B(n_2412),
.C(n_2405),
.Y(n_2801)
);

OAI32xp33_ASAP7_75t_L g2802 ( 
.A1(n_2766),
.A2(n_2757),
.A3(n_2780),
.B1(n_2760),
.B2(n_2770),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2787),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2769),
.B(n_2518),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2785),
.B(n_2558),
.Y(n_2805)
);

AOI22xp5_ASAP7_75t_L g2806 ( 
.A1(n_2761),
.A2(n_2526),
.B1(n_2558),
.B2(n_2471),
.Y(n_2806)
);

OR2x2_ASAP7_75t_L g2807 ( 
.A(n_2768),
.B(n_2467),
.Y(n_2807)
);

INVxp67_ASAP7_75t_L g2808 ( 
.A(n_2781),
.Y(n_2808)
);

NAND3xp33_ASAP7_75t_L g2809 ( 
.A(n_2771),
.B(n_2412),
.C(n_2502),
.Y(n_2809)
);

INVx1_ASAP7_75t_SL g2810 ( 
.A(n_2783),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_SL g2811 ( 
.A(n_2784),
.B(n_2502),
.Y(n_2811)
);

OR2x2_ASAP7_75t_L g2812 ( 
.A(n_2773),
.B(n_2467),
.Y(n_2812)
);

OAI21xp5_ASAP7_75t_SL g2813 ( 
.A1(n_2797),
.A2(n_2776),
.B(n_2775),
.Y(n_2813)
);

AOI21xp5_ASAP7_75t_L g2814 ( 
.A1(n_2788),
.A2(n_2786),
.B(n_2764),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2800),
.Y(n_2815)
);

NOR2xp33_ASAP7_75t_L g2816 ( 
.A(n_2807),
.B(n_2467),
.Y(n_2816)
);

OAI21xp5_ASAP7_75t_SL g2817 ( 
.A1(n_2806),
.A2(n_2481),
.B(n_2471),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2790),
.Y(n_2818)
);

OAI21xp5_ASAP7_75t_SL g2819 ( 
.A1(n_2799),
.A2(n_2481),
.B(n_2471),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2810),
.Y(n_2820)
);

AOI21xp5_ASAP7_75t_L g2821 ( 
.A1(n_2811),
.A2(n_2481),
.B(n_2784),
.Y(n_2821)
);

NOR2x1_ASAP7_75t_L g2822 ( 
.A(n_2803),
.B(n_2306),
.Y(n_2822)
);

INVxp67_ASAP7_75t_L g2823 ( 
.A(n_2805),
.Y(n_2823)
);

AOI221xp5_ASAP7_75t_L g2824 ( 
.A1(n_2796),
.A2(n_2404),
.B1(n_2394),
.B2(n_2357),
.C(n_2406),
.Y(n_2824)
);

BUFx2_ASAP7_75t_L g2825 ( 
.A(n_2812),
.Y(n_2825)
);

AOI221xp5_ASAP7_75t_L g2826 ( 
.A1(n_2792),
.A2(n_2404),
.B1(n_2357),
.B2(n_2408),
.C(n_2385),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2795),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2789),
.B(n_2382),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2804),
.Y(n_2829)
);

AOI221xp5_ASAP7_75t_L g2830 ( 
.A1(n_2801),
.A2(n_2385),
.B1(n_2435),
.B2(n_2422),
.C(n_2383),
.Y(n_2830)
);

BUFx2_ASAP7_75t_L g2831 ( 
.A(n_2794),
.Y(n_2831)
);

NAND2xp33_ASAP7_75t_R g2832 ( 
.A(n_2825),
.B(n_2791),
.Y(n_2832)
);

OAI221xp5_ASAP7_75t_L g2833 ( 
.A1(n_2820),
.A2(n_2798),
.B1(n_2801),
.B2(n_2809),
.C(n_2793),
.Y(n_2833)
);

O2A1O1Ixp5_ASAP7_75t_L g2834 ( 
.A1(n_2814),
.A2(n_2802),
.B(n_2809),
.C(n_2808),
.Y(n_2834)
);

AOI221xp5_ASAP7_75t_L g2835 ( 
.A1(n_2815),
.A2(n_2376),
.B1(n_2430),
.B2(n_2421),
.C(n_2285),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2823),
.B(n_2818),
.Y(n_2836)
);

AOI22xp5_ASAP7_75t_L g2837 ( 
.A1(n_2822),
.A2(n_2427),
.B1(n_2387),
.B2(n_2246),
.Y(n_2837)
);

AOI21xp5_ASAP7_75t_L g2838 ( 
.A1(n_2821),
.A2(n_2387),
.B(n_2316),
.Y(n_2838)
);

AOI222xp33_ASAP7_75t_L g2839 ( 
.A1(n_2826),
.A2(n_2316),
.B1(n_2378),
.B2(n_2252),
.C1(n_2308),
.C2(n_2303),
.Y(n_2839)
);

NOR3xp33_ASAP7_75t_L g2840 ( 
.A(n_2827),
.B(n_2291),
.C(n_2310),
.Y(n_2840)
);

NAND4xp75_ASAP7_75t_L g2841 ( 
.A(n_2829),
.B(n_72),
.C(n_70),
.D(n_71),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2831),
.Y(n_2842)
);

NOR4xp25_ASAP7_75t_L g2843 ( 
.A(n_2813),
.B(n_2310),
.C(n_2220),
.D(n_2222),
.Y(n_2843)
);

AOI222xp33_ASAP7_75t_L g2844 ( 
.A1(n_2824),
.A2(n_2303),
.B1(n_2302),
.B2(n_2222),
.C1(n_2220),
.C2(n_2211),
.Y(n_2844)
);

AOI22x1_ASAP7_75t_SL g2845 ( 
.A1(n_2842),
.A2(n_2832),
.B1(n_2834),
.B2(n_2833),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2836),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2841),
.Y(n_2847)
);

INVxp67_ASAP7_75t_L g2848 ( 
.A(n_2844),
.Y(n_2848)
);

O2A1O1Ixp33_ASAP7_75t_SL g2849 ( 
.A1(n_2838),
.A2(n_2816),
.B(n_2819),
.C(n_2828),
.Y(n_2849)
);

AO22x1_ASAP7_75t_L g2850 ( 
.A1(n_2840),
.A2(n_2817),
.B1(n_2835),
.B2(n_2843),
.Y(n_2850)
);

OAI22xp5_ASAP7_75t_L g2851 ( 
.A1(n_2837),
.A2(n_2830),
.B1(n_2211),
.B2(n_2290),
.Y(n_2851)
);

AOI22xp5_ASAP7_75t_L g2852 ( 
.A1(n_2839),
.A2(n_2290),
.B1(n_2281),
.B2(n_2301),
.Y(n_2852)
);

AO22x1_ASAP7_75t_L g2853 ( 
.A1(n_2842),
.A2(n_77),
.B1(n_74),
.B2(n_76),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2836),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2836),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2836),
.Y(n_2856)
);

A2O1A1Ixp33_ASAP7_75t_SL g2857 ( 
.A1(n_2842),
.A2(n_81),
.B(n_78),
.C(n_80),
.Y(n_2857)
);

NOR2xp33_ASAP7_75t_SL g2858 ( 
.A(n_2846),
.B(n_2281),
.Y(n_2858)
);

OAI21xp33_ASAP7_75t_L g2859 ( 
.A1(n_2854),
.A2(n_2281),
.B(n_2275),
.Y(n_2859)
);

OAI21x1_ASAP7_75t_L g2860 ( 
.A1(n_2847),
.A2(n_2856),
.B(n_2855),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2845),
.Y(n_2861)
);

AOI22xp5_ASAP7_75t_L g2862 ( 
.A1(n_2848),
.A2(n_2281),
.B1(n_2301),
.B2(n_671),
.Y(n_2862)
);

OA22x2_ASAP7_75t_L g2863 ( 
.A1(n_2851),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_2863)
);

AOI221xp5_ASAP7_75t_L g2864 ( 
.A1(n_2849),
.A2(n_2850),
.B1(n_2857),
.B2(n_2853),
.C(n_2852),
.Y(n_2864)
);

AOI22xp33_ASAP7_75t_L g2865 ( 
.A1(n_2848),
.A2(n_860),
.B1(n_893),
.B2(n_871),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2853),
.B(n_84),
.Y(n_2866)
);

OAI211xp5_ASAP7_75t_SL g2867 ( 
.A1(n_2846),
.A2(n_87),
.B(n_85),
.C(n_86),
.Y(n_2867)
);

OAI31xp33_ASAP7_75t_L g2868 ( 
.A1(n_2846),
.A2(n_89),
.A3(n_85),
.B(n_88),
.Y(n_2868)
);

NOR2xp33_ASAP7_75t_L g2869 ( 
.A(n_2845),
.B(n_88),
.Y(n_2869)
);

AOI221xp5_ASAP7_75t_L g2870 ( 
.A1(n_2848),
.A2(n_90),
.B1(n_91),
.B2(n_95),
.C(n_96),
.Y(n_2870)
);

OAI211xp5_ASAP7_75t_L g2871 ( 
.A1(n_2846),
.A2(n_97),
.B(n_90),
.C(n_96),
.Y(n_2871)
);

AOI22xp5_ASAP7_75t_L g2872 ( 
.A1(n_2846),
.A2(n_1303),
.B1(n_860),
.B2(n_893),
.Y(n_2872)
);

AOI221xp5_ASAP7_75t_L g2873 ( 
.A1(n_2848),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.C(n_101),
.Y(n_2873)
);

NOR2x1_ASAP7_75t_L g2874 ( 
.A(n_2846),
.B(n_99),
.Y(n_2874)
);

OAI21x1_ASAP7_75t_SL g2875 ( 
.A1(n_2866),
.A2(n_101),
.B(n_102),
.Y(n_2875)
);

OAI211xp5_ASAP7_75t_SL g2876 ( 
.A1(n_2861),
.A2(n_104),
.B(n_102),
.C(n_103),
.Y(n_2876)
);

OAI21xp5_ASAP7_75t_L g2877 ( 
.A1(n_2869),
.A2(n_871),
.B(n_860),
.Y(n_2877)
);

AOI21xp5_ASAP7_75t_SL g2878 ( 
.A1(n_2864),
.A2(n_104),
.B(n_107),
.Y(n_2878)
);

OAI211xp5_ASAP7_75t_SL g2879 ( 
.A1(n_2865),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_2879)
);

OAI311xp33_ASAP7_75t_L g2880 ( 
.A1(n_2862),
.A2(n_112),
.A3(n_113),
.B1(n_114),
.C1(n_115),
.Y(n_2880)
);

NAND3xp33_ASAP7_75t_SL g2881 ( 
.A(n_2870),
.B(n_113),
.C(n_115),
.Y(n_2881)
);

CKINVDCx16_ASAP7_75t_R g2882 ( 
.A(n_2874),
.Y(n_2882)
);

BUFx2_ASAP7_75t_L g2883 ( 
.A(n_2860),
.Y(n_2883)
);

OAI22xp33_ASAP7_75t_L g2884 ( 
.A1(n_2863),
.A2(n_871),
.B1(n_893),
.B2(n_860),
.Y(n_2884)
);

AND2x4_ASAP7_75t_L g2885 ( 
.A(n_2872),
.B(n_116),
.Y(n_2885)
);

OAI22xp5_ASAP7_75t_L g2886 ( 
.A1(n_2873),
.A2(n_860),
.B1(n_893),
.B2(n_871),
.Y(n_2886)
);

AOI221xp5_ASAP7_75t_L g2887 ( 
.A1(n_2871),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.C(n_120),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2858),
.B(n_2868),
.Y(n_2888)
);

BUFx6f_ASAP7_75t_L g2889 ( 
.A(n_2867),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2882),
.B(n_2859),
.Y(n_2890)
);

NAND3xp33_ASAP7_75t_L g2891 ( 
.A(n_2883),
.B(n_893),
.C(n_871),
.Y(n_2891)
);

NOR3xp33_ASAP7_75t_L g2892 ( 
.A(n_2877),
.B(n_117),
.C(n_118),
.Y(n_2892)
);

AND3x2_ASAP7_75t_L g2893 ( 
.A(n_2878),
.B(n_2887),
.C(n_2888),
.Y(n_2893)
);

NOR2x1_ASAP7_75t_L g2894 ( 
.A(n_2876),
.B(n_121),
.Y(n_2894)
);

AOI21xp5_ASAP7_75t_L g2895 ( 
.A1(n_2884),
.A2(n_122),
.B(n_123),
.Y(n_2895)
);

AND2x2_ASAP7_75t_L g2896 ( 
.A(n_2889),
.B(n_123),
.Y(n_2896)
);

NOR2x1_ASAP7_75t_L g2897 ( 
.A(n_2881),
.B(n_124),
.Y(n_2897)
);

AOI222xp33_ASAP7_75t_L g2898 ( 
.A1(n_2889),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.C1(n_128),
.C2(n_129),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2875),
.B(n_126),
.Y(n_2899)
);

NOR2x1_ASAP7_75t_L g2900 ( 
.A(n_2879),
.B(n_2886),
.Y(n_2900)
);

NAND3x1_ASAP7_75t_L g2901 ( 
.A(n_2880),
.B(n_129),
.C(n_130),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2901),
.Y(n_2902)
);

HB1xp67_ASAP7_75t_L g2903 ( 
.A(n_2894),
.Y(n_2903)
);

AND2x4_ASAP7_75t_L g2904 ( 
.A(n_2896),
.B(n_2885),
.Y(n_2904)
);

NAND3xp33_ASAP7_75t_L g2905 ( 
.A(n_2899),
.B(n_839),
.C(n_1103),
.Y(n_2905)
);

NOR2x1_ASAP7_75t_L g2906 ( 
.A(n_2890),
.B(n_133),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2897),
.Y(n_2907)
);

NOR2xp33_ASAP7_75t_L g2908 ( 
.A(n_2893),
.B(n_133),
.Y(n_2908)
);

CKINVDCx5p33_ASAP7_75t_R g2909 ( 
.A(n_2895),
.Y(n_2909)
);

NAND2x1_ASAP7_75t_L g2910 ( 
.A(n_2900),
.B(n_134),
.Y(n_2910)
);

NAND4xp25_ASAP7_75t_SL g2911 ( 
.A(n_2898),
.B(n_134),
.C(n_135),
.D(n_136),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2892),
.B(n_135),
.Y(n_2912)
);

AND2x4_ASAP7_75t_L g2913 ( 
.A(n_2907),
.B(n_2891),
.Y(n_2913)
);

OAI22xp5_ASAP7_75t_L g2914 ( 
.A1(n_2902),
.A2(n_1173),
.B1(n_1176),
.B2(n_1226),
.Y(n_2914)
);

OAI22xp5_ASAP7_75t_L g2915 ( 
.A1(n_2908),
.A2(n_1173),
.B1(n_1176),
.B2(n_1226),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_2903),
.B(n_139),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_L g2917 ( 
.A(n_2906),
.B(n_2910),
.Y(n_2917)
);

AOI311xp33_ASAP7_75t_L g2918 ( 
.A1(n_2912),
.A2(n_139),
.A3(n_141),
.B(n_142),
.C(n_143),
.Y(n_2918)
);

NOR3xp33_ASAP7_75t_L g2919 ( 
.A(n_2904),
.B(n_144),
.C(n_145),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_L g2920 ( 
.A(n_2904),
.B(n_144),
.Y(n_2920)
);

NOR2xp67_ASAP7_75t_L g2921 ( 
.A(n_2911),
.B(n_145),
.Y(n_2921)
);

AOI221xp5_ASAP7_75t_SL g2922 ( 
.A1(n_2909),
.A2(n_146),
.B1(n_149),
.B2(n_150),
.C(n_151),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2905),
.B(n_146),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2910),
.Y(n_2924)
);

NAND3xp33_ASAP7_75t_SL g2925 ( 
.A(n_2902),
.B(n_150),
.C(n_152),
.Y(n_2925)
);

AOI22xp33_ASAP7_75t_L g2926 ( 
.A1(n_2902),
.A2(n_839),
.B1(n_1121),
.B2(n_1117),
.Y(n_2926)
);

NAND4xp25_ASAP7_75t_L g2927 ( 
.A(n_2908),
.B(n_153),
.C(n_154),
.D(n_157),
.Y(n_2927)
);

AND2x2_ASAP7_75t_SL g2928 ( 
.A(n_2924),
.B(n_2917),
.Y(n_2928)
);

NOR3xp33_ASAP7_75t_SL g2929 ( 
.A(n_2925),
.B(n_2927),
.C(n_2923),
.Y(n_2929)
);

OR5x1_ASAP7_75t_L g2930 ( 
.A(n_2921),
.B(n_158),
.C(n_159),
.D(n_160),
.E(n_166),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2920),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2916),
.Y(n_2932)
);

XNOR2xp5_ASAP7_75t_L g2933 ( 
.A(n_2919),
.B(n_2915),
.Y(n_2933)
);

XNOR2x1_ASAP7_75t_L g2934 ( 
.A(n_2913),
.B(n_158),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2914),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_2918),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2928),
.Y(n_2937)
);

AOI32xp33_ASAP7_75t_L g2938 ( 
.A1(n_2936),
.A2(n_2926),
.A3(n_2922),
.B1(n_168),
.B2(n_169),
.Y(n_2938)
);

OAI22xp5_ASAP7_75t_SL g2939 ( 
.A1(n_2930),
.A2(n_159),
.B1(n_167),
.B2(n_171),
.Y(n_2939)
);

AO22x2_ASAP7_75t_L g2940 ( 
.A1(n_2934),
.A2(n_167),
.B1(n_171),
.B2(n_172),
.Y(n_2940)
);

OAI22xp5_ASAP7_75t_L g2941 ( 
.A1(n_2931),
.A2(n_1264),
.B1(n_1226),
.B2(n_1176),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2932),
.Y(n_2942)
);

AOI22xp33_ASAP7_75t_L g2943 ( 
.A1(n_2935),
.A2(n_1114),
.B1(n_1117),
.B2(n_1121),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2929),
.Y(n_2944)
);

AOI22xp5_ASAP7_75t_L g2945 ( 
.A1(n_2933),
.A2(n_1303),
.B1(n_1240),
.B2(n_1243),
.Y(n_2945)
);

OAI22xp5_ASAP7_75t_L g2946 ( 
.A1(n_2928),
.A2(n_1264),
.B1(n_1226),
.B2(n_1176),
.Y(n_2946)
);

AOI22xp5_ASAP7_75t_L g2947 ( 
.A1(n_2928),
.A2(n_1293),
.B1(n_1240),
.B2(n_1243),
.Y(n_2947)
);

AO22x2_ASAP7_75t_L g2948 ( 
.A1(n_2934),
.A2(n_174),
.B1(n_175),
.B2(n_177),
.Y(n_2948)
);

INVxp67_ASAP7_75t_L g2949 ( 
.A(n_2928),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2928),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2928),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2928),
.Y(n_2952)
);

NAND4xp75_ASAP7_75t_L g2953 ( 
.A(n_2928),
.B(n_174),
.C(n_179),
.D(n_181),
.Y(n_2953)
);

NOR4xp25_ASAP7_75t_L g2954 ( 
.A(n_2932),
.B(n_182),
.C(n_183),
.D(n_1085),
.Y(n_2954)
);

AOI22xp5_ASAP7_75t_L g2955 ( 
.A1(n_2928),
.A2(n_1293),
.B1(n_1291),
.B2(n_1266),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2928),
.Y(n_2956)
);

OAI22xp5_ASAP7_75t_SL g2957 ( 
.A1(n_2930),
.A2(n_182),
.B1(n_183),
.B2(n_839),
.Y(n_2957)
);

OAI22xp5_ASAP7_75t_L g2958 ( 
.A1(n_2928),
.A2(n_1264),
.B1(n_1291),
.B2(n_1262),
.Y(n_2958)
);

AOI22xp5_ASAP7_75t_L g2959 ( 
.A1(n_2949),
.A2(n_1262),
.B1(n_1266),
.B2(n_1012),
.Y(n_2959)
);

AOI22xp33_ASAP7_75t_L g2960 ( 
.A1(n_2937),
.A2(n_1121),
.B1(n_1114),
.B2(n_1117),
.Y(n_2960)
);

HB1xp67_ASAP7_75t_L g2961 ( 
.A(n_2950),
.Y(n_2961)
);

INVx2_ASAP7_75t_L g2962 ( 
.A(n_2951),
.Y(n_2962)
);

AND2x2_ASAP7_75t_L g2963 ( 
.A(n_2952),
.B(n_186),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_L g2964 ( 
.A(n_2956),
.B(n_2942),
.Y(n_2964)
);

OAI31xp33_ASAP7_75t_SL g2965 ( 
.A1(n_2944),
.A2(n_422),
.A3(n_193),
.B(n_198),
.Y(n_2965)
);

INVx3_ASAP7_75t_SL g2966 ( 
.A(n_2948),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2940),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2940),
.Y(n_2968)
);

AOI22xp33_ASAP7_75t_L g2969 ( 
.A1(n_2939),
.A2(n_1114),
.B1(n_1117),
.B2(n_1121),
.Y(n_2969)
);

AOI22xp5_ASAP7_75t_L g2970 ( 
.A1(n_2953),
.A2(n_1012),
.B1(n_1046),
.B2(n_1080),
.Y(n_2970)
);

BUFx2_ASAP7_75t_L g2971 ( 
.A(n_2957),
.Y(n_2971)
);

OAI31xp33_ASAP7_75t_L g2972 ( 
.A1(n_2958),
.A2(n_1085),
.A3(n_1084),
.B(n_1080),
.Y(n_2972)
);

AOI22xp5_ASAP7_75t_L g2973 ( 
.A1(n_2941),
.A2(n_1012),
.B1(n_1046),
.B2(n_1078),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2938),
.B(n_190),
.Y(n_2974)
);

OAI22xp33_ASAP7_75t_L g2975 ( 
.A1(n_2945),
.A2(n_1264),
.B1(n_1282),
.B2(n_1278),
.Y(n_2975)
);

OAI22xp5_ASAP7_75t_L g2976 ( 
.A1(n_2943),
.A2(n_1012),
.B1(n_1282),
.B2(n_1278),
.Y(n_2976)
);

AOI211xp5_ASAP7_75t_L g2977 ( 
.A1(n_2954),
.A2(n_1121),
.B(n_1114),
.C(n_1117),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2947),
.Y(n_2978)
);

OAI22xp5_ASAP7_75t_L g2979 ( 
.A1(n_2955),
.A2(n_1310),
.B1(n_1282),
.B2(n_1278),
.Y(n_2979)
);

OAI31xp33_ASAP7_75t_SL g2980 ( 
.A1(n_2946),
.A2(n_199),
.A3(n_201),
.B(n_204),
.Y(n_2980)
);

AO22x2_ASAP7_75t_L g2981 ( 
.A1(n_2937),
.A2(n_1084),
.B1(n_1078),
.B2(n_1077),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2937),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2937),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2937),
.Y(n_2984)
);

OAI22x1_ASAP7_75t_L g2985 ( 
.A1(n_2966),
.A2(n_839),
.B1(n_209),
.B2(n_212),
.Y(n_2985)
);

AOI22xp5_ASAP7_75t_L g2986 ( 
.A1(n_2961),
.A2(n_1310),
.B1(n_1248),
.B2(n_1247),
.Y(n_2986)
);

OAI211xp5_ASAP7_75t_SL g2987 ( 
.A1(n_2964),
.A2(n_206),
.B(n_214),
.C(n_215),
.Y(n_2987)
);

AOI211xp5_ASAP7_75t_L g2988 ( 
.A1(n_2983),
.A2(n_2984),
.B(n_2982),
.C(n_2962),
.Y(n_2988)
);

XOR2xp5_ASAP7_75t_L g2989 ( 
.A(n_2967),
.B(n_217),
.Y(n_2989)
);

AOI22xp33_ASAP7_75t_L g2990 ( 
.A1(n_2971),
.A2(n_1114),
.B1(n_839),
.B2(n_1074),
.Y(n_2990)
);

AO22x2_ASAP7_75t_L g2991 ( 
.A1(n_2968),
.A2(n_1077),
.B1(n_1060),
.B2(n_1056),
.Y(n_2991)
);

INVx2_ASAP7_75t_L g2992 ( 
.A(n_2963),
.Y(n_2992)
);

OAI22xp5_ASAP7_75t_L g2993 ( 
.A1(n_2969),
.A2(n_1310),
.B1(n_1248),
.B2(n_1247),
.Y(n_2993)
);

OAI22x1_ASAP7_75t_L g2994 ( 
.A1(n_2974),
.A2(n_2978),
.B1(n_2970),
.B2(n_2965),
.Y(n_2994)
);

XOR2xp5_ASAP7_75t_L g2995 ( 
.A(n_2979),
.B(n_219),
.Y(n_2995)
);

AOI22xp5_ASAP7_75t_L g2996 ( 
.A1(n_2975),
.A2(n_1248),
.B1(n_1247),
.B2(n_1235),
.Y(n_2996)
);

OAI22xp5_ASAP7_75t_SL g2997 ( 
.A1(n_2977),
.A2(n_839),
.B1(n_1060),
.B2(n_1056),
.Y(n_2997)
);

AOI211xp5_ASAP7_75t_L g2998 ( 
.A1(n_2980),
.A2(n_1074),
.B(n_1054),
.C(n_1033),
.Y(n_2998)
);

AOI322xp5_ASAP7_75t_L g2999 ( 
.A1(n_2960),
.A2(n_1054),
.A3(n_1043),
.B1(n_1033),
.B2(n_1235),
.C1(n_1189),
.C2(n_230),
.Y(n_2999)
);

OAI22xp5_ASAP7_75t_L g3000 ( 
.A1(n_2973),
.A2(n_1235),
.B1(n_1189),
.B2(n_1074),
.Y(n_3000)
);

AOI21xp33_ASAP7_75t_L g3001 ( 
.A1(n_2972),
.A2(n_220),
.B(n_221),
.Y(n_3001)
);

XNOR2xp5_ASAP7_75t_L g3002 ( 
.A(n_2981),
.B(n_225),
.Y(n_3002)
);

AOI22xp5_ASAP7_75t_L g3003 ( 
.A1(n_2976),
.A2(n_1189),
.B1(n_1043),
.B2(n_1074),
.Y(n_3003)
);

AOI22xp33_ASAP7_75t_L g3004 ( 
.A1(n_2981),
.A2(n_1074),
.B1(n_1052),
.B2(n_1019),
.Y(n_3004)
);

NAND4xp25_ASAP7_75t_SL g3005 ( 
.A(n_2959),
.B(n_226),
.C(n_228),
.D(n_231),
.Y(n_3005)
);

AOI22xp33_ASAP7_75t_L g3006 ( 
.A1(n_2961),
.A2(n_1052),
.B1(n_1019),
.B2(n_1021),
.Y(n_3006)
);

AOI21xp33_ASAP7_75t_L g3007 ( 
.A1(n_2961),
.A2(n_237),
.B(n_243),
.Y(n_3007)
);

OAI22xp33_ASAP7_75t_L g3008 ( 
.A1(n_2961),
.A2(n_1021),
.B1(n_1052),
.B2(n_1048),
.Y(n_3008)
);

NAND4xp25_ASAP7_75t_SL g3009 ( 
.A(n_2964),
.B(n_248),
.C(n_249),
.D(n_251),
.Y(n_3009)
);

AOI31xp33_ASAP7_75t_L g3010 ( 
.A1(n_2988),
.A2(n_252),
.A3(n_253),
.B(n_254),
.Y(n_3010)
);

AOI22xp33_ASAP7_75t_L g3011 ( 
.A1(n_2992),
.A2(n_1052),
.B1(n_1021),
.B2(n_1048),
.Y(n_3011)
);

AOI22xp33_ASAP7_75t_L g3012 ( 
.A1(n_3005),
.A2(n_1052),
.B1(n_1021),
.B2(n_1047),
.Y(n_3012)
);

AOI22xp33_ASAP7_75t_L g3013 ( 
.A1(n_2987),
.A2(n_1021),
.B1(n_1047),
.B2(n_1039),
.Y(n_3013)
);

AOI31xp33_ASAP7_75t_L g3014 ( 
.A1(n_2989),
.A2(n_257),
.A3(n_259),
.B(n_260),
.Y(n_3014)
);

AOI31xp33_ASAP7_75t_L g3015 ( 
.A1(n_3002),
.A2(n_261),
.A3(n_265),
.B(n_266),
.Y(n_3015)
);

AOI22xp33_ASAP7_75t_L g3016 ( 
.A1(n_2994),
.A2(n_1050),
.B1(n_1039),
.B2(n_1038),
.Y(n_3016)
);

AOI22xp33_ASAP7_75t_L g3017 ( 
.A1(n_2985),
.A2(n_1050),
.B1(n_1038),
.B2(n_1035),
.Y(n_3017)
);

AOI31xp33_ASAP7_75t_L g3018 ( 
.A1(n_2998),
.A2(n_269),
.A3(n_270),
.B(n_272),
.Y(n_3018)
);

AOI31xp33_ASAP7_75t_L g3019 ( 
.A1(n_3001),
.A2(n_273),
.A3(n_274),
.B(n_277),
.Y(n_3019)
);

AOI22xp33_ASAP7_75t_L g3020 ( 
.A1(n_2995),
.A2(n_1035),
.B1(n_1032),
.B2(n_1026),
.Y(n_3020)
);

AOI31xp33_ASAP7_75t_L g3021 ( 
.A1(n_3007),
.A2(n_279),
.A3(n_282),
.B(n_285),
.Y(n_3021)
);

AOI31xp33_ASAP7_75t_L g3022 ( 
.A1(n_2990),
.A2(n_286),
.A3(n_293),
.B(n_298),
.Y(n_3022)
);

HB1xp67_ASAP7_75t_L g3023 ( 
.A(n_3020),
.Y(n_3023)
);

OAI22xp5_ASAP7_75t_L g3024 ( 
.A1(n_3012),
.A2(n_2986),
.B1(n_2996),
.B2(n_3003),
.Y(n_3024)
);

INVx2_ASAP7_75t_L g3025 ( 
.A(n_3015),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_3019),
.Y(n_3026)
);

AOI22x1_ASAP7_75t_L g3027 ( 
.A1(n_3016),
.A2(n_2991),
.B1(n_2997),
.B2(n_2999),
.Y(n_3027)
);

HB1xp67_ASAP7_75t_L g3028 ( 
.A(n_3017),
.Y(n_3028)
);

OAI22xp5_ASAP7_75t_SL g3029 ( 
.A1(n_3013),
.A2(n_3006),
.B1(n_3004),
.B2(n_2993),
.Y(n_3029)
);

AOI22xp5_ASAP7_75t_L g3030 ( 
.A1(n_3011),
.A2(n_3009),
.B1(n_3000),
.B2(n_2991),
.Y(n_3030)
);

XNOR2x1_ASAP7_75t_L g3031 ( 
.A(n_3025),
.B(n_3014),
.Y(n_3031)
);

OAI21xp5_ASAP7_75t_L g3032 ( 
.A1(n_3026),
.A2(n_3021),
.B(n_3018),
.Y(n_3032)
);

AOI22xp33_ASAP7_75t_L g3033 ( 
.A1(n_3028),
.A2(n_3008),
.B1(n_3022),
.B2(n_3010),
.Y(n_3033)
);

AOI21xp5_ASAP7_75t_L g3034 ( 
.A1(n_3023),
.A2(n_3029),
.B(n_3024),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_3027),
.Y(n_3035)
);

OAI21xp5_ASAP7_75t_SL g3036 ( 
.A1(n_3030),
.A2(n_299),
.B(n_302),
.Y(n_3036)
);

OR2x6_ASAP7_75t_L g3037 ( 
.A(n_3025),
.B(n_1032),
.Y(n_3037)
);

AOI21xp33_ASAP7_75t_L g3038 ( 
.A1(n_3035),
.A2(n_307),
.B(n_309),
.Y(n_3038)
);

INVxp67_ASAP7_75t_L g3039 ( 
.A(n_3034),
.Y(n_3039)
);

OAI21x1_ASAP7_75t_L g3040 ( 
.A1(n_3032),
.A2(n_1026),
.B(n_1007),
.Y(n_3040)
);

NAND3xp33_ASAP7_75t_L g3041 ( 
.A(n_3031),
.B(n_1007),
.C(n_1000),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_3039),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_3040),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_3041),
.Y(n_3044)
);

OAI21x1_ASAP7_75t_L g3045 ( 
.A1(n_3042),
.A2(n_3033),
.B(n_3036),
.Y(n_3045)
);

AOI221xp5_ASAP7_75t_L g3046 ( 
.A1(n_3045),
.A2(n_3043),
.B1(n_3044),
.B2(n_3038),
.C(n_3037),
.Y(n_3046)
);

AOI211xp5_ASAP7_75t_L g3047 ( 
.A1(n_3046),
.A2(n_3037),
.B(n_319),
.C(n_320),
.Y(n_3047)
);


endmodule