module real_jpeg_5661_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_288;
wire n_78;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B1(n_23),
.B2(n_25),
.Y(n_19)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_1),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_1),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_1),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_1),
.Y(n_284)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_1),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_1),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_2),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_2),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_2),
.A2(n_55),
.B1(n_205),
.B2(n_275),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_2),
.A2(n_205),
.B1(n_286),
.B2(n_391),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g451 ( 
.A1(n_2),
.A2(n_205),
.B1(n_452),
.B2(n_454),
.Y(n_451)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_3),
.Y(n_191)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_3),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_3),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_4),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_4),
.A2(n_50),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_4),
.A2(n_50),
.B1(n_135),
.B2(n_137),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_4),
.A2(n_50),
.B1(n_286),
.B2(n_288),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_5),
.A2(n_43),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_5),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_5),
.A2(n_190),
.B1(n_259),
.B2(n_261),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g402 ( 
.A1(n_5),
.A2(n_190),
.B1(n_403),
.B2(n_404),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_5),
.A2(n_190),
.B1(n_425),
.B2(n_428),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_8),
.Y(n_119)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_8),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_8),
.Y(n_385)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_9),
.Y(n_95)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_10),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_10),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_10),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_11),
.A2(n_218),
.B1(n_220),
.B2(n_223),
.Y(n_217)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_11),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_11),
.A2(n_223),
.B1(n_261),
.B2(n_272),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_11),
.A2(n_182),
.B1(n_223),
.B2(n_306),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_L g365 ( 
.A1(n_11),
.A2(n_223),
.B1(n_366),
.B2(n_367),
.Y(n_365)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_12),
.Y(n_84)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_13),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_13),
.A2(n_163),
.B1(n_220),
.B2(n_379),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_13),
.B(n_385),
.C(n_386),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_13),
.B(n_91),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_13),
.B(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_13),
.B(n_133),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_13),
.B(n_213),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_14),
.A2(n_59),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_14),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_14),
.A2(n_76),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_14),
.A2(n_76),
.B1(n_219),
.B2(n_227),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_14),
.A2(n_76),
.B1(n_349),
.B2(n_350),
.Y(n_348)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_16),
.A2(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_16),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_16),
.A2(n_73),
.B1(n_170),
.B2(n_175),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_16),
.A2(n_73),
.B1(n_226),
.B2(n_231),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_16),
.A2(n_73),
.B1(n_210),
.B2(n_323),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_17),
.A2(n_54),
.B1(n_58),
.B2(n_61),
.Y(n_53)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_17),
.A2(n_61),
.B1(n_101),
.B2(n_103),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_17),
.A2(n_61),
.B1(n_170),
.B2(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_17),
.A2(n_61),
.B1(n_331),
.B2(n_332),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_18),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_18),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_18),
.A2(n_194),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_18),
.A2(n_194),
.B1(n_246),
.B2(n_248),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g397 ( 
.A1(n_18),
.A2(n_194),
.B1(n_307),
.B2(n_398),
.Y(n_397)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_63),
.B(n_529),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_51),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_27),
.B(n_51),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_38),
.B(n_45),
.Y(n_27)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_28),
.B(n_193),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_28),
.B(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_29),
.A2(n_52),
.B1(n_189),
.B2(n_274),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_29),
.B(n_163),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_34),
.Y(n_153)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_34),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_36),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_36),
.Y(n_207)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_36),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_36),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_38),
.B(n_193),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_38),
.A2(n_251),
.B(n_255),
.Y(n_250)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_42),
.Y(n_157)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_43),
.Y(n_195)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_44),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_44),
.B(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_52),
.B1(n_53),
.B2(n_62),
.Y(n_51)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_51),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_51),
.B(n_65),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_62),
.B1(n_69),
.B2(n_74),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_52),
.A2(n_53),
.B1(n_62),
.B2(n_74),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_52),
.A2(n_256),
.B(n_274),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_52),
.A2(n_62),
.B1(n_69),
.B2(n_501),
.Y(n_500)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_57),
.Y(n_254)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_62),
.A2(n_189),
.B(n_192),
.Y(n_188)
);

AO21x1_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_142),
.B(n_528),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_138),
.C(n_139),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_66),
.A2(n_67),
.B1(n_524),
.B2(n_525),
.Y(n_523)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_77),
.C(n_109),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_68),
.B(n_516),
.Y(n_515)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_77),
.A2(n_109),
.B1(n_110),
.B2(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_77),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_100),
.B1(n_105),
.B2(n_106),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g140 ( 
.A(n_78),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_78),
.A2(n_105),
.B1(n_202),
.B2(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_78),
.A2(n_105),
.B1(n_271),
.B2(n_322),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_78),
.A2(n_100),
.B1(n_105),
.B2(n_505),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_91),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_83),
.Y(n_465)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_85),
.Y(n_213)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_86),
.Y(n_353)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_89),
.Y(n_349)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_90),
.Y(n_204)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_90),
.Y(n_260)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_91),
.A2(n_140),
.B(n_141),
.Y(n_139)
);

AOI22x1_ASAP7_75t_L g268 ( 
.A1(n_91),
.A2(n_140),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_91),
.A2(n_140),
.B1(n_347),
.B2(n_348),
.Y(n_346)
);

AO22x2_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_94),
.B1(n_96),
.B2(n_98),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_94),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_95),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_95),
.Y(n_247)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_95),
.Y(n_405)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_95),
.Y(n_468)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_114),
.B1(n_117),
.B2(n_120),
.Y(n_113)
);

INVx11_ASAP7_75t_L g403 ( 
.A(n_96),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_97),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_97),
.Y(n_234)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_98),
.Y(n_469)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_101),
.Y(n_261)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_105),
.B(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_105),
.A2(n_258),
.B(n_303),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_109),
.A2(n_110),
.B1(n_503),
.B2(n_504),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_109),
.B(n_500),
.C(n_503),
.Y(n_511)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_132),
.B(n_134),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_111),
.A2(n_132),
.B1(n_217),
.B2(n_224),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_111),
.A2(n_378),
.B(n_380),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_111),
.A2(n_132),
.B1(n_402),
.B2(n_451),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_111),
.A2(n_380),
.B(n_451),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_112),
.B(n_245),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_112),
.A2(n_133),
.B1(n_225),
.B2(n_280),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_112),
.A2(n_133),
.B1(n_280),
.B2(n_330),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_112),
.A2(n_133),
.B1(n_330),
.B2(n_356),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_123),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_123),
.A2(n_244),
.B(n_402),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_129),
.B2(n_131),
.Y(n_123)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_127),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_128),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_130),
.Y(n_287)
);

BUFx5_ASAP7_75t_L g429 ( 
.A(n_130),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_132),
.A2(n_217),
.B(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_133),
.B(n_245),
.Y(n_380)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_134),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_136),
.Y(n_333)
);

INVx5_ASAP7_75t_L g453 ( 
.A(n_136),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_138),
.B(n_139),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_140),
.A2(n_201),
.B(n_208),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_140),
.B(n_269),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_140),
.A2(n_208),
.B(n_457),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_522),
.B(n_527),
.Y(n_142)
);

AOI21x1_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_494),
.B(n_519),
.Y(n_143)
);

OAI311xp33_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_315),
.A3(n_371),
.B1(n_488),
.C1(n_493),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_293),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_147),
.A2(n_490),
.B(n_491),
.Y(n_489)
);

NOR2x1_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_262),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_148),
.B(n_262),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_214),
.C(n_242),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_149),
.B(n_313),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_186),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_150),
.B(n_187),
.C(n_200),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_164),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_151),
.A2(n_164),
.B1(n_165),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_151),
.Y(n_300)
);

OAI32xp33_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_154),
.A3(n_155),
.B1(n_158),
.B2(n_162),
.Y(n_151)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_156),
.B(n_159),
.Y(n_158)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_SL g251 ( 
.A1(n_162),
.A2(n_163),
.B(n_252),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_163),
.A2(n_166),
.B(n_394),
.Y(n_421)
);

OAI21xp33_ASAP7_75t_SL g457 ( 
.A1(n_163),
.A2(n_323),
.B(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_173),
.B1(n_176),
.B2(n_179),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_166),
.A2(n_237),
.B1(n_282),
.B2(n_285),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_166),
.A2(n_285),
.B(n_335),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_166),
.A2(n_390),
.B(n_394),
.Y(n_389)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_167),
.A2(n_180),
.B1(n_236),
.B2(n_240),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_167),
.A2(n_174),
.B1(n_305),
.B2(n_310),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_167),
.B(n_397),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_167),
.A2(n_438),
.B1(n_439),
.B2(n_440),
.Y(n_437)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_169),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_169),
.Y(n_420)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_169),
.Y(n_432)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_171),
.Y(n_175)
);

BUFx8_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g290 ( 
.A(n_172),
.Y(n_290)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_172),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_172),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_185),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_199),
.B2(n_200),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_191),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_192),
.B(n_364),
.Y(n_363)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_209),
.Y(n_269)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_214),
.A2(n_215),
.B1(n_242),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_235),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_216),
.B(n_235),
.Y(n_266)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx4_ASAP7_75t_SL g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_230),
.Y(n_383)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_234),
.Y(n_379)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx4_ASAP7_75t_L g398 ( 
.A(n_238),
.Y(n_398)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_239),
.Y(n_387)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_242),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_249),
.C(n_257),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_243),
.B(n_257),
.Y(n_296)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

AOI32xp33_ASAP7_75t_L g463 ( 
.A1(n_247),
.A2(n_261),
.A3(n_459),
.B1(n_464),
.B2(n_466),
.Y(n_463)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_248),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_249),
.A2(n_250),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_263),
.B(n_278),
.C(n_291),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_278),
.B1(n_291),
.B2(n_292),
.Y(n_264)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_265),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_266),
.B(n_268),
.C(n_277),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_273),
.B1(n_276),
.B2(n_277),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_268),
.Y(n_276)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_273),
.Y(n_277)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_278),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_281),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_279),
.B(n_281),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_312),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_294),
.B(n_312),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_298),
.C(n_301),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_295),
.B(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_296),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_298),
.A2(n_299),
.B1(n_301),
.B2(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_301),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.C(n_311),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g478 ( 
.A(n_302),
.B(n_479),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_304),
.B(n_311),
.Y(n_479)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_305),
.Y(n_462)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx4_ASAP7_75t_SL g307 ( 
.A(n_308),
.Y(n_307)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp33_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_368),
.Y(n_315)
);

A2O1A1Ixp33_ASAP7_75t_SL g488 ( 
.A1(n_316),
.A2(n_368),
.B(n_489),
.C(n_492),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_340),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_317),
.B(n_340),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_327),
.C(n_339),
.Y(n_317)
);

FAx1_ASAP7_75t_SL g370 ( 
.A(n_318),
.B(n_327),
.CI(n_339),
.CON(n_370),
.SN(n_370)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_321),
.C(n_326),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_326),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_322),
.Y(n_347)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_328),
.A2(n_329),
.B1(n_334),
.B2(n_338),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_329),
.B(n_334),
.Y(n_360)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_334),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_334),
.A2(n_338),
.B1(n_362),
.B2(n_363),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_334),
.A2(n_360),
.B(n_363),
.Y(n_497)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_341),
.B(n_344),
.C(n_358),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_344),
.B1(n_358),
.B2(n_359),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_354),
.B(n_357),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_346),
.B(n_355),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_348),
.Y(n_505)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

FAx1_ASAP7_75t_SL g496 ( 
.A(n_357),
.B(n_497),
.CI(n_498),
.CON(n_496),
.SN(n_496)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_357),
.B(n_497),
.C(n_498),
.Y(n_518)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_365),
.Y(n_501)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_366),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_369),
.B(n_370),
.Y(n_492)
);

BUFx24_ASAP7_75t_SL g532 ( 
.A(n_370),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_372),
.A2(n_482),
.B(n_487),
.Y(n_371)
);

AO21x1_ASAP7_75t_SL g372 ( 
.A1(n_373),
.A2(n_471),
.B(n_481),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_374),
.A2(n_445),
.B(n_470),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_375),
.A2(n_408),
.B(n_444),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_388),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_376),
.B(n_388),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_381),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_377),
.A2(n_381),
.B1(n_382),
.B2(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_377),
.Y(n_442)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_399),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_389),
.B(n_400),
.C(n_407),
.Y(n_446)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_390),
.Y(n_439)
);

INVx6_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_397),
.Y(n_394)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_400),
.A2(n_401),
.B1(n_406),
.B2(n_407),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_403),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_409),
.A2(n_436),
.B(n_443),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_410),
.A2(n_422),
.B(n_435),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_421),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_418),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_419),
.Y(n_440)
);

INVx8_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_423),
.B(n_434),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_423),
.B(n_434),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_424),
.A2(n_430),
.B(n_433),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_424),
.Y(n_438)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx5_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx5_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_432),
.A2(n_433),
.B(n_462),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_441),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_437),
.B(n_441),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_446),
.B(n_447),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_460),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_449),
.A2(n_450),
.B1(n_455),
.B2(n_456),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_450),
.B(n_455),
.C(n_460),
.Y(n_472)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVxp33_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_463),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_461),
.B(n_463),
.Y(n_477)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

NAND2xp33_ASAP7_75t_SL g466 ( 
.A(n_467),
.B(n_469),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_472),
.B(n_473),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_474),
.A2(n_475),
.B1(n_478),
.B2(n_480),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_476),
.B(n_477),
.C(n_480),
.Y(n_483)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_478),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_484),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_483),
.B(n_484),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_508),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_496),
.B(n_507),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_496),
.B(n_507),
.Y(n_520)
);

BUFx24_ASAP7_75t_SL g531 ( 
.A(n_496),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_499),
.A2(n_500),
.B1(n_502),
.B2(n_506),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_499),
.A2(n_500),
.B1(n_514),
.B2(n_515),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_499),
.B(n_510),
.C(n_514),
.Y(n_526)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_502),
.Y(n_506)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_508),
.A2(n_520),
.B(n_521),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_509),
.B(n_518),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_509),
.B(n_518),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_510),
.A2(n_511),
.B1(n_512),
.B2(n_513),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_526),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_523),
.B(n_526),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_525),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_530),
.Y(n_529)
);


endmodule