module real_jpeg_21555_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_110;
wire n_205;
wire n_61;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_228;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_259;
wire n_103;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_210;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

INVx13_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_1),
.A2(n_30),
.B1(n_36),
.B2(n_37),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_2),
.A2(n_65),
.B1(n_72),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_2),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_2),
.A2(n_52),
.B1(n_54),
.B2(n_96),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_2),
.A2(n_36),
.B1(n_37),
.B2(n_96),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_96),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_3),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_4),
.Y(n_144)
);

AOI21xp33_ASAP7_75t_L g145 ( 
.A1(n_4),
.A2(n_52),
.B(n_70),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_4),
.A2(n_65),
.B1(n_72),
.B2(n_144),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_4),
.B(n_75),
.Y(n_193)
);

A2O1A1O1Ixp25_ASAP7_75t_L g204 ( 
.A1(n_4),
.A2(n_36),
.B(n_40),
.C(n_205),
.D(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_4),
.B(n_36),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_4),
.B(n_60),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_4),
.A2(n_25),
.B(n_220),
.Y(n_237)
);

A2O1A1O1Ixp25_ASAP7_75t_L g250 ( 
.A1(n_4),
.A2(n_54),
.B(n_55),
.C(n_154),
.D(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_4),
.B(n_54),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_5),
.A2(n_65),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_5),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_5),
.A2(n_52),
.B1(n_54),
.B2(n_73),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_73),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_5),
.A2(n_36),
.B1(n_37),
.B2(n_73),
.Y(n_249)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_7),
.B(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_7),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_7),
.A2(n_26),
.B1(n_148),
.B2(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_7),
.B(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_8),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_35)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_8),
.A2(n_38),
.B1(n_52),
.B2(n_54),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_38),
.Y(n_148)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_10),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_53),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_10),
.A2(n_53),
.B1(n_65),
.B2(n_72),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_53),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_11),
.A2(n_65),
.B1(n_72),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_11),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_11),
.A2(n_52),
.B1(n_54),
.B2(n_77),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_11),
.A2(n_36),
.B1(n_37),
.B2(n_77),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_77),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_13),
.A2(n_36),
.B1(n_37),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_46),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_13),
.A2(n_46),
.B1(n_52),
.B2(n_54),
.Y(n_114)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_131),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_129),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_104),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_20),
.B(n_104),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.C(n_85),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_21),
.A2(n_22),
.B1(n_78),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_48),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_23),
.B(n_50),
.C(n_62),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_24),
.B(n_34),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_25),
.A2(n_32),
.B(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_25),
.A2(n_29),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_25),
.A2(n_31),
.B1(n_88),
.B2(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_25),
.A2(n_219),
.B(n_220),
.Y(n_218)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_26),
.A2(n_225),
.B1(n_227),
.B2(n_228),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_26),
.B(n_221),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_27),
.A2(n_28),
.B1(n_41),
.B2(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_27),
.B(n_41),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_27),
.B(n_239),
.Y(n_238)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_28),
.A2(n_42),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_31),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_31),
.B(n_144),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_39),
.B1(n_45),
.B2(n_47),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_35),
.A2(n_39),
.B1(n_47),
.B2(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_37),
.B1(n_56),
.B2(n_57),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_36),
.B(n_56),
.Y(n_257)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

O2A1O1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_41),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_37),
.A2(n_59),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_39),
.A2(n_45),
.B1(n_47),
.B2(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_39),
.A2(n_47),
.B1(n_217),
.B2(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_39),
.A2(n_249),
.B(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_40),
.A2(n_43),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_40),
.B(n_170),
.Y(n_169)
);

CKINVDCx9p33_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_47),
.A2(n_92),
.B(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_47),
.B(n_171),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_47),
.A2(n_169),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_47),
.B(n_144),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_62),
.B2(n_63),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_55),
.B1(n_60),
.B2(n_61),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_51),
.Y(n_99)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_SL g55 ( 
.A1(n_52),
.A2(n_56),
.B(n_59),
.C(n_60),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_56),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_54),
.B1(n_67),
.B2(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_55),
.A2(n_60),
.B1(n_61),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_55),
.Y(n_152)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_71),
.B(n_74),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_64),
.A2(n_69),
.B1(n_71),
.B2(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_64),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_67),
.B(n_68),
.C(n_69),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_67),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_65),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_65),
.A2(n_67),
.B(n_144),
.C(n_145),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_69),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g140 ( 
.A1(n_69),
.A2(n_95),
.B(n_124),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_74),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_78),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_82),
.B2(n_84),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_79),
.A2(n_80),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_82),
.Y(n_119)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_81),
.A2(n_226),
.B(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_81),
.A2(n_235),
.B(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_82),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_83),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_85),
.B(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_93),
.C(n_97),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_87),
.B(n_91),
.Y(n_165)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_93),
.A2(n_94),
.B1(n_97),
.B2(n_98),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B(n_101),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_100),
.B(n_103),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_100),
.A2(n_151),
.B1(n_152),
.B2(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_100),
.A2(n_101),
.B(n_177),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_127),
.B2(n_128),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_116),
.B2(n_117),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_113),
.B(n_115),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_113),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_126),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_125),
.A2(n_173),
.B(n_174),
.Y(n_172)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_158),
.B(n_283),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_155),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_133),
.B(n_155),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.C(n_137),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_136),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_137),
.A2(n_138),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.C(n_149),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_140),
.B1(n_149),
.B2(n_150),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_146),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B(n_153),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_197),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI21xp33_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_181),
.B(n_196),
.Y(n_160)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_161),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_178),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_178),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.C(n_166),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_166),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_172),
.C(n_175),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_167),
.A2(n_168),
.B1(n_175),
.B2(n_176),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_182),
.B(n_184),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.C(n_189),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_185),
.B(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_187),
.A2(n_189),
.B1(n_190),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_187),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.C(n_194),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_191),
.A2(n_192),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_193),
.B(n_194),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_195),
.Y(n_259)
);

NOR3xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_281),
.C(n_282),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_275),
.B(n_280),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_262),
.B(n_274),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_243),
.B(n_261),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_222),
.B(n_242),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_211),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_203),
.B(n_211),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_204),
.A2(n_207),
.B1(n_208),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_204),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_205),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_206),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_218),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_216),
.C(n_218),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_219),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_231),
.B(n_241),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_229),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_224),
.B(n_229),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_236),
.B(n_240),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_233),
.B(n_234),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_244),
.B(n_245),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_254),
.B2(n_260),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_250),
.B1(n_252),
.B2(n_253),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_248),
.Y(n_253)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_250),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_253),
.C(n_260),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_251),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_254),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_258),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_263),
.B(n_264),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_270),
.C(n_272),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_266),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_272),
.B2(n_273),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_269),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_270),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_276),
.B(n_277),
.Y(n_280)
);


endmodule