module fake_jpeg_1746_n_632 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_632);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_632;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_5),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_61),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_63),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_65),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_66),
.Y(n_187)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g127 ( 
.A(n_67),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_68),
.Y(n_167)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx10_ASAP7_75t_L g153 ( 
.A(n_70),
.Y(n_153)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_73),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_27),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_74),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_22),
.B(n_9),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_75),
.B(n_81),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g165 ( 
.A(n_76),
.Y(n_165)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_77),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_78),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_82),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_27),
.Y(n_83)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_85),
.Y(n_193)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_86),
.B(n_87),
.Y(n_143)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_89),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

INVx4_ASAP7_75t_SL g92 ( 
.A(n_25),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_92),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_93),
.Y(n_197)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_32),
.B(n_10),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_45),
.C(n_26),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_95),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_96),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_27),
.Y(n_98)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

BUFx8_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_100),
.Y(n_186)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_101),
.Y(n_157)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_30),
.Y(n_103)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_8),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_104),
.A2(n_107),
.B(n_108),
.C(n_115),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_105),
.Y(n_173)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_8),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_11),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_24),
.Y(n_110)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_56),
.B(n_11),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_111),
.B(n_26),
.Y(n_172)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_25),
.Y(n_113)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_113),
.Y(n_171)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_30),
.Y(n_114)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_114),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_35),
.B(n_7),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_24),
.Y(n_116)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_116),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_44),
.Y(n_117)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_117),
.Y(n_200)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_37),
.Y(n_118)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_118),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_44),
.Y(n_119)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_119),
.Y(n_204)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_25),
.Y(n_120)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_120),
.Y(n_194)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_25),
.Y(n_121)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_121),
.Y(n_198)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_122),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_50),
.Y(n_123)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_132),
.B(n_172),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_92),
.A2(n_37),
.B1(n_45),
.B2(n_51),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g214 ( 
.A1(n_135),
.A2(n_169),
.B1(n_174),
.B2(n_27),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_115),
.B(n_41),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_139),
.B(n_90),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_61),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_145),
.B(n_152),
.Y(n_208)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_149),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_62),
.Y(n_152)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_83),
.Y(n_155)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_155),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_64),
.A2(n_37),
.B1(n_51),
.B2(n_42),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_163),
.A2(n_168),
.B1(n_135),
.B2(n_169),
.Y(n_217)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_166),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_111),
.A2(n_19),
.B1(n_20),
.B2(n_52),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_100),
.A2(n_51),
.B1(n_52),
.B2(n_50),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_94),
.A2(n_123),
.B1(n_119),
.B2(n_117),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_170),
.A2(n_34),
.B1(n_55),
.B2(n_24),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_172),
.B(n_199),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_104),
.A2(n_50),
.B1(n_52),
.B2(n_42),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_107),
.B(n_58),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_178),
.Y(n_215)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_70),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_183),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_108),
.B(n_39),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_185),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_103),
.B(n_39),
.Y(n_185)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_70),
.Y(n_190)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_68),
.B(n_35),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_191),
.B(n_19),
.Y(n_253)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_121),
.Y(n_195)
);

INVxp67_ASAP7_75t_SL g212 ( 
.A(n_195),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_76),
.B(n_58),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_196),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_73),
.A2(n_41),
.B1(n_53),
.B2(n_48),
.Y(n_199)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_105),
.Y(n_202)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_205),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_143),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_206),
.B(n_226),
.Y(n_300)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_174),
.A2(n_97),
.B1(n_95),
.B2(n_93),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_207),
.A2(n_217),
.B1(n_221),
.B2(n_175),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_209),
.B(n_223),
.Y(n_287)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_210),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_211),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_214),
.A2(n_243),
.B1(n_271),
.B2(n_142),
.Y(n_295)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_151),
.Y(n_216)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_216),
.Y(n_280)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_218),
.Y(n_281)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_158),
.Y(n_220)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_220),
.Y(n_292)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_163),
.A2(n_85),
.B1(n_78),
.B2(n_21),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_222),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_125),
.B(n_48),
.Y(n_223)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_134),
.Y(n_225)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_225),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_143),
.Y(n_226)
);

OA22x2_ASAP7_75t_L g227 ( 
.A1(n_148),
.A2(n_177),
.B1(n_147),
.B2(n_141),
.Y(n_227)
);

OA22x2_ASAP7_75t_L g317 ( 
.A1(n_227),
.A2(n_165),
.B1(n_181),
.B2(n_13),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_126),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_228),
.Y(n_283)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_229),
.Y(n_308)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_198),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_230),
.Y(n_341)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_192),
.Y(n_231)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_231),
.Y(n_312)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_127),
.Y(n_233)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_233),
.Y(n_313)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_176),
.Y(n_234)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_234),
.Y(n_318)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_171),
.Y(n_235)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_235),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_236),
.B(n_251),
.Y(n_305)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_127),
.Y(n_237)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_237),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_161),
.A2(n_53),
.B1(n_21),
.B2(n_40),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_238),
.A2(n_245),
.B1(n_252),
.B2(n_264),
.Y(n_322)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_176),
.Y(n_239)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_239),
.Y(n_340)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_240),
.Y(n_334)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_128),
.Y(n_241)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_241),
.Y(n_338)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_144),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_242),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_146),
.A2(n_90),
.B1(n_80),
.B2(n_76),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_125),
.A2(n_20),
.B1(n_19),
.B2(n_40),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_156),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_246),
.B(n_249),
.Y(n_311)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_133),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_247),
.Y(n_288)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_137),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_248),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_156),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_196),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_250),
.B(n_253),
.Y(n_339)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_140),
.Y(n_251)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_126),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_254),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_178),
.A2(n_34),
.B1(n_55),
.B2(n_20),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_255),
.B(n_274),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_130),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_256),
.Y(n_298)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_150),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_263),
.Y(n_285)
);

INVx8_ASAP7_75t_L g258 ( 
.A(n_130),
.Y(n_258)
);

BUFx24_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_167),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_259),
.Y(n_310)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_164),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_260),
.B(n_262),
.Y(n_314)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_180),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_136),
.B(n_12),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_131),
.A2(n_80),
.B1(n_34),
.B2(n_12),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_189),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_265),
.B(n_270),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_167),
.B(n_12),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_268),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_153),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_160),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_273),
.Y(n_301)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_131),
.Y(n_270)
);

INVx8_ASAP7_75t_L g271 ( 
.A(n_175),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_124),
.B(n_34),
.C(n_12),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_124),
.C(n_187),
.Y(n_286)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_173),
.Y(n_273)
);

FAx1_ASAP7_75t_SL g274 ( 
.A(n_153),
.B(n_34),
.CI(n_7),
.CON(n_274),
.SN(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_160),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_275),
.B(n_278),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_138),
.B(n_7),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_173),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_279),
.B(n_2),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_286),
.B(n_304),
.Y(n_358)
);

OAI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_154),
.B1(n_203),
.B2(n_197),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_289),
.A2(n_290),
.B1(n_293),
.B2(n_325),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_252),
.A2(n_204),
.B1(n_200),
.B2(n_203),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_207),
.A2(n_214),
.B(n_266),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_294),
.A2(n_296),
.B(n_342),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_295),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_215),
.A2(n_162),
.B1(n_179),
.B2(n_129),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_213),
.B(n_204),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_299),
.B(n_303),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_227),
.B(n_200),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_236),
.B(n_165),
.C(n_153),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_227),
.B(n_165),
.C(n_193),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_307),
.B(n_317),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_221),
.A2(n_197),
.B1(n_193),
.B2(n_181),
.Y(n_309)
);

OAI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_309),
.A2(n_228),
.B1(n_259),
.B2(n_256),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_208),
.B(n_0),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_320),
.B(n_321),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_274),
.B(n_0),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_277),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_274),
.B(n_1),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_326),
.B(n_329),
.Y(n_367)
);

FAx1_ASAP7_75t_L g327 ( 
.A(n_255),
.B(n_1),
.CI(n_2),
.CON(n_327),
.SN(n_327)
);

AOI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_327),
.A2(n_304),
.B(n_317),
.Y(n_380)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_328),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_248),
.B(n_272),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_224),
.B(n_3),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_330),
.B(n_3),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_214),
.A2(n_14),
.B1(n_17),
.B2(n_16),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_331),
.A2(n_342),
.B1(n_211),
.B2(n_244),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_261),
.B(n_6),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_336),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_279),
.A2(n_6),
.B1(n_13),
.B2(n_15),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_339),
.B(n_230),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_343),
.B(n_359),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_335),
.Y(n_347)
);

INVx3_ASAP7_75t_SL g430 ( 
.A(n_347),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_314),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_348),
.B(n_352),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_294),
.A2(n_273),
.B1(n_270),
.B2(n_212),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_349),
.A2(n_362),
.B1(n_372),
.B2(n_374),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_293),
.A2(n_238),
.B1(n_243),
.B2(n_254),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_350),
.A2(n_360),
.B1(n_365),
.B2(n_370),
.Y(n_395)
);

AOI32xp33_ASAP7_75t_L g352 ( 
.A1(n_321),
.A2(n_276),
.A3(n_244),
.B1(n_205),
.B2(n_242),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_308),
.Y(n_354)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_354),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_307),
.A2(n_212),
.B1(n_234),
.B2(n_239),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_355),
.A2(n_380),
.B(n_324),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_L g419 ( 
.A1(n_356),
.A2(n_357),
.B1(n_283),
.B2(n_335),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_299),
.B(n_251),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_333),
.A2(n_271),
.B1(n_258),
.B2(n_276),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_287),
.B(n_219),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_361),
.B(n_364),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_303),
.A2(n_219),
.B1(n_232),
.B2(n_15),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_341),
.Y(n_363)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_363),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_323),
.B(n_291),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_333),
.A2(n_232),
.B1(n_4),
.B2(n_5),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g366 ( 
.A(n_326),
.B(n_327),
.Y(n_366)
);

CKINVDCx14_ASAP7_75t_R g413 ( 
.A(n_366),
.Y(n_413)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_308),
.Y(n_368)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_368),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_369),
.B(n_373),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_329),
.A2(n_331),
.B1(n_322),
.B2(n_286),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_290),
.A2(n_6),
.B1(n_18),
.B2(n_3),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_285),
.B(n_4),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_327),
.A2(n_4),
.B1(n_18),
.B2(n_305),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_300),
.B(n_305),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_375),
.B(n_389),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_337),
.B(n_320),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_376),
.B(n_377),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_330),
.B(n_305),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_325),
.A2(n_317),
.B1(n_306),
.B2(n_311),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_378),
.A2(n_384),
.B1(n_324),
.B2(n_302),
.Y(n_418)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_341),
.Y(n_379)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_379),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_313),
.B(n_316),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_381),
.B(n_387),
.Y(n_433)
);

INVx3_ASAP7_75t_SL g382 ( 
.A(n_283),
.Y(n_382)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_382),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_317),
.A2(n_306),
.B1(n_296),
.B2(n_298),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_383),
.A2(n_391),
.B1(n_315),
.B2(n_332),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_337),
.A2(n_310),
.B1(n_301),
.B2(n_316),
.Y(n_384)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_312),
.Y(n_386)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_386),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_312),
.B(n_313),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_302),
.Y(n_388)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_388),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_280),
.B(n_281),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g429 ( 
.A(n_390),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_280),
.A2(n_281),
.B1(n_297),
.B2(n_292),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_324),
.Y(n_392)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_392),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_391),
.Y(n_393)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_393),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_371),
.A2(n_340),
.B(n_318),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_394),
.A2(n_396),
.B(n_404),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_371),
.A2(n_340),
.B(n_318),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_358),
.B(n_367),
.C(n_370),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_397),
.B(n_398),
.C(n_402),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_358),
.B(n_292),
.Y(n_398)
);

FAx1_ASAP7_75t_SL g401 ( 
.A(n_367),
.B(n_297),
.CI(n_314),
.CON(n_401),
.SN(n_401)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_401),
.B(n_353),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_377),
.B(n_319),
.C(n_314),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_390),
.A2(n_385),
.B(n_380),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_410),
.A2(n_417),
.B(n_434),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_344),
.B(n_319),
.C(n_288),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_414),
.B(n_402),
.C(n_397),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_347),
.Y(n_415)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_415),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_366),
.A2(n_288),
.B(n_338),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_418),
.A2(n_425),
.B1(n_431),
.B2(n_382),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_419),
.A2(n_421),
.B1(n_422),
.B2(n_424),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_385),
.A2(n_315),
.B1(n_332),
.B2(n_334),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_385),
.A2(n_344),
.B1(n_346),
.B2(n_383),
.Y(n_424)
);

OAI22x1_ASAP7_75t_SL g425 ( 
.A1(n_346),
.A2(n_282),
.B1(n_334),
.B2(n_338),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_387),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_427),
.B(n_359),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_366),
.A2(n_282),
.B1(n_284),
.B2(n_378),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_381),
.Y(n_432)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_432),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_380),
.A2(n_284),
.B(n_348),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_347),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_435),
.B(n_382),
.Y(n_439)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_400),
.Y(n_437)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_437),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_439),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_440),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_433),
.B(n_369),
.Y(n_441)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_441),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_433),
.B(n_351),
.Y(n_442)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_442),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_427),
.B(n_432),
.Y(n_443)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_443),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_429),
.A2(n_375),
.B(n_349),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_444),
.A2(n_450),
.B(n_456),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_420),
.B(n_343),
.Y(n_445)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_445),
.A2(n_449),
.B(n_472),
.Y(n_502)
);

NAND4xp25_ASAP7_75t_SL g446 ( 
.A(n_421),
.B(n_384),
.C(n_374),
.D(n_373),
.Y(n_446)
);

INVx13_ASAP7_75t_L g500 ( 
.A(n_446),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_398),
.B(n_351),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_447),
.B(n_448),
.C(n_451),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_429),
.A2(n_360),
.B1(n_350),
.B2(n_365),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_426),
.B(n_353),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_424),
.A2(n_362),
.B1(n_372),
.B2(n_392),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_452),
.A2(n_470),
.B1(n_395),
.B2(n_425),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_404),
.B(n_413),
.C(n_426),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_454),
.B(n_455),
.C(n_458),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_413),
.B(n_414),
.C(n_434),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_431),
.A2(n_345),
.B1(n_357),
.B2(n_352),
.Y(n_456)
);

XNOR2x1_ASAP7_75t_L g457 ( 
.A(n_417),
.B(n_354),
.Y(n_457)
);

XOR2x2_ASAP7_75t_SL g486 ( 
.A(n_457),
.B(n_401),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_410),
.B(n_368),
.C(n_386),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_420),
.B(n_376),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_459),
.B(n_406),
.Y(n_501)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_400),
.Y(n_460)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_460),
.Y(n_497)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_408),
.Y(n_462)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_462),
.Y(n_498)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_408),
.Y(n_463)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_463),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_428),
.A2(n_389),
.B(n_363),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_464),
.A2(n_473),
.B(n_423),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_428),
.B(n_388),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_465),
.B(n_467),
.C(n_469),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_466),
.B(n_412),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_403),
.B(n_379),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_393),
.B(n_284),
.C(n_407),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_405),
.B(n_403),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_405),
.A2(n_401),
.B(n_416),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_436),
.A2(n_418),
.B1(n_407),
.B2(n_399),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_480),
.A2(n_485),
.B(n_493),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_484),
.A2(n_499),
.B1(n_480),
.B2(n_491),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_468),
.A2(n_394),
.B(n_396),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_486),
.B(n_437),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_456),
.A2(n_395),
.B1(n_422),
.B2(n_399),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_488),
.A2(n_491),
.B1(n_478),
.B2(n_483),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_438),
.B(n_416),
.C(n_411),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_489),
.B(n_490),
.C(n_504),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_438),
.B(n_411),
.C(n_423),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_491),
.A2(n_452),
.B1(n_453),
.B2(n_462),
.Y(n_519)
);

NOR2x1_ASAP7_75t_L g493 ( 
.A(n_454),
.B(n_440),
.Y(n_493)
);

INVxp67_ASAP7_75t_SL g512 ( 
.A(n_494),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_469),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_495),
.B(n_471),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_440),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_496),
.B(n_501),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_464),
.A2(n_412),
.B1(n_430),
.B2(n_406),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_442),
.B(n_409),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_503),
.B(n_463),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_448),
.B(n_409),
.C(n_415),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_447),
.B(n_435),
.C(n_430),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_505),
.B(n_506),
.C(n_482),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_455),
.B(n_430),
.C(n_458),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_476),
.Y(n_507)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_507),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_485),
.A2(n_468),
.B(n_461),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_508),
.A2(n_525),
.B(n_477),
.Y(n_554)
);

XOR2x2_ASAP7_75t_L g509 ( 
.A(n_481),
.B(n_465),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_509),
.B(n_510),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_SL g510 ( 
.A(n_481),
.B(n_451),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_SL g540 ( 
.A(n_510),
.B(n_522),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_493),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_511),
.B(n_524),
.Y(n_537)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_476),
.Y(n_513)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_513),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g514 ( 
.A(n_499),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_514),
.B(n_494),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_492),
.A2(n_443),
.B1(n_473),
.B2(n_466),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_515),
.A2(n_518),
.B1(n_520),
.B2(n_531),
.Y(n_550)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_474),
.Y(n_516)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_516),
.Y(n_548)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_474),
.Y(n_517)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_517),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_492),
.A2(n_461),
.B1(n_450),
.B2(n_444),
.Y(n_518)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_519),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_484),
.A2(n_441),
.B1(n_467),
.B2(n_457),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_487),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_478),
.A2(n_446),
.B(n_460),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_497),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_526),
.B(n_527),
.Y(n_539)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_497),
.Y(n_527)
);

CKINVDCx14_ASAP7_75t_R g557 ( 
.A(n_528),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_529),
.B(n_530),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_479),
.B(n_471),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_533),
.A2(n_488),
.B1(n_500),
.B2(n_475),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_534),
.B(n_506),
.C(n_504),
.Y(n_545)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_498),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_535),
.B(n_483),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_538),
.B(n_545),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_541),
.B(n_522),
.Y(n_562)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_543),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_534),
.B(n_490),
.C(n_479),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_546),
.B(n_551),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_547),
.A2(n_519),
.B1(n_531),
.B2(n_512),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_530),
.B(n_495),
.C(n_489),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_532),
.B(n_505),
.C(n_482),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_552),
.B(n_556),
.C(n_558),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_554),
.A2(n_524),
.B(n_520),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_523),
.B(n_475),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_555),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_532),
.B(n_477),
.C(n_486),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_509),
.B(n_487),
.C(n_502),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_511),
.B(n_498),
.C(n_500),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_559),
.B(n_507),
.C(n_513),
.Y(n_571)
);

NOR2xp67_ASAP7_75t_L g589 ( 
.A(n_562),
.B(n_579),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_550),
.A2(n_515),
.B1(n_525),
.B2(n_533),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_563),
.A2(n_578),
.B1(n_543),
.B2(n_542),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_536),
.B(n_521),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_564),
.B(n_567),
.Y(n_583)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_565),
.Y(n_588)
);

INVxp33_ASAP7_75t_SL g566 ( 
.A(n_555),
.Y(n_566)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_566),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_536),
.B(n_521),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_552),
.B(n_518),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_568),
.B(n_569),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_551),
.B(n_508),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_570),
.B(n_576),
.Y(n_592)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_571),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_545),
.B(n_529),
.C(n_517),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_573),
.B(n_577),
.Y(n_580)
);

FAx1_ASAP7_75t_SL g576 ( 
.A(n_556),
.B(n_516),
.CI(n_526),
.CON(n_576),
.SN(n_576)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_546),
.B(n_527),
.C(n_535),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_558),
.A2(n_537),
.B(n_554),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_557),
.B(n_553),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_569),
.B(n_537),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_581),
.B(n_563),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_575),
.B(n_559),
.C(n_540),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_582),
.B(n_585),
.Y(n_608)
);

NOR2xp67_ASAP7_75t_SL g584 ( 
.A(n_560),
.B(n_540),
.Y(n_584)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_584),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_577),
.B(n_553),
.C(n_547),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_561),
.B(n_539),
.Y(n_587)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_587),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_568),
.B(n_542),
.C(n_544),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_590),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_SL g601 ( 
.A1(n_591),
.A2(n_565),
.B1(n_576),
.B2(n_544),
.Y(n_601)
);

NOR2x1_ASAP7_75t_L g595 ( 
.A(n_574),
.B(n_539),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_595),
.A2(n_570),
.B(n_571),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_594),
.B(n_573),
.C(n_572),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_596),
.B(n_597),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_SL g597 ( 
.A(n_580),
.B(n_560),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_586),
.B(n_590),
.C(n_581),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_599),
.B(n_601),
.Y(n_611)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_600),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_603),
.B(n_605),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_586),
.B(n_564),
.C(n_567),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_585),
.B(n_562),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_SL g615 ( 
.A(n_606),
.B(n_607),
.Y(n_615)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_587),
.Y(n_607)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_599),
.B(n_582),
.Y(n_610)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_610),
.Y(n_620)
);

O2A1O1Ixp33_ASAP7_75t_SL g613 ( 
.A1(n_602),
.A2(n_592),
.B(n_593),
.C(n_595),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_L g621 ( 
.A1(n_613),
.A2(n_600),
.B(n_601),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_604),
.B(n_588),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_614),
.B(n_616),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_596),
.B(n_583),
.C(n_592),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_617),
.A2(n_598),
.B(n_589),
.Y(n_618)
);

OAI21xp5_ASAP7_75t_L g625 ( 
.A1(n_618),
.A2(n_613),
.B(n_611),
.Y(n_625)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_610),
.B(n_608),
.Y(n_619)
);

XOR2xp5_ASAP7_75t_L g626 ( 
.A(n_619),
.B(n_612),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_SL g624 ( 
.A1(n_621),
.A2(n_622),
.B(n_616),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_SL g622 ( 
.A(n_609),
.B(n_615),
.Y(n_622)
);

AOI21x1_ASAP7_75t_L g627 ( 
.A1(n_624),
.A2(n_625),
.B(n_623),
.Y(n_627)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_626),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_SL g629 ( 
.A1(n_627),
.A2(n_620),
.B1(n_576),
.B2(n_605),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_SL g630 ( 
.A1(n_629),
.A2(n_628),
.B(n_583),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_L g631 ( 
.A1(n_630),
.A2(n_548),
.B1(n_549),
.B2(n_627),
.Y(n_631)
);

XOR2xp5_ASAP7_75t_L g632 ( 
.A(n_631),
.B(n_548),
.Y(n_632)
);


endmodule