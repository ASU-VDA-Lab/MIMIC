module fake_jpeg_12497_n_134 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_134);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx10_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_59),
.Y(n_76)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_66),
.Y(n_70)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_SL g73 ( 
.A(n_65),
.B(n_67),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_50),
.B(n_1),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_53),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_75),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_64),
.B(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_80),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_43),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_57),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_78),
.A2(n_44),
.B(n_55),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_81),
.Y(n_100)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_83),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_70),
.B(n_42),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_44),
.B1(n_57),
.B2(n_59),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_94),
.B1(n_4),
.B2(n_6),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_90),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_49),
.B1(n_51),
.B2(n_55),
.Y(n_88)
);

AO21x2_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_4),
.B(n_7),
.Y(n_111)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_92),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_56),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_93),
.B(n_68),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_49),
.B1(n_46),
.B2(n_3),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_54),
.B1(n_2),
.B2(n_3),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_109),
.B1(n_10),
.B2(n_15),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_40),
.C(n_12),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_92),
.A2(n_68),
.B(n_54),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_107),
.B(n_96),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_85),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_103),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_88),
.A2(n_1),
.B(n_2),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_22),
.Y(n_110)
);

NAND2x1p5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_16),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_111),
.A2(n_7),
.B(n_8),
.Y(n_115)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_112),
.A2(n_113),
.B1(n_117),
.B2(n_121),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_101),
.A2(n_111),
.B1(n_88),
.B2(n_100),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_114),
.A2(n_115),
.B1(n_118),
.B2(n_119),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_108),
.Y(n_119)
);

AOI322xp5_ASAP7_75t_SL g125 ( 
.A1(n_120),
.A2(n_110),
.A3(n_20),
.B1(n_23),
.B2(n_24),
.C1(n_25),
.C2(n_26),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_17),
.C(n_18),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_119),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_116),
.Y(n_126)
);

NOR3xp33_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_102),
.C(n_27),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_127),
.C(n_128),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_116),
.C(n_105),
.Y(n_127)
);

NOR2x1_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_123),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_SL g131 ( 
.A1(n_130),
.A2(n_111),
.B(n_125),
.Y(n_131)
);

AOI21x1_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_19),
.B(n_31),
.Y(n_132)
);

NAND4xp25_ASAP7_75t_SL g133 ( 
.A(n_132),
.B(n_34),
.C(n_35),
.D(n_36),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_38),
.Y(n_134)
);


endmodule