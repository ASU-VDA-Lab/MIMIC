module real_aes_3773_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_319;
wire n_112;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_119;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_653;
wire n_290;
wire n_365;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_183;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_500;
wire n_307;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g402 ( .A(n_0), .Y(n_402) );
AOI22x1_ASAP7_75t_L g183 ( .A1(n_1), .A2(n_40), .B1(n_184), .B2(n_189), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_2), .B(n_259), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_3), .B(n_289), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_4), .A2(n_30), .B1(n_301), .B2(n_348), .Y(n_347) );
AOI211xp5_ASAP7_75t_L g98 ( .A1(n_5), .A2(n_99), .B(n_124), .C(n_161), .Y(n_98) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_6), .A2(n_10), .B1(n_126), .B2(n_131), .Y(n_125) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_7), .A2(n_32), .B1(n_319), .B2(n_359), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_8), .A2(n_51), .B1(n_364), .B2(n_379), .Y(n_386) );
INVx1_ASAP7_75t_L g397 ( .A(n_9), .Y(n_397) );
INVx1_ASAP7_75t_L g121 ( .A(n_11), .Y(n_121) );
INVxp67_ASAP7_75t_L g150 ( .A(n_11), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_11), .B(n_60), .Y(n_157) );
AOI221xp5_ASAP7_75t_L g192 ( .A1(n_12), .A2(n_20), .B1(n_193), .B2(n_197), .C(n_200), .Y(n_192) );
INVx1_ASAP7_75t_L g400 ( .A(n_13), .Y(n_400) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_14), .A2(n_57), .B(n_252), .Y(n_251) );
OA21x2_ASAP7_75t_L g340 ( .A1(n_14), .A2(n_57), .B(n_252), .Y(n_340) );
NAND2xp5_ASAP7_75t_SL g117 ( .A(n_15), .B(n_106), .Y(n_117) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_16), .A2(n_54), .B1(n_364), .B2(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g394 ( .A(n_17), .Y(n_394) );
HB1xp67_ASAP7_75t_L g90 ( .A(n_18), .Y(n_90) );
BUFx3_ASAP7_75t_L g212 ( .A(n_19), .Y(n_212) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_21), .Y(n_106) );
AO22x1_ASAP7_75t_L g280 ( .A1(n_22), .A2(n_65), .B1(n_281), .B2(n_285), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_23), .Y(n_304) );
AND2x2_ASAP7_75t_L g318 ( .A(n_24), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_25), .B(n_285), .Y(n_311) );
AO22x1_ASAP7_75t_L g161 ( .A1(n_26), .A2(n_71), .B1(n_162), .B2(n_169), .Y(n_161) );
HB1xp67_ASAP7_75t_L g89 ( .A(n_27), .Y(n_89) );
AOI22x1_ASAP7_75t_L g363 ( .A1(n_27), .A2(n_75), .B1(n_343), .B2(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g107 ( .A(n_28), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_28), .B(n_59), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_29), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_31), .B(n_256), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g140 ( .A1(n_33), .A2(n_64), .B1(n_141), .B2(n_151), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_34), .B(n_263), .Y(n_262) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_35), .Y(n_82) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_36), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g252 ( .A(n_37), .Y(n_252) );
AO22x1_ASAP7_75t_L g200 ( .A1(n_38), .A2(n_53), .B1(n_201), .B2(n_203), .Y(n_200) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_39), .Y(n_223) );
AND2x4_ASAP7_75t_L g227 ( .A(n_39), .B(n_221), .Y(n_227) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_41), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_42), .Y(n_94) );
INVx2_ASAP7_75t_L g381 ( .A(n_43), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_44), .A2(n_95), .B1(n_96), .B2(n_647), .Y(n_646) );
CKINVDCx5p33_ASAP7_75t_R g647 ( .A(n_44), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_45), .A2(n_61), .B1(n_301), .B2(n_343), .Y(n_342) );
CKINVDCx14_ASAP7_75t_R g292 ( .A(n_46), .Y(n_292) );
AND2x2_ASAP7_75t_L g326 ( .A(n_47), .B(n_285), .Y(n_326) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_47), .Y(n_641) );
HB1xp67_ASAP7_75t_L g84 ( .A(n_48), .Y(n_84) );
OA22x2_ASAP7_75t_L g111 ( .A1(n_49), .A2(n_60), .B1(n_106), .B2(n_110), .Y(n_111) );
INVx1_ASAP7_75t_L g137 ( .A(n_49), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_50), .B(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_52), .B(n_249), .Y(n_248) );
AOI221xp5_ASAP7_75t_L g172 ( .A1(n_55), .A2(n_62), .B1(n_173), .B2(n_177), .C(n_182), .Y(n_172) );
NAND2x1p5_ASAP7_75t_L g329 ( .A(n_56), .B(n_276), .Y(n_329) );
CKINVDCx14_ASAP7_75t_R g368 ( .A(n_58), .Y(n_368) );
INVx1_ASAP7_75t_L g123 ( .A(n_59), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_59), .B(n_135), .Y(n_160) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_59), .Y(n_215) );
OAI21xp33_ASAP7_75t_L g138 ( .A1(n_60), .A2(n_66), .B(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_63), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g109 ( .A(n_66), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_66), .B(n_74), .Y(n_158) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_67), .Y(n_236) );
BUFx5_ASAP7_75t_L g260 ( .A(n_67), .Y(n_260) );
INVx1_ASAP7_75t_L g284 ( .A(n_67), .Y(n_284) );
INVx2_ASAP7_75t_L g404 ( .A(n_68), .Y(n_404) );
NAND2xp33_ASAP7_75t_L g322 ( .A(n_69), .B(n_323), .Y(n_322) );
INVx2_ASAP7_75t_SL g221 ( .A(n_70), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_72), .B(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_73), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_74), .B(n_116), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_76), .B(n_274), .Y(n_313) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_207), .B1(n_224), .B2(n_237), .C(n_639), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_92), .Y(n_78) );
OAI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_81), .B1(n_86), .B2(n_87), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
AOI22xp5_ASAP7_75t_L g81 ( .A1(n_82), .A2(n_83), .B1(n_84), .B2(n_85), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_82), .Y(n_85) );
CKINVDCx14_ASAP7_75t_R g83 ( .A(n_84), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_87), .Y(n_86) );
OAI22xp5_ASAP7_75t_L g87 ( .A1(n_88), .A2(n_89), .B1(n_90), .B2(n_91), .Y(n_87) );
CKINVDCx16_ASAP7_75t_R g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g91 ( .A(n_90), .Y(n_91) );
AOI22xp5_ASAP7_75t_L g92 ( .A1(n_93), .A2(n_95), .B1(n_96), .B2(n_206), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_93), .Y(n_206) );
INVx1_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_95), .A2(n_96), .B1(n_641), .B2(n_642), .Y(n_640) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
HB1xp67_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
NAND3xp33_ASAP7_75t_L g97 ( .A(n_98), .B(n_172), .C(n_192), .Y(n_97) );
HB1xp67_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx3_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_112), .Y(n_102) );
AND2x2_ASAP7_75t_L g196 ( .A(n_103), .B(n_181), .Y(n_196) );
AND2x2_ASAP7_75t_L g202 ( .A(n_103), .B(n_187), .Y(n_202) );
AND2x4_ASAP7_75t_L g204 ( .A(n_103), .B(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_111), .Y(n_103) );
INVx1_ASAP7_75t_L g130 ( .A(n_104), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
NAND2xp33_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
INVx2_ASAP7_75t_L g110 ( .A(n_106), .Y(n_110) );
INVx3_ASAP7_75t_L g116 ( .A(n_106), .Y(n_116) );
NAND2xp33_ASAP7_75t_L g122 ( .A(n_106), .B(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g139 ( .A(n_106), .Y(n_139) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_106), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_107), .B(n_137), .Y(n_136) );
INVxp67_ASAP7_75t_L g216 ( .A(n_107), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
OAI21xp5_ASAP7_75t_L g149 ( .A1(n_109), .A2(n_139), .B(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g129 ( .A(n_111), .B(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g148 ( .A(n_111), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g165 ( .A(n_111), .Y(n_165) );
AND2x4_ASAP7_75t_L g128 ( .A(n_112), .B(n_129), .Y(n_128) );
AND2x4_ASAP7_75t_L g132 ( .A(n_112), .B(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g176 ( .A(n_112), .B(n_164), .Y(n_176) );
AND2x4_ASAP7_75t_L g112 ( .A(n_113), .B(n_118), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g144 ( .A(n_114), .B(n_145), .Y(n_144) );
OR2x2_ASAP7_75t_L g167 ( .A(n_114), .B(n_168), .Y(n_167) );
AND2x4_ASAP7_75t_L g181 ( .A(n_114), .B(n_118), .Y(n_181) );
AND2x4_ASAP7_75t_L g187 ( .A(n_114), .B(n_188), .Y(n_187) );
AND2x4_ASAP7_75t_L g114 ( .A(n_115), .B(n_117), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_116), .B(n_121), .Y(n_120) );
INVxp67_ASAP7_75t_L g135 ( .A(n_116), .Y(n_135) );
NAND3xp33_ASAP7_75t_L g159 ( .A(n_117), .B(n_134), .C(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g168 ( .A(n_119), .Y(n_168) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_122), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_140), .Y(n_124) );
INVx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g199 ( .A(n_129), .B(n_181), .Y(n_199) );
AND2x4_ASAP7_75t_L g164 ( .A(n_130), .B(n_165), .Y(n_164) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x4_ASAP7_75t_L g171 ( .A(n_133), .B(n_166), .Y(n_171) );
AND2x4_ASAP7_75t_L g191 ( .A(n_133), .B(n_187), .Y(n_191) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_138), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
HB1xp67_ASAP7_75t_L g217 ( .A(n_137), .Y(n_217) );
INVx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx5_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_148), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
INVx1_ASAP7_75t_L g155 ( .A(n_146), .Y(n_155) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_147), .Y(n_213) );
INVx4_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx4_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AO21x2_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_159), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_164), .B(n_166), .Y(n_163) );
AND2x4_ASAP7_75t_L g180 ( .A(n_164), .B(n_181), .Y(n_180) );
AND2x4_ASAP7_75t_L g186 ( .A(n_164), .B(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g205 ( .A(n_167), .Y(n_205) );
INVx1_ASAP7_75t_L g188 ( .A(n_168), .Y(n_188) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx6_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
BUFx4f_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
BUFx12f_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
BUFx12f_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx4_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx8_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
BUFx3_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
BUFx3_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
BUFx8_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
BUFx3_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
BUFx10_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_210), .B(n_218), .Y(n_209) );
INVxp67_ASAP7_75t_SL g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g644 ( .A(n_211), .B(n_218), .Y(n_644) );
AOI211xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_214), .C(n_217), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_219), .B(n_222), .Y(n_218) );
OR2x2_ASAP7_75t_L g649 ( .A(n_219), .B(n_223), .Y(n_649) );
INVx1_ASAP7_75t_L g652 ( .A(n_219), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_219), .B(n_222), .Y(n_653) );
HB1xp67_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
HB1xp67_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
BUFx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_228), .Y(n_225) );
OAI21x1_ASAP7_75t_L g299 ( .A1(n_226), .A2(n_300), .B(n_308), .Y(n_299) );
AO31x2_ASAP7_75t_L g356 ( .A1(n_226), .A2(n_357), .A3(n_366), .B(n_367), .Y(n_356) );
AO31x2_ASAP7_75t_L g421 ( .A1(n_226), .A2(n_357), .A3(n_366), .B(n_367), .Y(n_421) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx3_ASAP7_75t_L g270 ( .A(n_227), .Y(n_270) );
INVx1_ASAP7_75t_L g273 ( .A(n_227), .Y(n_273) );
INVx3_ASAP7_75t_L g341 ( .A(n_227), .Y(n_341) );
OA21x2_ASAP7_75t_L g651 ( .A1(n_228), .A2(n_652), .B(n_653), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_229), .B(n_233), .Y(n_228) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_230), .B(n_303), .Y(n_302) );
OAI22x1_ASAP7_75t_L g357 ( .A1(n_230), .A2(n_358), .B1(n_362), .B2(n_363), .Y(n_357) );
INVx4_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_231), .A2(n_255), .B(n_258), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_231), .A2(n_301), .B1(n_302), .B2(n_305), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_231), .B(n_339), .Y(n_338) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_232), .Y(n_268) );
INVxp67_ASAP7_75t_L g324 ( .A(n_232), .Y(n_324) );
INVx1_ASAP7_75t_L g346 ( .A(n_232), .Y(n_346) );
INVx4_ASAP7_75t_L g376 ( .A(n_232), .Y(n_376) );
INVx3_ASAP7_75t_L g385 ( .A(n_232), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_232), .B(n_394), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_232), .B(n_397), .Y(n_396) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g310 ( .A(n_235), .Y(n_310) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx6_ASAP7_75t_L g257 ( .A(n_236), .Y(n_257) );
INVx3_ASAP7_75t_L g264 ( .A(n_236), .Y(n_264) );
INVx2_ASAP7_75t_L g307 ( .A(n_236), .Y(n_307) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NOR2x1p5_ASAP7_75t_L g239 ( .A(n_240), .B(n_541), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NOR3xp33_ASAP7_75t_L g241 ( .A(n_242), .B(n_459), .C(n_504), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_435), .Y(n_242) );
AOI211x1_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_371), .B(n_405), .C(n_426), .Y(n_243) );
OAI21xp5_ASAP7_75t_SL g244 ( .A1(n_245), .A2(n_295), .B(n_353), .Y(n_244) );
OR2x2_ASAP7_75t_L g450 ( .A(n_245), .B(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g537 ( .A(n_246), .B(n_538), .Y(n_537) );
AOI211xp5_ASAP7_75t_L g570 ( .A1(n_246), .A2(n_571), .B(n_572), .C(n_573), .Y(n_570) );
AND2x2_ASAP7_75t_L g582 ( .A(n_246), .B(n_451), .Y(n_582) );
AND2x2_ASAP7_75t_L g585 ( .A(n_246), .B(n_416), .Y(n_585) );
AND2x2_ASAP7_75t_L g615 ( .A(n_246), .B(n_440), .Y(n_615) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_271), .Y(n_246) );
INVx3_ASAP7_75t_L g425 ( .A(n_247), .Y(n_425) );
INVx2_ASAP7_75t_L g455 ( .A(n_247), .Y(n_455) );
AND2x2_ASAP7_75t_L g498 ( .A(n_247), .B(n_414), .Y(n_498) );
AND2x4_ASAP7_75t_L g247 ( .A(n_248), .B(n_253), .Y(n_247) );
NOR2x1_ASAP7_75t_L g269 ( .A(n_249), .B(n_270), .Y(n_269) );
INVx3_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_250), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx4_ASAP7_75t_L g277 ( .A(n_251), .Y(n_277) );
BUFx3_ASAP7_75t_L g294 ( .A(n_251), .Y(n_294) );
OAI21x1_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_261), .B(n_269), .Y(n_253) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g320 ( .A(n_257), .Y(n_320) );
INVx1_ASAP7_75t_L g323 ( .A(n_257), .Y(n_323) );
INVx2_ASAP7_75t_L g301 ( .A(n_259), .Y(n_301) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g266 ( .A(n_260), .Y(n_266) );
INVx2_ASAP7_75t_L g285 ( .A(n_260), .Y(n_285) );
INVx2_ASAP7_75t_L g365 ( .A(n_260), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_265), .B(n_267), .Y(n_261) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g289 ( .A(n_264), .Y(n_289) );
INVx2_ASAP7_75t_L g349 ( .A(n_264), .Y(n_349) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g279 ( .A(n_268), .Y(n_279) );
INVx2_ASAP7_75t_SL g290 ( .A(n_268), .Y(n_290) );
INVxp67_ASAP7_75t_L g312 ( .A(n_268), .Y(n_312) );
INVx2_ASAP7_75t_L g334 ( .A(n_270), .Y(n_334) );
INVx2_ASAP7_75t_SL g414 ( .A(n_271), .Y(n_414) );
AND2x2_ASAP7_75t_L g424 ( .A(n_271), .B(n_425), .Y(n_424) );
OAI21x1_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_278), .B(n_291), .Y(n_271) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_272), .A2(n_278), .B(n_291), .Y(n_463) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_273), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g380 ( .A(n_275), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g333 ( .A(n_277), .Y(n_333) );
AOI21x1_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_280), .B(n_286), .Y(n_278) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g361 ( .A(n_284), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_285), .A2(n_310), .B1(n_399), .B2(n_401), .Y(n_398) );
AOI21x1_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_288), .B(n_290), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_290), .B(n_329), .Y(n_330) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
NOR2xp67_ASAP7_75t_SL g367 ( .A(n_293), .B(n_368), .Y(n_367) );
INVx3_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OA21x2_ASAP7_75t_L g298 ( .A1(n_294), .A2(n_299), .B(n_313), .Y(n_298) );
OA21x2_ASAP7_75t_L g370 ( .A1(n_294), .A2(n_299), .B(n_313), .Y(n_370) );
NOR2x1_ASAP7_75t_SL g499 ( .A(n_295), .B(n_500), .Y(n_499) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_314), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_296), .B(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g576 ( .A(n_296), .B(n_553), .Y(n_576) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g445 ( .A(n_297), .B(n_336), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_297), .B(n_410), .Y(n_477) );
AND2x2_ASAP7_75t_L g618 ( .A(n_297), .B(n_356), .Y(n_618) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g419 ( .A(n_298), .Y(n_419) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_298), .Y(n_521) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_311), .B(n_312), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_310), .B(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_336), .Y(n_314) );
INVx1_ASAP7_75t_L g408 ( .A(n_315), .Y(n_408) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g354 ( .A(n_316), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g458 ( .A(n_316), .Y(n_458) );
INVxp67_ASAP7_75t_L g591 ( .A(n_316), .Y(n_591) );
AO21x2_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_325), .B(n_331), .Y(n_316) );
AO21x2_ASAP7_75t_L g432 ( .A1(n_317), .A2(n_325), .B(n_331), .Y(n_432) );
OAI21x1_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_321), .B(n_324), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_319), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g343 ( .A(n_323), .Y(n_343) );
OAI21x1_ASAP7_75t_SL g325 ( .A1(n_326), .A2(n_327), .B(n_330), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g335 ( .A(n_329), .Y(n_335) );
AOI21xp33_ASAP7_75t_SL g331 ( .A1(n_332), .A2(n_334), .B(n_335), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND3xp33_ASAP7_75t_SL g375 ( .A(n_334), .B(n_376), .C(n_377), .Y(n_375) );
NAND3xp33_ASAP7_75t_L g383 ( .A(n_334), .B(n_377), .C(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g369 ( .A(n_336), .B(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g410 ( .A(n_336), .Y(n_410) );
INVx1_ASAP7_75t_L g417 ( .A(n_336), .Y(n_417) );
INVx1_ASAP7_75t_L g635 ( .A(n_336), .Y(n_635) );
NAND2x1p5_ASAP7_75t_L g336 ( .A(n_337), .B(n_344), .Y(n_336) );
AND2x2_ASAP7_75t_L g472 ( .A(n_337), .B(n_344), .Y(n_472) );
OR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_342), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_339), .B(n_346), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g352 ( .A(n_340), .Y(n_352) );
INVx2_ASAP7_75t_L g377 ( .A(n_340), .Y(n_377) );
OA21x2_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_347), .B(n_350), .Y(n_344) );
INVx1_ASAP7_75t_L g362 ( .A(n_346), .Y(n_362) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g379 ( .A(n_349), .Y(n_379) );
INVx1_ASAP7_75t_L g366 ( .A(n_351), .Y(n_366) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_369), .Y(n_353) );
INVx1_ASAP7_75t_L g479 ( .A(n_354), .Y(n_479) );
INVx2_ASAP7_75t_L g434 ( .A(n_355), .Y(n_434) );
INVx1_ASAP7_75t_L g448 ( .A(n_355), .Y(n_448) );
AND2x2_ASAP7_75t_L g481 ( .A(n_355), .B(n_410), .Y(n_481) );
INVx3_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_369), .B(n_457), .Y(n_487) );
AND2x2_ASAP7_75t_L g590 ( .A(n_369), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g474 ( .A(n_370), .B(n_432), .Y(n_474) );
AND2x2_ASAP7_75t_L g589 ( .A(n_370), .B(n_472), .Y(n_589) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_372), .B(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g563 ( .A(n_372), .B(n_424), .Y(n_563) );
INVx2_ASAP7_75t_L g572 ( .A(n_372), .Y(n_572) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_387), .Y(n_372) );
INVx1_ASAP7_75t_L g412 ( .A(n_373), .Y(n_412) );
NOR2x1_ASAP7_75t_L g428 ( .A(n_373), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g440 ( .A(n_373), .B(n_388), .Y(n_440) );
INVx1_ASAP7_75t_L g452 ( .A(n_373), .Y(n_452) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_373), .Y(n_466) );
INVx1_ASAP7_75t_L g497 ( .A(n_373), .Y(n_497) );
INVx2_ASAP7_75t_L g503 ( .A(n_373), .Y(n_503) );
AND2x2_ASAP7_75t_L g546 ( .A(n_373), .B(n_425), .Y(n_546) );
OR2x6_ASAP7_75t_L g373 ( .A(n_374), .B(n_382), .Y(n_373) );
OAI21x1_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_378), .B(n_380), .Y(n_374) );
NOR2xp33_ASAP7_75t_SL g399 ( .A(n_376), .B(n_400), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_376), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g390 ( .A(n_377), .Y(n_390) );
NOR2xp67_ASAP7_75t_L g382 ( .A(n_383), .B(n_386), .Y(n_382) );
INVx3_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g502 ( .A(n_387), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g413 ( .A(n_388), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g429 ( .A(n_388), .Y(n_429) );
OR2x2_ASAP7_75t_L g462 ( .A(n_388), .B(n_463), .Y(n_462) );
INVxp67_ASAP7_75t_L g540 ( .A(n_388), .Y(n_540) );
INVx1_ASAP7_75t_L g574 ( .A(n_388), .Y(n_574) );
AO21x2_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .B(n_403), .Y(n_388) );
NAND3xp33_ASAP7_75t_SL g391 ( .A(n_392), .B(n_395), .C(n_398), .Y(n_391) );
OAI32xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_409), .A3(n_411), .B1(n_415), .B2(n_422), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g605 ( .A(n_408), .B(n_477), .Y(n_605) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
AND2x2_ASAP7_75t_L g507 ( .A(n_412), .B(n_508), .Y(n_507) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_412), .Y(n_548) );
AND2x4_ASAP7_75t_L g545 ( .A(n_413), .B(n_546), .Y(n_545) );
BUFx3_ASAP7_75t_L g556 ( .A(n_413), .Y(n_556) );
INVx1_ASAP7_75t_L g517 ( .A(n_414), .Y(n_517) );
OR2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_418), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g511 ( .A(n_417), .Y(n_511) );
INVx1_ASAP7_75t_L g578 ( .A(n_417), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
AND2x4_ASAP7_75t_L g431 ( .A(n_419), .B(n_432), .Y(n_431) );
INVxp67_ASAP7_75t_SL g601 ( .A(n_419), .Y(n_601) );
INVx1_ASAP7_75t_L g561 ( .A(n_420), .Y(n_561) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g457 ( .A(n_421), .B(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g536 ( .A(n_421), .B(n_432), .Y(n_536) );
OR2x2_ASAP7_75t_L g553 ( .A(n_421), .B(n_432), .Y(n_553) );
INVx1_ASAP7_75t_L g569 ( .A(n_423), .Y(n_569) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x4_ASAP7_75t_L g427 ( .A(n_424), .B(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g438 ( .A(n_424), .Y(n_438) );
AND2x2_ASAP7_75t_L g501 ( .A(n_424), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g516 ( .A(n_425), .Y(n_516) );
AND2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_430), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_427), .A2(n_587), .B1(n_588), .B2(n_590), .Y(n_586) );
INVx2_ASAP7_75t_L g599 ( .A(n_427), .Y(n_599) );
INVx2_ASAP7_75t_L g568 ( .A(n_428), .Y(n_568) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_433), .Y(n_430) );
AND2x4_ASAP7_75t_SL g447 ( .A(n_431), .B(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_431), .B(n_481), .Y(n_495) );
BUFx3_ASAP7_75t_L g529 ( .A(n_431), .Y(n_529) );
INVx1_ASAP7_75t_L g491 ( .A(n_433), .Y(n_491) );
AND2x2_ASAP7_75t_L g562 ( .A(n_433), .B(n_445), .Y(n_562) );
AND2x2_ASAP7_75t_L g583 ( .A(n_433), .B(n_474), .Y(n_583) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g443 ( .A(n_434), .Y(n_443) );
AND2x2_ASAP7_75t_L g526 ( .A(n_434), .B(n_471), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_441), .B(n_449), .Y(n_435) );
INVx2_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g579 ( .A(n_437), .Y(n_579) );
OR2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_440), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_440), .B(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_442), .B(n_446), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_443), .B(n_585), .Y(n_609) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_446), .A2(n_450), .B1(n_453), .B2(n_456), .Y(n_449) );
INVx2_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
NAND2xp67_ASAP7_75t_L g509 ( .A(n_447), .B(n_510), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_447), .A2(n_631), .B1(n_637), .B2(n_638), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_448), .B(n_623), .Y(n_629) );
OR2x2_ASAP7_75t_L g514 ( .A(n_451), .B(n_515), .Y(n_514) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_451), .Y(n_611) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g488 ( .A(n_452), .B(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g567 ( .A(n_454), .B(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g571 ( .A(n_454), .Y(n_571) );
AND2x2_ASAP7_75t_L g573 ( .A(n_454), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g461 ( .A(n_455), .B(n_462), .Y(n_461) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_455), .Y(n_484) );
AND2x2_ASAP7_75t_L g523 ( .A(n_455), .B(n_497), .Y(n_523) );
AND2x2_ASAP7_75t_L g555 ( .A(n_457), .B(n_535), .Y(n_555) );
AND2x4_ASAP7_75t_L g588 ( .A(n_457), .B(n_589), .Y(n_588) );
INVx3_ASAP7_75t_L g606 ( .A(n_457), .Y(n_606) );
BUFx3_ASAP7_75t_L g637 ( .A(n_457), .Y(n_637) );
INVx1_ASAP7_75t_L g522 ( .A(n_458), .Y(n_522) );
OAI211xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_467), .B(n_482), .C(n_493), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_464), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_461), .A2(n_613), .B1(n_614), .B2(n_616), .Y(n_612) );
INVx1_ASAP7_75t_L g485 ( .A(n_462), .Y(n_485) );
INVx2_ASAP7_75t_L g489 ( .A(n_462), .Y(n_489) );
BUFx2_ASAP7_75t_L g508 ( .A(n_463), .Y(n_508) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g604 ( .A(n_466), .B(n_489), .Y(n_604) );
NOR3xp33_ASAP7_75t_L g467 ( .A(n_468), .B(n_475), .C(n_478), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_473), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g535 ( .A(n_471), .Y(n_535) );
INVx2_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g492 ( .A(n_473), .Y(n_492) );
INVx1_ASAP7_75t_L g525 ( .A(n_473), .Y(n_525) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVxp67_ASAP7_75t_L g560 ( .A(n_477), .Y(n_560) );
NAND2xp33_ASAP7_75t_SL g478 ( .A(n_479), .B(n_480), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_479), .B(n_539), .Y(n_584) );
NOR2x1_ASAP7_75t_R g528 ( .A(n_480), .B(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_481), .B(n_520), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_486), .B1(n_488), .B2(n_490), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g638 ( .A(n_488), .B(n_633), .Y(n_638) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_491), .B(n_601), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_496), .B(n_499), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
INVx2_ASAP7_75t_L g624 ( .A(n_498), .Y(n_624) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OAI211xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_509), .B(n_512), .C(n_527), .Y(n_504) );
INVxp67_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g533 ( .A(n_508), .Y(n_533) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g551 ( .A(n_511), .B(n_552), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_518), .B1(n_523), .B2(n_524), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NOR2xp67_ASAP7_75t_SL g597 ( .A(n_515), .B(n_574), .Y(n_597) );
OR2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g550 ( .A(n_516), .Y(n_550) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
INVx1_ASAP7_75t_L g617 ( .A(n_522), .Y(n_617) );
NAND2x2_ASAP7_75t_L g625 ( .A(n_523), .B(n_556), .Y(n_625) );
OAI21xp33_ASAP7_75t_L g554 ( .A1(n_524), .A2(n_555), .B(n_556), .Y(n_554) );
AND2x4_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_530), .B1(n_534), .B2(n_537), .Y(n_527) );
INVx2_ASAP7_75t_L g622 ( .A(n_529), .Y(n_622) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVxp67_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
AND2x2_ASAP7_75t_L g577 ( .A(n_536), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g626 ( .A(n_536), .Y(n_626) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_592), .Y(n_541) );
NOR2x1p5_ASAP7_75t_L g542 ( .A(n_543), .B(n_564), .Y(n_542) );
NAND3xp33_ASAP7_75t_SL g543 ( .A(n_544), .B(n_554), .C(n_557), .Y(n_543) );
OAI21xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_547), .B(n_551), .Y(n_544) );
INVx2_ASAP7_75t_L g628 ( .A(n_545), .Y(n_628) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g633 ( .A(n_550), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OAI21xp33_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_562), .B(n_563), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
NAND2x1p5_ASAP7_75t_L g596 ( .A(n_562), .B(n_597), .Y(n_596) );
NAND2x1p5_ASAP7_75t_L g564 ( .A(n_565), .B(n_580), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_575), .B1(n_577), .B2(n_579), .Y(n_565) );
AO21x1_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_569), .B(n_570), .Y(n_566) );
OR2x2_ASAP7_75t_L g623 ( .A(n_568), .B(n_624), .Y(n_623) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_573), .Y(n_587) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_586), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_583), .B1(n_584), .B2(n_585), .Y(n_581) );
NOR2x1_ASAP7_75t_L g592 ( .A(n_593), .B(n_619), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_607), .Y(n_593) );
NOR3xp33_ASAP7_75t_L g594 ( .A(n_595), .B(n_598), .C(n_602), .Y(n_594) );
INVxp67_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_599), .A2(n_603), .B1(n_605), .B2(n_606), .Y(n_602) );
INVx1_ASAP7_75t_L g613 ( .A(n_601), .Y(n_613) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_SL g636 ( .A(n_604), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_610), .B(n_612), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVxp67_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_616), .B(n_628), .Y(n_627) );
NAND2x1p5_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_630), .Y(n_619) );
NOR3xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_627), .C(n_629), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_623), .B1(n_625), .B2(n_626), .Y(n_621) );
NOR2xp67_ASAP7_75t_L g631 ( .A(n_632), .B(n_636), .Y(n_631) );
INVx2_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI222xp33_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_642), .B1(n_643), .B2(n_645), .C1(n_648), .C2(n_650), .Y(n_639) );
CKINVDCx5p33_ASAP7_75t_R g642 ( .A(n_641), .Y(n_642) );
INVx1_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
BUFx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
endmodule