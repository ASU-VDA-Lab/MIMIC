module fake_netlist_1_442_n_44 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_44);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_44;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
BUFx2_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_4), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_5), .Y(n_13) );
INVx5_ASAP7_75t_L g14 ( .A(n_6), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_2), .B(n_6), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_8), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_1), .Y(n_17) );
AND3x1_ASAP7_75t_L g18 ( .A(n_15), .B(n_0), .C(n_1), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_11), .B(n_0), .Y(n_19) );
BUFx12f_ASAP7_75t_L g20 ( .A(n_11), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_12), .B(n_2), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_14), .Y(n_22) );
NAND2xp5_ASAP7_75t_SL g23 ( .A(n_14), .B(n_3), .Y(n_23) );
OAI22x1_ASAP7_75t_L g24 ( .A1(n_18), .A2(n_17), .B1(n_13), .B2(n_15), .Y(n_24) );
AND2x4_ASAP7_75t_L g25 ( .A(n_18), .B(n_14), .Y(n_25) );
OAI22xp33_ASAP7_75t_SL g26 ( .A1(n_19), .A2(n_14), .B1(n_16), .B2(n_7), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_22), .Y(n_27) );
BUFx3_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
OAI31xp33_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_23), .A3(n_21), .B(n_22), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_27), .Y(n_30) );
AOI22xp33_ASAP7_75t_L g31 ( .A1(n_28), .A2(n_25), .B1(n_24), .B2(n_20), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_31), .B(n_20), .Y(n_33) );
AOI21xp33_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_29), .B(n_28), .Y(n_34) );
OR2x2_ASAP7_75t_L g35 ( .A(n_32), .B(n_28), .Y(n_35) );
NAND2xp33_ASAP7_75t_L g36 ( .A(n_35), .B(n_30), .Y(n_36) );
O2A1O1Ixp33_ASAP7_75t_L g37 ( .A1(n_34), .A2(n_29), .B(n_28), .C(n_30), .Y(n_37) );
AO22x2_ASAP7_75t_L g38 ( .A1(n_33), .A2(n_28), .B1(n_29), .B2(n_7), .Y(n_38) );
AND2x2_ASAP7_75t_L g39 ( .A(n_38), .B(n_14), .Y(n_39) );
INVxp67_ASAP7_75t_SL g40 ( .A(n_36), .Y(n_40) );
NOR3xp33_ASAP7_75t_L g41 ( .A(n_37), .B(n_14), .C(n_5), .Y(n_41) );
OAI22xp5_ASAP7_75t_L g42 ( .A1(n_40), .A2(n_38), .B1(n_3), .B2(n_10), .Y(n_42) );
NAND2xp5_ASAP7_75t_L g43 ( .A(n_39), .B(n_9), .Y(n_43) );
OAI22xp5_ASAP7_75t_L g44 ( .A1(n_42), .A2(n_39), .B1(n_41), .B2(n_43), .Y(n_44) );
endmodule