module fake_jpeg_1199_n_188 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_188);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_24),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

BUFx4f_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_68),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_60),
.B1(n_48),
.B2(n_61),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_77),
.A2(n_83),
.B1(n_65),
.B2(n_48),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_84),
.Y(n_91)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_56),
.B1(n_65),
.B2(n_47),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_78),
.B1(n_81),
.B2(n_74),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_47),
.B1(n_53),
.B2(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_89),
.B1(n_97),
.B2(n_100),
.Y(n_105)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_68),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_90),
.B(n_96),
.Y(n_115)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_52),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_80),
.A2(n_65),
.B1(n_52),
.B2(n_64),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_54),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_55),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_76),
.A2(n_65),
.B1(n_62),
.B2(n_53),
.Y(n_100)
);

NOR3xp33_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_64),
.C(n_59),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_70),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_89),
.B(n_93),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_121),
.C(n_43),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_118),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_54),
.B1(n_59),
.B2(n_62),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_108),
.B1(n_114),
.B2(n_58),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_95),
.B1(n_89),
.B2(n_93),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_92),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_57),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_57),
.B1(n_55),
.B2(n_49),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_49),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_46),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_70),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_39),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_70),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_129),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_124),
.A2(n_126),
.B1(n_133),
.B2(n_4),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_58),
.C(n_45),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_131),
.C(n_135),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_44),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_132),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_9),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_119),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_116),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_137),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_42),
.C(n_41),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_40),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_109),
.B1(n_103),
.B2(n_117),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_134),
.A2(n_135),
.B1(n_120),
.B2(n_5),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_106),
.A2(n_38),
.B1(n_37),
.B2(n_36),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_113),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_102),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_120),
.B1(n_112),
.B2(n_6),
.Y(n_145)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_33),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_30),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_SL g142 ( 
.A1(n_122),
.A2(n_127),
.A3(n_123),
.B1(n_132),
.B2(n_136),
.C1(n_125),
.C2(n_140),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_142),
.B(n_149),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_133),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_143),
.B(n_144),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_133),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_152),
.B1(n_155),
.B2(n_153),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_150),
.Y(n_160)
);

NOR3xp33_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_156),
.C(n_10),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_4),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_134),
.A2(n_5),
.B(n_6),
.Y(n_153)
);

AOI32xp33_ASAP7_75t_L g166 ( 
.A1(n_153),
.A2(n_154),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_7),
.B(n_8),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_138),
.A2(n_126),
.B1(n_10),
.B2(n_11),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_158),
.A2(n_162),
.B1(n_15),
.B2(n_16),
.Y(n_174)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_159),
.A2(n_163),
.B1(n_164),
.B2(n_166),
.Y(n_173)
);

AOI221xp5_ASAP7_75t_L g169 ( 
.A1(n_161),
.A2(n_154),
.B1(n_148),
.B2(n_157),
.C(n_156),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_147),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_164),
.A2(n_146),
.B1(n_155),
.B2(n_157),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_169),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_165),
.A2(n_150),
.B(n_27),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_172),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_25),
.C(n_13),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_174),
.C(n_163),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_160),
.A2(n_12),
.B1(n_15),
.B2(n_16),
.Y(n_172)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_175),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_170),
.C(n_173),
.Y(n_177)
);

NAND4xp25_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_168),
.C(n_176),
.D(n_178),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_179),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_172),
.C(n_159),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_180),
.B1(n_167),
.B2(n_19),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_17),
.C(n_18),
.Y(n_184)
);

MAJx2_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_19),
.C(n_20),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_20),
.B(n_21),
.Y(n_186)
);

AOI221xp5_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.C(n_24),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_22),
.Y(n_188)
);


endmodule