module fake_jpeg_11052_n_155 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_155);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_155;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_29),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_23),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

INVx11_ASAP7_75t_SL g55 ( 
.A(n_30),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_16),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_24),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_7),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_19),
.B1(n_46),
.B2(n_45),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_74),
.A2(n_51),
.B1(n_60),
.B2(n_64),
.Y(n_87)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_0),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_76),
.B(n_80),
.Y(n_83)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_55),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_55),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_66),
.B(n_4),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_62),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_49),
.B1(n_56),
.B2(n_52),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_66),
.B(n_69),
.C(n_67),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_95),
.B(n_3),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_90),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_59),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_94),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_58),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_49),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_111),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_87),
.A2(n_56),
.B1(n_60),
.B2(n_64),
.Y(n_98)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_105),
.B1(n_107),
.B2(n_110),
.Y(n_123)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_54),
.B(n_20),
.C(n_21),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_3),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_106),
.B(n_109),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_18),
.B1(n_42),
.B2(n_39),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_4),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_17),
.B1(n_35),
.B2(n_34),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_84),
.A2(n_5),
.B(n_6),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_12),
.C(n_32),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_114),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_48),
.B1(n_28),
.B2(n_27),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_22),
.B1(n_10),
.B2(n_11),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_82),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_91),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_9),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_103),
.B(n_5),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_108),
.B(n_6),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_26),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_122),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_106),
.B(n_7),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_125),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_99),
.B(n_8),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_101),
.B(n_8),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_100),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_130),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_113),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_133),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_132),
.A2(n_123),
.B1(n_120),
.B2(n_124),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_105),
.B(n_10),
.Y(n_133)
);

AO22x1_ASAP7_75t_L g136 ( 
.A1(n_124),
.A2(n_11),
.B1(n_131),
.B2(n_118),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_136),
.B(n_138),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_128),
.C(n_126),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_139),
.A2(n_143),
.B(n_142),
.Y(n_146)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

INVxp67_ASAP7_75t_SL g145 ( 
.A(n_141),
.Y(n_145)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_146),
.B(n_139),
.Y(n_148)
);

NAND4xp25_ASAP7_75t_SL g147 ( 
.A(n_136),
.B(n_127),
.C(n_132),
.D(n_140),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_147),
.B(n_142),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_148),
.B(n_149),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_145),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_148),
.B1(n_150),
.B2(n_144),
.Y(n_153)
);

NAND3xp33_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_135),
.C(n_134),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_137),
.Y(n_155)
);


endmodule