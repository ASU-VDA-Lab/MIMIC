module real_jpeg_2739_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_284, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_284;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_110;
wire n_61;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_70;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_41;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_167;
wire n_128;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

INVx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_1),
.A2(n_73),
.B1(n_74),
.B2(n_163),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_1),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_1),
.A2(n_62),
.B1(n_63),
.B2(n_163),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_1),
.A2(n_44),
.B1(n_45),
.B2(n_163),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_1),
.A2(n_31),
.B1(n_34),
.B2(n_163),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_3),
.A2(n_73),
.B1(n_74),
.B2(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_3),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_3),
.A2(n_62),
.B1(n_63),
.B2(n_134),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_134),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_3),
.A2(n_31),
.B1(n_34),
.B2(n_134),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_4),
.A2(n_44),
.B1(n_45),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_4),
.A2(n_53),
.B1(n_62),
.B2(n_63),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_4),
.A2(n_31),
.B1(n_34),
.B2(n_53),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_5),
.A2(n_31),
.B1(n_34),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_5),
.A2(n_38),
.B1(n_62),
.B2(n_63),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_5),
.A2(n_38),
.B1(n_44),
.B2(n_45),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_5),
.A2(n_38),
.B1(n_73),
.B2(n_74),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_6),
.A2(n_44),
.B1(n_45),
.B2(n_51),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_6),
.A2(n_51),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_6),
.A2(n_31),
.B1(n_34),
.B2(n_51),
.Y(n_151)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_8),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_9),
.A2(n_73),
.B1(n_74),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_9),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_9),
.A2(n_62),
.B1(n_63),
.B2(n_80),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_80),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_9),
.A2(n_31),
.B1(n_34),
.B2(n_80),
.Y(n_223)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_12),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_12),
.B(n_82),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_12),
.B(n_62),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_12),
.A2(n_73),
.B(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_12),
.B(n_34),
.C(n_47),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_12),
.A2(n_44),
.B1(n_45),
.B2(n_154),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_12),
.B(n_110),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_12),
.B(n_28),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_12),
.B(n_55),
.Y(n_238)
);

AOI21xp33_ASAP7_75t_L g253 ( 
.A1(n_12),
.A2(n_62),
.B(n_187),
.Y(n_253)
);

BUFx10_ASAP7_75t_L g76 ( 
.A(n_13),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_14),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_14),
.A2(n_33),
.B1(n_73),
.B2(n_74),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_14),
.A2(n_33),
.B1(n_44),
.B2(n_45),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_14),
.A2(n_33),
.B1(n_62),
.B2(n_63),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_137),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_135),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_113),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_19),
.B(n_113),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_84),
.B2(n_85),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_56),
.C(n_70),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_22),
.A2(n_23),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_40),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_35),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_26),
.A2(n_39),
.B(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_34),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_27),
.A2(n_30),
.B(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_27),
.A2(n_36),
.B(n_151),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_27),
.A2(n_90),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_28),
.B(n_37),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_28),
.A2(n_39),
.B1(n_126),
.B2(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_28),
.A2(n_39),
.B1(n_154),
.B2(n_234),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_28),
.A2(n_39),
.B1(n_234),
.B2(n_237),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_30),
.A2(n_90),
.B(n_127),
.Y(n_189)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_31),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_34),
.B(n_232),
.Y(n_231)
);

INVxp33_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_40),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_50),
.B1(n_52),
.B2(n_54),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_41),
.A2(n_52),
.B(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_41),
.A2(n_92),
.B(n_105),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_41),
.A2(n_54),
.B1(n_183),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_42),
.B(n_93),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_42),
.A2(n_104),
.B(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_42),
.A2(n_55),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_42),
.A2(n_55),
.B1(n_220),
.B2(n_226),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_49),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_43)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_45),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_L g188 ( 
.A(n_44),
.B(n_58),
.C(n_63),
.Y(n_188)
);

CKINVDCx6p67_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_45),
.A2(n_59),
.B(n_186),
.C(n_188),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_45),
.B(n_216),
.Y(n_215)
);

BUFx4f_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_49),
.B(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_50),
.A2(n_54),
.B(n_107),
.Y(n_128)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_55),
.B(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_56),
.B(n_70),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_61),
.B(n_65),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_57),
.A2(n_68),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_57),
.A2(n_68),
.B1(n_174),
.B2(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_59),
.B1(n_62),
.B2(n_63),
.Y(n_69)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_61),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_63),
.B1(n_76),
.B2(n_77),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_62),
.B(n_74),
.C(n_77),
.Y(n_155)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_63),
.A2(n_76),
.B(n_153),
.C(n_155),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_66),
.B(n_110),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_67),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_67),
.A2(n_110),
.B1(n_158),
.B2(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_68),
.A2(n_130),
.B(n_131),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_68),
.A2(n_157),
.B(n_159),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_79),
.B(n_81),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_71),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_71),
.A2(n_78),
.B1(n_79),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_71),
.A2(n_78),
.B1(n_133),
.B2(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_71),
.A2(n_78),
.B1(n_162),
.B2(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_78),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_74),
.B(n_154),
.Y(n_153)
);

BUFx4f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_100),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_83),
.Y(n_98)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_101),
.B2(n_102),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_94),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_91),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_89),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_91),
.B1(n_95),
.B2(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_90),
.A2(n_125),
.B(n_127),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_91),
.Y(n_119)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_108),
.B(n_112),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_108),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_110),
.B(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.C(n_120),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_114),
.A2(n_117),
.B1(n_118),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_114),
.Y(n_167)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_120),
.A2(n_121),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_129),
.C(n_132),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_123),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_124),
.B(n_128),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_132),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_168),
.B(n_282),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_164),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_139),
.B(n_164),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.C(n_145),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_140),
.B(n_143),
.Y(n_265)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_145),
.B(n_265),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_156),
.C(n_161),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_146),
.A2(n_147),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_152),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_148),
.A2(n_149),
.B1(n_152),
.B2(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_152),
.Y(n_208)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_156),
.B(n_161),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

AOI321xp33_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_263),
.A3(n_274),
.B1(n_280),
.B2(n_281),
.C(n_284),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_209),
.B(n_262),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_190),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_171),
.B(n_190),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_181),
.C(n_184),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_172),
.B(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_177),
.C(n_180),
.Y(n_205)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_181),
.B(n_184),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_189),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_185),
.B(n_189),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_202),
.B2(n_203),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_191),
.B(n_204),
.C(n_207),
.Y(n_275)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_193),
.B(n_197),
.C(n_201),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_200),
.B2(n_201),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_257),
.B(n_261),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_247),
.B(n_256),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_228),
.B(n_246),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_221),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_221),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_214),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_225),
.C(n_227),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_223),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_226),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_240),
.B(n_245),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_235),
.B(n_239),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_238),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_237),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_244),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_248),
.B(n_249),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_252),
.C(n_254),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_260),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_266),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_271),
.C(n_273),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_267),
.A2(n_268),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_271),
.A2(n_272),
.B1(n_273),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_273),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_276),
.Y(n_280)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);


endmodule