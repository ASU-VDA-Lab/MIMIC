module fake_jpeg_2007_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx12_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_1),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_19),
.Y(n_31)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_9),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_18),
.A2(n_15),
.B1(n_11),
.B2(n_10),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_5),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_14),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_22),
.Y(n_32)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_15),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_8),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_27),
.Y(n_34)
);

AOI21xp33_ASAP7_75t_L g27 ( 
.A1(n_19),
.A2(n_8),
.B(n_11),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_29),
.A2(n_17),
.B1(n_18),
.B2(n_10),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_10),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_31),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_40),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_20),
.C(n_21),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_29),
.C(n_28),
.Y(n_43)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_37),
.C(n_33),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_SL g46 ( 
.A(n_41),
.B(n_36),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_34),
.B1(n_40),
.B2(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_48),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_34),
.C(n_46),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_49),
.C(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_44),
.B(n_35),
.Y(n_54)
);

AOI221xp5_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_26),
.B1(n_38),
.B2(n_39),
.C(n_45),
.Y(n_55)
);


endmodule