module fake_jpeg_9033_n_254 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_254);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_SL g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_39),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_30),
.B(n_0),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_30),
.B1(n_18),
.B2(n_19),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_39),
.B1(n_19),
.B2(n_18),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_37),
.B1(n_36),
.B2(n_38),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_46),
.B1(n_51),
.B2(n_24),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_20),
.B1(n_29),
.B2(n_17),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_52),
.B1(n_33),
.B2(n_25),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_17),
.B1(n_29),
.B2(n_26),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_24),
.B1(n_26),
.B2(n_20),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_36),
.B1(n_21),
.B2(n_27),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_57),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_54),
.Y(n_75)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_50),
.A2(n_38),
.B1(n_27),
.B2(n_21),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_59),
.A2(n_70),
.B1(n_78),
.B2(n_49),
.Y(n_91)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_63),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_51),
.A2(n_28),
.B1(n_18),
.B2(n_19),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_62),
.B(n_71),
.Y(n_100)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_58),
.B(n_23),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_68),
.Y(n_104)
);

CKINVDCx12_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_56),
.B1(n_55),
.B2(n_49),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_18),
.B1(n_19),
.B2(n_23),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_67),
.A2(n_79),
.B1(n_32),
.B2(n_48),
.Y(n_96)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_74),
.Y(n_105)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_12),
.C(n_13),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_73),
.Y(n_107)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_41),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_77),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_44),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_33),
.B1(n_32),
.B2(n_22),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_41),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_82),
.Y(n_89)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_41),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_85),
.Y(n_99)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_84),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_56),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_87),
.A2(n_88),
.B1(n_101),
.B2(n_107),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_33),
.B1(n_56),
.B2(n_49),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_0),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_94),
.B(n_64),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_109),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_1),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_96),
.B(n_35),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_74),
.A2(n_78),
.B1(n_70),
.B2(n_75),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_98),
.A2(n_108),
.B1(n_111),
.B2(n_48),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_37),
.B1(n_35),
.B2(n_34),
.Y(n_101)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_68),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_85),
.A2(n_11),
.B1(n_14),
.B2(n_3),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_134),
.B(n_100),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_83),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_115),
.B(n_118),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_93),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_116),
.B(n_122),
.Y(n_148)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_104),
.B(n_62),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_77),
.B(n_61),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_119),
.A2(n_136),
.B(n_37),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_82),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_120),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_125),
.B1(n_137),
.B2(n_108),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_84),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_73),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_124),
.C(n_130),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_35),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_93),
.Y(n_128)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_131),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_109),
.C(n_103),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_35),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_34),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_90),
.B(n_94),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_34),
.Y(n_135)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_88),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_107),
.B1(n_97),
.B2(n_100),
.Y(n_138)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_141),
.B(n_151),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_136),
.A2(n_87),
.B1(n_94),
.B2(n_101),
.Y(n_142)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_142),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_96),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_147),
.C(n_123),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_144),
.B(n_135),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_133),
.A2(n_106),
.B(n_16),
.Y(n_146)
);

HAxp5_ASAP7_75t_SL g182 ( 
.A(n_146),
.B(n_149),
.CON(n_182),
.SN(n_182)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_102),
.C(n_108),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_16),
.B(n_102),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_150),
.A2(n_157),
.B1(n_128),
.B2(n_116),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_134),
.A2(n_32),
.B(n_16),
.Y(n_151)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_131),
.A2(n_37),
.A3(n_48),
.B1(n_102),
.B2(n_16),
.Y(n_152)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_110),
.B1(n_37),
.B2(n_1),
.Y(n_154)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_121),
.A2(n_37),
.B1(n_2),
.B2(n_1),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_156),
.Y(n_179)
);

AOI22x1_ASAP7_75t_SL g157 ( 
.A1(n_119),
.A2(n_7),
.B1(n_13),
.B2(n_3),
.Y(n_157)
);

A2O1A1O1Ixp25_ASAP7_75t_L g161 ( 
.A1(n_120),
.A2(n_7),
.B(n_13),
.C(n_3),
.D(n_4),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_112),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_8),
.B1(n_12),
.B2(n_4),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_117),
.Y(n_165)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_115),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_169),
.C(n_180),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_167),
.B(n_173),
.Y(n_198)
);

NAND3xp33_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_132),
.C(n_113),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_184),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_113),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_174),
.A2(n_183),
.B1(n_181),
.B2(n_186),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_140),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_176),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_153),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_160),
.B(n_148),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_122),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_153),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_1),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_178),
.A2(n_142),
.B1(n_162),
.B2(n_144),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_187),
.A2(n_189),
.B1(n_197),
.B2(n_202),
.Y(n_215)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_178),
.A2(n_162),
.B1(n_163),
.B2(n_158),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_190),
.B(n_167),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_172),
.B(n_141),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_6),
.C(n_8),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_170),
.A2(n_138),
.B1(n_156),
.B2(n_160),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_192),
.A2(n_195),
.B1(n_196),
.B2(n_5),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_166),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_170),
.A2(n_163),
.B1(n_158),
.B2(n_147),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_186),
.A2(n_154),
.B1(n_143),
.B2(n_152),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_179),
.A2(n_145),
.B1(n_149),
.B2(n_161),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_184),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_185),
.A2(n_146),
.B1(n_145),
.B2(n_151),
.Y(n_200)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_181),
.A2(n_127),
.B1(n_2),
.B2(n_6),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_194),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_189),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_199),
.A2(n_185),
.B1(n_182),
.B2(n_169),
.Y(n_206)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_204),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_208),
.A2(n_210),
.B(n_211),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_209),
.B(n_203),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_196),
.A2(n_182),
.B(n_168),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_L g211 ( 
.A1(n_204),
.A2(n_172),
.B1(n_180),
.B2(n_2),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_213),
.A2(n_216),
.B1(n_202),
.B2(n_197),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_198),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_187),
.A2(n_9),
.B1(n_11),
.B2(n_14),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_218),
.A2(n_219),
.B(n_208),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_217),
.A2(n_192),
.B1(n_201),
.B2(n_191),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_220),
.A2(n_215),
.B1(n_216),
.B2(n_212),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_188),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_222),
.B(n_226),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_224),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_213),
.B(n_193),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_228),
.C(n_214),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_203),
.C(n_195),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_225),
.A2(n_217),
.B1(n_210),
.B2(n_212),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_229),
.A2(n_220),
.B1(n_228),
.B2(n_227),
.Y(n_241)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_230),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_233),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_226),
.Y(n_233)
);

NAND2xp33_ASAP7_75t_SL g234 ( 
.A(n_221),
.B(n_215),
.Y(n_234)
);

INVxp33_ASAP7_75t_L g242 ( 
.A(n_234),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_221),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_238),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_223),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_239),
.B(n_241),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_237),
.A2(n_230),
.B(n_236),
.Y(n_243)
);

AOI21xp33_ASAP7_75t_L g248 ( 
.A1(n_243),
.A2(n_240),
.B(n_242),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_234),
.C(n_233),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_229),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_247),
.A2(n_248),
.B(n_245),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_246),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_249),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_242),
.C(n_9),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_14),
.C(n_250),
.Y(n_253)
);

BUFx24_ASAP7_75t_SL g254 ( 
.A(n_253),
.Y(n_254)
);


endmodule