module fake_jpeg_1878_n_375 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_375);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_375;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_331;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_SL g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx2_ASAP7_75t_R g47 ( 
.A(n_27),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_47),
.B(n_63),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_49),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_19),
.B(n_7),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_51),
.B(n_57),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_52),
.Y(n_149)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_19),
.B(n_7),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_16),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_58),
.B(n_59),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_21),
.B(n_15),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g145 ( 
.A(n_60),
.Y(n_145)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_62),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_65),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_21),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_76),
.Y(n_115)
);

BUFx8_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_75),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_26),
.Y(n_76)
);

HAxp5_ASAP7_75t_SL g77 ( 
.A(n_33),
.B(n_0),
.CON(n_77),
.SN(n_77)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_0),
.B(n_1),
.Y(n_97)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_26),
.B(n_10),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_87),
.Y(n_118)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_90),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_89),
.Y(n_119)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_25),
.B(n_12),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_92),
.Y(n_121)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_17),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_17),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_93),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_94),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_28),
.B(n_10),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_95),
.B(n_12),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_97),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_48),
.A2(n_33),
.B1(n_23),
.B2(n_22),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_100),
.A2(n_47),
.B1(n_93),
.B2(n_68),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_89),
.A2(n_39),
.B1(n_44),
.B2(n_31),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_102),
.A2(n_106),
.B1(n_130),
.B2(n_136),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_50),
.A2(n_44),
.B1(n_36),
.B2(n_37),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_56),
.A2(n_42),
.B1(n_34),
.B2(n_32),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_109),
.A2(n_132),
.B1(n_9),
.B2(n_4),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_60),
.A2(n_42),
.B1(n_34),
.B2(n_28),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_110),
.A2(n_152),
.B1(n_80),
.B2(n_90),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_38),
.C(n_29),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_111),
.B(n_139),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_49),
.B(n_38),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_131),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_88),
.A2(n_37),
.B1(n_36),
.B2(n_29),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g131 ( 
.A(n_88),
.B(n_71),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_62),
.A2(n_45),
.B1(n_23),
.B2(n_22),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_71),
.A2(n_45),
.B1(n_2),
.B2(n_3),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_65),
.B(n_12),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_144),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_65),
.B(n_10),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_77),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_84),
.A2(n_52),
.B1(n_83),
.B2(n_82),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_99),
.Y(n_154)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_94),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_155),
.B(n_173),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_121),
.A2(n_148),
.B1(n_107),
.B2(n_138),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_156),
.A2(n_171),
.B1(n_186),
.B2(n_137),
.Y(n_220)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_113),
.Y(n_159)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_159),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_161),
.A2(n_185),
.B1(n_120),
.B2(n_103),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_115),
.B(n_86),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_162),
.Y(n_203)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_164),
.Y(n_199)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_108),
.Y(n_166)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_108),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_167),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_104),
.Y(n_168)
);

NAND3xp33_ASAP7_75t_L g229 ( 
.A(n_168),
.B(n_184),
.C(n_114),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_105),
.B(n_96),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_169),
.B(n_170),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_134),
.B(n_73),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_148),
.A2(n_107),
.B1(n_133),
.B2(n_149),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_98),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_174),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_111),
.B(n_1),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_122),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_175),
.Y(n_223)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_180),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_97),
.A2(n_81),
.B(n_53),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_177),
.A2(n_103),
.B(n_112),
.Y(n_221)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_122),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_178),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_181),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_183),
.Y(n_207)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_104),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_118),
.A2(n_69),
.B1(n_61),
.B2(n_8),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_2),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_187),
.B(n_188),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_119),
.B(n_4),
.Y(n_188)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_132),
.A2(n_5),
.B(n_6),
.C(n_131),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_189),
.B(n_198),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_101),
.B(n_5),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_191),
.Y(n_217)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_129),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_135),
.B(n_6),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_142),
.Y(n_224)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_143),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_194),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_135),
.B(n_117),
.Y(n_194)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_196),
.Y(n_225)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_98),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_151),
.B(n_127),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_142),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_150),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_232),
.C(n_189),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_206),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_155),
.A2(n_116),
.B1(n_145),
.B2(n_125),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_209),
.A2(n_213),
.B1(n_215),
.B2(n_220),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_182),
.A2(n_179),
.B(n_153),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_210),
.A2(n_168),
.B(n_164),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_L g213 ( 
.A1(n_160),
.A2(n_145),
.B1(n_137),
.B2(n_151),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_153),
.A2(n_127),
.B1(n_150),
.B2(n_143),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_229),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_221),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_224),
.B(n_158),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_173),
.A2(n_112),
.B1(n_123),
.B2(n_114),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_228),
.A2(n_196),
.B1(n_172),
.B2(n_159),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_191),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_165),
.B(n_123),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_157),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_156),
.B(n_124),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_214),
.A2(n_177),
.B1(n_179),
.B2(n_192),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_233),
.A2(n_249),
.B1(n_228),
.B2(n_232),
.Y(n_269)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_235),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_240),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_205),
.A2(n_171),
.B1(n_174),
.B2(n_183),
.Y(n_238)
);

BUFx24_ASAP7_75t_L g276 ( 
.A(n_238),
.Y(n_276)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_154),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_241),
.B(n_246),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_248),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_184),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_243),
.B(n_244),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_200),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_225),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_250),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_201),
.B(n_186),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_214),
.A2(n_181),
.B1(n_178),
.B2(n_166),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_224),
.B(n_193),
.Y(n_250)
);

XNOR2x1_ASAP7_75t_SL g275 ( 
.A(n_251),
.B(n_258),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_202),
.B(n_163),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_255),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_254),
.A2(n_205),
.B1(n_220),
.B2(n_204),
.Y(n_261)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_256),
.Y(n_264)
);

NOR2x1_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_195),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_124),
.C(n_176),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_210),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_237),
.A2(n_252),
.B1(n_257),
.B2(n_245),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_260),
.A2(n_267),
.B1(n_273),
.B2(n_280),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_261),
.A2(n_269),
.B1(n_272),
.B2(n_279),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_237),
.A2(n_221),
.B1(n_206),
.B2(n_216),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_258),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_233),
.A2(n_217),
.B1(n_209),
.B2(n_229),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_252),
.A2(n_217),
.B1(n_210),
.B2(n_207),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_218),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_278),
.C(n_259),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_218),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_245),
.A2(n_226),
.B1(n_207),
.B2(n_227),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_248),
.A2(n_215),
.B1(n_226),
.B2(n_227),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_255),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_235),
.Y(n_300)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_285),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_244),
.Y(n_287)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_287),
.Y(n_313)
);

BUFx12f_ASAP7_75t_SL g288 ( 
.A(n_275),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_288),
.Y(n_315)
);

INVx13_ASAP7_75t_L g289 ( 
.A(n_268),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_289),
.Y(n_310)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_268),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_291),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_270),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_263),
.B(n_274),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_299),
.Y(n_308)
);

NOR4xp25_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_236),
.C(n_257),
.D(n_251),
.Y(n_293)
);

OAI322xp33_ASAP7_75t_L g314 ( 
.A1(n_293),
.A2(n_250),
.A3(n_230),
.B1(n_239),
.B2(n_241),
.C1(n_276),
.C2(n_200),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_267),
.A2(n_260),
.B1(n_273),
.B2(n_277),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_294),
.A2(n_296),
.B1(n_303),
.B2(n_304),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_265),
.C(n_247),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_234),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_281),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_297),
.B(n_298),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_283),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_275),
.A2(n_258),
.B(n_256),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_300),
.B(n_301),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_266),
.B(n_246),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_249),
.Y(n_316)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_283),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_271),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_294),
.A2(n_269),
.B1(n_272),
.B2(n_280),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_307),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_284),
.A2(n_265),
.B1(n_278),
.B2(n_263),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_311),
.B(n_319),
.Y(n_336)
);

A2O1A1O1Ixp25_ASAP7_75t_L g323 ( 
.A1(n_314),
.A2(n_293),
.B(n_299),
.C(n_287),
.D(n_296),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_320),
.C(n_291),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_286),
.A2(n_276),
.B1(n_254),
.B2(n_223),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_321),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_204),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_219),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_286),
.A2(n_276),
.B1(n_223),
.B2(n_211),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_307),
.Y(n_337)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_313),
.Y(n_324)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_324),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_326),
.B(n_329),
.C(n_330),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_306),
.A2(n_313),
.B(n_315),
.Y(n_328)
);

OAI21x1_ASAP7_75t_SL g343 ( 
.A1(n_328),
.A2(n_333),
.B(n_334),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_295),
.C(n_303),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_304),
.C(n_290),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_285),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_330),
.Y(n_344)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_322),
.Y(n_332)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_332),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_305),
.A2(n_288),
.B(n_297),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_321),
.A2(n_289),
.B(n_211),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_309),
.Y(n_335)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_335),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_337),
.A2(n_344),
.B(n_329),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_333),
.A2(n_318),
.B1(n_312),
.B2(n_310),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_339),
.B(n_347),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_328),
.A2(n_310),
.B1(n_309),
.B2(n_316),
.Y(n_341)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_341),
.Y(n_349)
);

BUFx24_ASAP7_75t_SL g346 ( 
.A(n_323),
.Y(n_346)
);

INVx5_ASAP7_75t_L g354 ( 
.A(n_346),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_326),
.B(n_308),
.C(n_311),
.Y(n_347)
);

NAND2xp33_ASAP7_75t_L g348 ( 
.A(n_339),
.B(n_327),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_348),
.B(n_352),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_342),
.B(n_336),
.Y(n_351)
);

MAJx2_ASAP7_75t_L g356 ( 
.A(n_351),
.B(n_347),
.C(n_308),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_337),
.A2(n_325),
.B(n_334),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_342),
.B(n_336),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_353),
.B(n_327),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_355),
.A2(n_325),
.B1(n_340),
.B2(n_338),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_356),
.B(n_360),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_358),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_345),
.Y(n_359)
);

A2O1A1Ixp33_ASAP7_75t_SL g363 ( 
.A1(n_359),
.A2(n_343),
.B(n_353),
.C(n_351),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_350),
.B(n_354),
.Y(n_361)
);

AO21x1_ASAP7_75t_L g367 ( 
.A1(n_361),
.A2(n_362),
.B(n_354),
.Y(n_367)
);

CKINVDCx14_ASAP7_75t_R g362 ( 
.A(n_350),
.Y(n_362)
);

AOI322xp5_ASAP7_75t_L g369 ( 
.A1(n_363),
.A2(n_222),
.A3(n_167),
.B1(n_175),
.B2(n_212),
.C1(n_141),
.C2(n_219),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_357),
.A2(n_359),
.B(n_362),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_364),
.B(n_367),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_369),
.A2(n_212),
.B(n_222),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_365),
.B(n_366),
.C(n_363),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_370),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_371),
.B(n_368),
.C(n_222),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_373),
.A2(n_372),
.B(n_141),
.Y(n_374)
);

BUFx24_ASAP7_75t_SL g375 ( 
.A(n_374),
.Y(n_375)
);


endmodule