module real_aes_9222_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_753;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g116 ( .A(n_0), .Y(n_116) );
INVx1_ASAP7_75t_L g509 ( .A(n_1), .Y(n_509) );
INVx1_ASAP7_75t_L g269 ( .A(n_2), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_3), .A2(n_39), .B1(n_188), .B2(n_537), .Y(n_536) );
AOI21xp33_ASAP7_75t_L g176 ( .A1(n_4), .A2(n_177), .B(n_178), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_5), .B(n_175), .Y(n_486) );
AND2x6_ASAP7_75t_L g150 ( .A(n_6), .B(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_7), .A2(n_245), .B(n_246), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_8), .B(n_40), .Y(n_117) );
INVx1_ASAP7_75t_L g185 ( .A(n_9), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_10), .B(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g147 ( .A(n_11), .Y(n_147) );
INVx1_ASAP7_75t_L g505 ( .A(n_12), .Y(n_505) );
INVx1_ASAP7_75t_L g251 ( .A(n_13), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_14), .B(n_153), .Y(n_543) );
AOI222xp33_ASAP7_75t_SL g454 ( .A1(n_15), .A2(n_112), .B1(n_455), .B2(n_456), .C1(n_465), .C2(n_752), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_16), .B(n_143), .Y(n_514) );
XNOR2xp5_ASAP7_75t_L g125 ( .A(n_17), .B(n_126), .Y(n_125) );
AO32x2_ASAP7_75t_L g534 ( .A1(n_17), .A2(n_142), .A3(n_175), .B1(n_497), .B2(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_18), .B(n_188), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_19), .B(n_196), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_20), .B(n_143), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_21), .A2(n_51), .B1(n_188), .B2(n_537), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_22), .B(n_177), .Y(n_205) );
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_23), .A2(n_78), .B1(n_153), .B2(n_188), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_24), .B(n_188), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_25), .B(n_173), .Y(n_199) );
OAI22xp5_ASAP7_75t_SL g456 ( .A1(n_26), .A2(n_457), .B1(n_458), .B2(n_464), .Y(n_456) );
INVx1_ASAP7_75t_L g464 ( .A(n_26), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_27), .A2(n_249), .B(n_250), .C(n_252), .Y(n_248) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_28), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_29), .B(n_190), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_30), .B(n_183), .Y(n_270) );
INVx1_ASAP7_75t_L g161 ( .A(n_31), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_32), .B(n_190), .Y(n_531) );
INVx2_ASAP7_75t_L g155 ( .A(n_33), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_34), .B(n_188), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_35), .B(n_190), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_36), .A2(n_105), .B1(n_118), .B2(n_756), .Y(n_104) );
AOI22xp5_ASAP7_75t_L g130 ( .A1(n_37), .A2(n_43), .B1(n_131), .B2(n_132), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_37), .Y(n_132) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_38), .A2(n_150), .B(n_162), .C(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g159 ( .A(n_41), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_42), .B(n_183), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_43), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_44), .B(n_188), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_45), .A2(n_88), .B1(n_213), .B2(n_537), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_46), .B(n_188), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_47), .B(n_188), .Y(n_506) );
CKINVDCx16_ASAP7_75t_R g165 ( .A(n_48), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_49), .B(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_50), .B(n_177), .Y(n_239) );
AOI22xp33_ASAP7_75t_SL g518 ( .A1(n_52), .A2(n_61), .B1(n_153), .B2(n_188), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g152 ( .A1(n_53), .A2(n_153), .B1(n_156), .B2(n_162), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_54), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_55), .B(n_188), .Y(n_496) );
CKINVDCx16_ASAP7_75t_R g266 ( .A(n_56), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_57), .B(n_188), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_58), .A2(n_182), .B(n_184), .C(n_187), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_59), .Y(n_226) );
INVx1_ASAP7_75t_L g179 ( .A(n_60), .Y(n_179) );
INVx1_ASAP7_75t_L g151 ( .A(n_62), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_63), .B(n_188), .Y(n_510) );
INVx1_ASAP7_75t_L g146 ( .A(n_64), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_65), .Y(n_123) );
AO32x2_ASAP7_75t_L g554 ( .A1(n_66), .A2(n_175), .A3(n_231), .B1(n_497), .B2(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g494 ( .A(n_67), .Y(n_494) );
OAI22xp5_ASAP7_75t_SL g128 ( .A1(n_68), .A2(n_129), .B1(n_130), .B2(n_133), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_68), .Y(n_133) );
INVx1_ASAP7_75t_L g526 ( .A(n_69), .Y(n_526) );
A2O1A1Ixp33_ASAP7_75t_SL g195 ( .A1(n_70), .A2(n_187), .B(n_196), .C(n_197), .Y(n_195) );
INVxp67_ASAP7_75t_L g198 ( .A(n_71), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_72), .B(n_153), .Y(n_527) );
INVx1_ASAP7_75t_L g110 ( .A(n_73), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_74), .Y(n_170) );
INVx1_ASAP7_75t_L g219 ( .A(n_75), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_76), .A2(n_102), .B1(n_462), .B2(n_463), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_76), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_77), .B(n_452), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_79), .A2(n_150), .B(n_162), .C(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_80), .B(n_537), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_81), .B(n_153), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_82), .B(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g144 ( .A(n_83), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_84), .B(n_196), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_85), .B(n_153), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_86), .A2(n_150), .B(n_162), .C(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g113 ( .A(n_87), .Y(n_113) );
OR2x2_ASAP7_75t_L g450 ( .A(n_87), .B(n_114), .Y(n_450) );
OR2x2_ASAP7_75t_L g468 ( .A(n_87), .B(n_115), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_89), .A2(n_103), .B1(n_153), .B2(n_154), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_90), .B(n_190), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g273 ( .A(n_91), .Y(n_273) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_92), .A2(n_150), .B(n_162), .C(n_234), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_93), .Y(n_241) );
INVx1_ASAP7_75t_L g194 ( .A(n_94), .Y(n_194) );
CKINVDCx16_ASAP7_75t_R g247 ( .A(n_95), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_96), .B(n_209), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_97), .A2(n_459), .B1(n_460), .B2(n_461), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_97), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_98), .B(n_153), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_99), .B(n_175), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_100), .B(n_110), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_101), .A2(n_177), .B(n_193), .Y(n_192) );
CKINVDCx16_ASAP7_75t_R g463 ( .A(n_102), .Y(n_463) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx12_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_108), .Y(n_756) );
OR2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
INVx3_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
NOR2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OR2x2_ASAP7_75t_L g751 ( .A(n_113), .B(n_115), .Y(n_751) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
OA21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_124), .B(n_453), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g755 ( .A(n_123), .Y(n_755) );
OAI21x1_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_447), .B(n_451), .Y(n_124) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_128), .B1(n_134), .B2(n_135), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_128), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_130), .Y(n_129) );
OAI22xp5_ASAP7_75t_SL g465 ( .A1(n_134), .A2(n_466), .B1(n_469), .B2(n_749), .Y(n_465) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OAI22xp5_ASAP7_75t_SL g752 ( .A1(n_135), .A2(n_466), .B1(n_753), .B2(n_754), .Y(n_752) );
AND3x1_ASAP7_75t_L g135 ( .A(n_136), .B(n_372), .C(n_421), .Y(n_135) );
NOR3xp33_ASAP7_75t_SL g136 ( .A(n_137), .B(n_279), .C(n_317), .Y(n_136) );
OAI222xp33_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_200), .B1(n_254), .B2(n_260), .C1(n_274), .C2(n_277), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_171), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_139), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_139), .B(n_322), .Y(n_413) );
BUFx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OR2x2_ASAP7_75t_L g290 ( .A(n_140), .B(n_191), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_140), .B(n_172), .Y(n_298) );
AND2x2_ASAP7_75t_L g333 ( .A(n_140), .B(n_310), .Y(n_333) );
OR2x2_ASAP7_75t_L g357 ( .A(n_140), .B(n_172), .Y(n_357) );
OR2x2_ASAP7_75t_L g365 ( .A(n_140), .B(n_264), .Y(n_365) );
AND2x2_ASAP7_75t_L g368 ( .A(n_140), .B(n_191), .Y(n_368) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
OR2x2_ASAP7_75t_L g262 ( .A(n_141), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g276 ( .A(n_141), .B(n_191), .Y(n_276) );
AND2x2_ASAP7_75t_L g326 ( .A(n_141), .B(n_264), .Y(n_326) );
AND2x2_ASAP7_75t_L g339 ( .A(n_141), .B(n_172), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_141), .B(n_425), .Y(n_446) );
AO21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_148), .B(n_169), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_142), .B(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g214 ( .A(n_142), .Y(n_214) );
AO21x2_ASAP7_75t_L g264 ( .A1(n_142), .A2(n_265), .B(n_272), .Y(n_264) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_143), .Y(n_175) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
AND2x2_ASAP7_75t_SL g190 ( .A(n_144), .B(n_145), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
OAI22xp33_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_152), .B1(n_165), .B2(n_166), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_L g178 ( .A1(n_149), .A2(n_179), .B(n_180), .C(n_181), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_149), .A2(n_180), .B(n_194), .C(n_195), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_149), .A2(n_180), .B(n_247), .C(n_248), .Y(n_246) );
INVx4_ASAP7_75t_SL g149 ( .A(n_150), .Y(n_149) );
NAND2x1p5_ASAP7_75t_L g166 ( .A(n_150), .B(n_167), .Y(n_166) );
AND2x4_ASAP7_75t_L g177 ( .A(n_150), .B(n_167), .Y(n_177) );
OAI21xp5_ASAP7_75t_L g477 ( .A1(n_150), .A2(n_478), .B(n_481), .Y(n_477) );
BUFx3_ASAP7_75t_L g497 ( .A(n_150), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g503 ( .A1(n_150), .A2(n_504), .B(n_508), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_150), .A2(n_525), .B(n_528), .Y(n_524) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_150), .A2(n_541), .B(n_545), .Y(n_540) );
INVx2_ASAP7_75t_L g271 ( .A(n_153), .Y(n_271) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g163 ( .A(n_155), .Y(n_163) );
INVx1_ASAP7_75t_L g168 ( .A(n_155), .Y(n_168) );
OAI22xp5_ASAP7_75t_SL g156 ( .A1(n_157), .A2(n_159), .B1(n_160), .B2(n_161), .Y(n_156) );
INVx2_ASAP7_75t_L g160 ( .A(n_157), .Y(n_160) );
INVx4_ASAP7_75t_L g249 ( .A(n_157), .Y(n_249) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g164 ( .A(n_158), .Y(n_164) );
AND2x2_ASAP7_75t_L g167 ( .A(n_158), .B(n_168), .Y(n_167) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_158), .Y(n_183) );
INVx3_ASAP7_75t_L g186 ( .A(n_158), .Y(n_186) );
INVx1_ASAP7_75t_L g196 ( .A(n_158), .Y(n_196) );
INVx5_ASAP7_75t_L g180 ( .A(n_162), .Y(n_180) );
AND2x6_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_163), .Y(n_188) );
BUFx3_ASAP7_75t_L g213 ( .A(n_163), .Y(n_213) );
INVx1_ASAP7_75t_L g537 ( .A(n_163), .Y(n_537) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_166), .A2(n_219), .B(n_220), .Y(n_218) );
OAI21xp5_ASAP7_75t_L g265 ( .A1(n_166), .A2(n_266), .B(n_267), .Y(n_265) );
INVx1_ASAP7_75t_L g484 ( .A(n_168), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_L g364 ( .A1(n_171), .A2(n_365), .B(n_366), .C(n_369), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_171), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_171), .B(n_309), .Y(n_431) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_191), .Y(n_171) );
AND2x2_ASAP7_75t_SL g275 ( .A(n_172), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g289 ( .A(n_172), .Y(n_289) );
AND2x2_ASAP7_75t_L g316 ( .A(n_172), .B(n_310), .Y(n_316) );
INVx1_ASAP7_75t_SL g324 ( .A(n_172), .Y(n_324) );
AND2x2_ASAP7_75t_L g347 ( .A(n_172), .B(n_348), .Y(n_347) );
BUFx2_ASAP7_75t_L g425 ( .A(n_172), .Y(n_425) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_176), .B(n_189), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NOR2xp33_ASAP7_75t_SL g215 ( .A(n_174), .B(n_216), .Y(n_215) );
NAND3xp33_ASAP7_75t_L g515 ( .A(n_174), .B(n_497), .C(n_516), .Y(n_515) );
AO21x1_ASAP7_75t_L g560 ( .A1(n_174), .A2(n_516), .B(n_561), .Y(n_560) );
INVx4_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
OA21x2_ASAP7_75t_L g191 ( .A1(n_175), .A2(n_192), .B(n_199), .Y(n_191) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_175), .A2(n_477), .B(n_486), .Y(n_476) );
BUFx2_ASAP7_75t_L g245 ( .A(n_177), .Y(n_245) );
O2A1O1Ixp5_ASAP7_75t_L g493 ( .A1(n_182), .A2(n_494), .B(n_495), .C(n_496), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_182), .A2(n_546), .B(n_547), .Y(n_545) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx4_ASAP7_75t_L g237 ( .A(n_183), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_183), .A2(n_485), .B1(n_517), .B2(n_518), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_183), .A2(n_485), .B1(n_536), .B2(n_538), .Y(n_535) );
OAI22xp5_ASAP7_75t_SL g555 ( .A1(n_183), .A2(n_186), .B1(n_556), .B2(n_557), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_186), .B(n_198), .Y(n_197) );
INVx5_ASAP7_75t_L g209 ( .A(n_186), .Y(n_209) );
O2A1O1Ixp5_ASAP7_75t_SL g525 ( .A1(n_187), .A2(n_209), .B(n_526), .C(n_527), .Y(n_525) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_188), .Y(n_238) );
INVx1_ASAP7_75t_L g227 ( .A(n_190), .Y(n_227) );
INVx2_ASAP7_75t_L g231 ( .A(n_190), .Y(n_231) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_190), .A2(n_244), .B(n_253), .Y(n_243) );
OA21x2_ASAP7_75t_L g523 ( .A1(n_190), .A2(n_524), .B(n_531), .Y(n_523) );
OA21x2_ASAP7_75t_L g539 ( .A1(n_190), .A2(n_540), .B(n_548), .Y(n_539) );
BUFx2_ASAP7_75t_L g261 ( .A(n_191), .Y(n_261) );
INVx1_ASAP7_75t_L g323 ( .A(n_191), .Y(n_323) );
INVx3_ASAP7_75t_L g348 ( .A(n_191), .Y(n_348) );
INVx1_ASAP7_75t_L g544 ( .A(n_196), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_200), .B(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_228), .Y(n_200) );
INVx1_ASAP7_75t_L g344 ( .A(n_201), .Y(n_344) );
OAI32xp33_ASAP7_75t_L g350 ( .A1(n_201), .A2(n_289), .A3(n_351), .B1(n_352), .B2(n_353), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_201), .A2(n_355), .B1(n_358), .B2(n_363), .Y(n_354) );
INVx4_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g292 ( .A(n_202), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g370 ( .A(n_202), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g440 ( .A(n_202), .B(n_386), .Y(n_440) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_217), .Y(n_202) );
AND2x2_ASAP7_75t_L g255 ( .A(n_203), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g285 ( .A(n_203), .Y(n_285) );
INVx1_ASAP7_75t_L g304 ( .A(n_203), .Y(n_304) );
OR2x2_ASAP7_75t_L g312 ( .A(n_203), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g319 ( .A(n_203), .B(n_293), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_203), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g340 ( .A(n_203), .B(n_258), .Y(n_340) );
INVx3_ASAP7_75t_L g362 ( .A(n_203), .Y(n_362) );
AND2x2_ASAP7_75t_L g387 ( .A(n_203), .B(n_259), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_203), .B(n_352), .Y(n_435) );
OR2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_215), .Y(n_203) );
AOI21xp5_ASAP7_75t_SL g204 ( .A1(n_205), .A2(n_206), .B(n_214), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_210), .B(n_211), .Y(n_207) );
O2A1O1Ixp33_ASAP7_75t_L g268 ( .A1(n_209), .A2(n_269), .B(n_270), .C(n_271), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_209), .A2(n_479), .B(n_480), .Y(n_478) );
INVx2_ASAP7_75t_L g485 ( .A(n_209), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_209), .A2(n_491), .B(n_492), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_211), .A2(n_222), .B(n_223), .Y(n_221) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g252 ( .A(n_213), .Y(n_252) );
INVx1_ASAP7_75t_L g224 ( .A(n_214), .Y(n_224) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_214), .A2(n_489), .B(n_498), .Y(n_488) );
OA21x2_ASAP7_75t_L g502 ( .A1(n_214), .A2(n_503), .B(n_511), .Y(n_502) );
INVx2_ASAP7_75t_L g259 ( .A(n_217), .Y(n_259) );
AND2x2_ASAP7_75t_L g391 ( .A(n_217), .B(n_229), .Y(n_391) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_224), .B(n_225), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_227), .B(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_227), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g433 ( .A(n_228), .Y(n_433) );
OR2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_242), .Y(n_228) );
INVx1_ASAP7_75t_L g278 ( .A(n_229), .Y(n_278) );
AND2x2_ASAP7_75t_L g305 ( .A(n_229), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_229), .B(n_259), .Y(n_313) );
AND2x2_ASAP7_75t_L g371 ( .A(n_229), .B(n_294), .Y(n_371) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g257 ( .A(n_230), .Y(n_257) );
AND2x2_ASAP7_75t_L g284 ( .A(n_230), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g293 ( .A(n_230), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_230), .B(n_259), .Y(n_359) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_240), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_239), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_238), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_242), .B(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g306 ( .A(n_242), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_242), .B(n_259), .Y(n_352) );
AND2x2_ASAP7_75t_L g361 ( .A(n_242), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g386 ( .A(n_242), .Y(n_386) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g258 ( .A(n_243), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g294 ( .A(n_243), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_249), .B(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g507 ( .A(n_249), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_249), .A2(n_529), .B(n_530), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_254), .A2(n_264), .B1(n_423), .B2(n_426), .Y(n_422) );
INVx1_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
OAI21xp5_ASAP7_75t_SL g445 ( .A1(n_256), .A2(n_367), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_257), .B(n_362), .Y(n_379) );
INVx1_ASAP7_75t_L g404 ( .A(n_257), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_258), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g331 ( .A(n_258), .B(n_284), .Y(n_331) );
INVx2_ASAP7_75t_L g287 ( .A(n_259), .Y(n_287) );
INVx1_ASAP7_75t_L g337 ( .A(n_259), .Y(n_337) );
OAI221xp5_ASAP7_75t_L g428 ( .A1(n_260), .A2(n_412), .B1(n_429), .B2(n_432), .C(n_434), .Y(n_428) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx1_ASAP7_75t_L g299 ( .A(n_261), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_261), .B(n_310), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_262), .B(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g353 ( .A(n_262), .B(n_299), .Y(n_353) );
INVx3_ASAP7_75t_SL g394 ( .A(n_262), .Y(n_394) );
AND2x2_ASAP7_75t_L g338 ( .A(n_263), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g367 ( .A(n_263), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_263), .B(n_276), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_263), .B(n_322), .Y(n_408) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx3_ASAP7_75t_L g310 ( .A(n_264), .Y(n_310) );
OAI322xp33_ASAP7_75t_L g405 ( .A1(n_264), .A2(n_336), .A3(n_358), .B1(n_406), .B2(n_408), .C1(n_409), .C2(n_410), .Y(n_405) );
O2A1O1Ixp33_ASAP7_75t_L g504 ( .A1(n_271), .A2(n_505), .B(n_506), .C(n_507), .Y(n_504) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AOI21xp33_ASAP7_75t_L g429 ( .A1(n_275), .A2(n_278), .B(n_430), .Y(n_429) );
NOR2xp33_ASAP7_75t_SL g355 ( .A(n_276), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g377 ( .A(n_276), .B(n_289), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_276), .B(n_316), .Y(n_392) );
INVxp67_ASAP7_75t_L g343 ( .A(n_278), .Y(n_343) );
AOI211xp5_ASAP7_75t_L g349 ( .A1(n_278), .A2(n_350), .B(n_354), .C(n_364), .Y(n_349) );
OAI221xp5_ASAP7_75t_SL g279 ( .A1(n_280), .A2(n_288), .B1(n_291), .B2(n_295), .C(n_300), .Y(n_279) );
INVxp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_286), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g303 ( .A(n_287), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g420 ( .A(n_287), .Y(n_420) );
OAI221xp5_ASAP7_75t_L g436 ( .A1(n_288), .A2(n_437), .B1(n_442), .B2(n_443), .C(n_445), .Y(n_436) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_289), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_SL g336 ( .A(n_289), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_289), .B(n_367), .Y(n_374) );
AND2x2_ASAP7_75t_L g416 ( .A(n_289), .B(n_394), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_290), .B(n_315), .Y(n_314) );
OAI22xp33_ASAP7_75t_L g411 ( .A1(n_290), .A2(n_302), .B1(n_412), .B2(n_413), .Y(n_411) );
OR2x2_ASAP7_75t_L g442 ( .A(n_290), .B(n_310), .Y(n_442) );
CKINVDCx16_ASAP7_75t_R g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g419 ( .A(n_293), .Y(n_419) );
AND2x2_ASAP7_75t_L g444 ( .A(n_293), .B(n_387), .Y(n_444) );
INVxp67_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NOR2xp33_ASAP7_75t_SL g296 ( .A(n_297), .B(n_299), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g308 ( .A(n_298), .B(n_309), .Y(n_308) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_307), .B1(n_311), .B2(n_314), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx1_ASAP7_75t_L g375 ( .A(n_303), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_303), .B(n_343), .Y(n_410) );
AOI322xp5_ASAP7_75t_L g334 ( .A1(n_305), .A2(n_335), .A3(n_337), .B1(n_338), .B2(n_340), .C1(n_341), .C2(n_345), .Y(n_334) );
INVxp67_ASAP7_75t_L g328 ( .A(n_306), .Y(n_328) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_308), .A2(n_313), .B1(n_330), .B2(n_332), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_309), .B(n_322), .Y(n_409) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_310), .B(n_348), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_310), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g406 ( .A(n_312), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
NAND3xp33_ASAP7_75t_SL g317 ( .A(n_318), .B(n_334), .C(n_349), .Y(n_317) );
AOI221xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_320), .B1(n_325), .B2(n_327), .C(n_329), .Y(n_318) );
AND2x2_ASAP7_75t_L g325 ( .A(n_321), .B(n_326), .Y(n_325) );
INVx3_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
AND2x2_ASAP7_75t_L g335 ( .A(n_326), .B(n_336), .Y(n_335) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_328), .Y(n_407) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_333), .B(n_347), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_336), .B(n_394), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_337), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g412 ( .A(n_340), .Y(n_412) );
AND2x2_ASAP7_75t_L g427 ( .A(n_340), .B(n_404), .Y(n_427) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AOI211xp5_ASAP7_75t_L g421 ( .A1(n_351), .A2(n_422), .B(n_428), .C(n_436), .Y(n_421) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g390 ( .A(n_361), .B(n_391), .Y(n_390) );
NAND2x1_ASAP7_75t_SL g432 ( .A(n_362), .B(n_433), .Y(n_432) );
CKINVDCx16_ASAP7_75t_R g402 ( .A(n_365), .Y(n_402) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g397 ( .A(n_371), .Y(n_397) );
AND2x2_ASAP7_75t_L g401 ( .A(n_371), .B(n_387), .Y(n_401) );
NOR5xp2_ASAP7_75t_L g372 ( .A(n_373), .B(n_388), .C(n_405), .D(n_411), .E(n_414), .Y(n_372) );
OAI221xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B1(n_376), .B2(n_378), .C(n_380), .Y(n_373) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_377), .B(n_435), .Y(n_434) );
INVxp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g403 ( .A(n_387), .B(n_404), .Y(n_403) );
OAI221xp5_ASAP7_75t_SL g388 ( .A1(n_389), .A2(n_392), .B1(n_393), .B2(n_395), .C(n_398), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_401), .B1(n_402), .B2(n_403), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g441 ( .A(n_401), .Y(n_441) );
AOI211xp5_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_417), .B(n_419), .C(n_420), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVxp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_441), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
CKINVDCx14_ASAP7_75t_R g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g452 ( .A(n_450), .Y(n_452) );
NAND3xp33_ASAP7_75t_L g453 ( .A(n_451), .B(n_454), .C(n_755), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
CKINVDCx14_ASAP7_75t_R g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g753 ( .A(n_469), .Y(n_753) );
NAND2x1p5_ASAP7_75t_L g469 ( .A(n_470), .B(n_673), .Y(n_469) );
AND2x2_ASAP7_75t_SL g470 ( .A(n_471), .B(n_631), .Y(n_470) );
NOR4xp25_ASAP7_75t_L g471 ( .A(n_472), .B(n_571), .C(n_607), .D(n_621), .Y(n_471) );
OAI221xp5_ASAP7_75t_SL g472 ( .A1(n_473), .A2(n_519), .B1(n_549), .B2(n_558), .C(n_562), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_473), .B(n_706), .Y(n_705) );
OR2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_499), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_487), .Y(n_475) );
AND2x2_ASAP7_75t_L g568 ( .A(n_476), .B(n_488), .Y(n_568) );
INVx3_ASAP7_75t_L g576 ( .A(n_476), .Y(n_576) );
AND2x2_ASAP7_75t_L g630 ( .A(n_476), .B(n_502), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_476), .B(n_501), .Y(n_666) );
AND2x2_ASAP7_75t_L g724 ( .A(n_476), .B(n_586), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B(n_485), .Y(n_481) );
INVx2_ASAP7_75t_L g495 ( .A(n_484), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_485), .A2(n_495), .B(n_509), .C(n_510), .Y(n_508) );
AND2x2_ASAP7_75t_L g559 ( .A(n_487), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g573 ( .A(n_487), .B(n_502), .Y(n_573) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_488), .B(n_502), .Y(n_588) );
AND2x2_ASAP7_75t_L g600 ( .A(n_488), .B(n_576), .Y(n_600) );
OR2x2_ASAP7_75t_L g602 ( .A(n_488), .B(n_560), .Y(n_602) );
AND2x2_ASAP7_75t_L g637 ( .A(n_488), .B(n_560), .Y(n_637) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_488), .Y(n_682) );
INVx1_ASAP7_75t_L g690 ( .A(n_488), .Y(n_690) );
OAI21xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_493), .B(n_497), .Y(n_489) );
OAI221xp5_ASAP7_75t_L g607 ( .A1(n_499), .A2(n_608), .B1(n_612), .B2(n_616), .C(n_617), .Y(n_607) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g567 ( .A(n_500), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_512), .Y(n_500) );
INVx2_ASAP7_75t_L g566 ( .A(n_501), .Y(n_566) );
AND2x2_ASAP7_75t_L g619 ( .A(n_501), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g638 ( .A(n_501), .B(n_576), .Y(n_638) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g701 ( .A(n_502), .B(n_576), .Y(n_701) );
AND2x2_ASAP7_75t_L g623 ( .A(n_512), .B(n_568), .Y(n_623) );
OAI322xp33_ASAP7_75t_L g691 ( .A1(n_512), .A2(n_647), .A3(n_692), .B1(n_694), .B2(n_697), .C1(n_699), .C2(n_703), .Y(n_691) );
INVx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NOR2x1_ASAP7_75t_L g574 ( .A(n_513), .B(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g587 ( .A(n_513), .Y(n_587) );
AND2x2_ASAP7_75t_L g696 ( .A(n_513), .B(n_576), .Y(n_696) );
AND2x2_ASAP7_75t_L g728 ( .A(n_513), .B(n_600), .Y(n_728) );
OR2x2_ASAP7_75t_L g731 ( .A(n_513), .B(n_732), .Y(n_731) );
AND2x4_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g561 ( .A(n_514), .Y(n_561) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_532), .Y(n_520) );
INVx1_ASAP7_75t_L g744 ( .A(n_521), .Y(n_744) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_L g551 ( .A(n_522), .B(n_539), .Y(n_551) );
INVx2_ASAP7_75t_L g584 ( .A(n_522), .Y(n_584) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g606 ( .A(n_523), .Y(n_606) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_523), .Y(n_614) );
OR2x2_ASAP7_75t_L g738 ( .A(n_523), .B(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g563 ( .A(n_532), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g603 ( .A(n_532), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g655 ( .A(n_532), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_539), .Y(n_532) );
AND2x2_ASAP7_75t_L g552 ( .A(n_533), .B(n_553), .Y(n_552) );
NOR2xp67_ASAP7_75t_L g610 ( .A(n_533), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g664 ( .A(n_533), .B(n_554), .Y(n_664) );
OR2x2_ASAP7_75t_L g672 ( .A(n_533), .B(n_606), .Y(n_672) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx2_ASAP7_75t_L g581 ( .A(n_534), .Y(n_581) );
AND2x2_ASAP7_75t_L g591 ( .A(n_534), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g615 ( .A(n_534), .B(n_539), .Y(n_615) );
AND2x2_ASAP7_75t_L g679 ( .A(n_534), .B(n_554), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_539), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_539), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g592 ( .A(n_539), .Y(n_592) );
INVx1_ASAP7_75t_L g597 ( .A(n_539), .Y(n_597) );
AND2x2_ASAP7_75t_L g609 ( .A(n_539), .B(n_610), .Y(n_609) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_539), .Y(n_687) );
INVx1_ASAP7_75t_L g739 ( .A(n_539), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_543), .B(n_544), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
AND2x2_ASAP7_75t_L g716 ( .A(n_550), .B(n_625), .Y(n_716) );
INVx2_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g643 ( .A(n_552), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g742 ( .A(n_552), .B(n_677), .Y(n_742) );
INVx1_ASAP7_75t_L g564 ( .A(n_553), .Y(n_564) );
AND2x2_ASAP7_75t_L g590 ( .A(n_553), .B(n_584), .Y(n_590) );
BUFx2_ASAP7_75t_L g649 ( .A(n_553), .Y(n_649) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_554), .Y(n_570) );
INVx1_ASAP7_75t_L g580 ( .A(n_554), .Y(n_580) );
NOR2xp67_ASAP7_75t_L g718 ( .A(n_558), .B(n_565), .Y(n_718) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AOI32xp33_ASAP7_75t_L g562 ( .A1(n_559), .A2(n_563), .A3(n_565), .B1(n_567), .B2(n_569), .Y(n_562) );
AND2x2_ASAP7_75t_L g702 ( .A(n_559), .B(n_575), .Y(n_702) );
AND2x2_ASAP7_75t_L g740 ( .A(n_559), .B(n_638), .Y(n_740) );
INVx1_ASAP7_75t_L g620 ( .A(n_560), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_564), .B(n_626), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_565), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_565), .B(n_568), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g719 ( .A(n_565), .B(n_637), .Y(n_719) );
OR2x2_ASAP7_75t_L g733 ( .A(n_565), .B(n_602), .Y(n_733) );
INVx3_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g660 ( .A(n_566), .B(n_568), .Y(n_660) );
OR2x2_ASAP7_75t_L g669 ( .A(n_566), .B(n_656), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_568), .B(n_619), .Y(n_641) );
INVx2_ASAP7_75t_L g656 ( .A(n_570), .Y(n_656) );
OR2x2_ASAP7_75t_L g671 ( .A(n_570), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g686 ( .A(n_570), .B(n_687), .Y(n_686) );
A2O1A1Ixp33_ASAP7_75t_L g743 ( .A1(n_570), .A2(n_663), .B(n_744), .C(n_745), .Y(n_743) );
OAI321xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_577), .A3(n_582), .B1(n_585), .B2(n_589), .C(n_593), .Y(n_571) );
INVx1_ASAP7_75t_L g684 ( .A(n_572), .Y(n_684) );
NAND2x1p5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
AND2x2_ASAP7_75t_L g695 ( .A(n_573), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g647 ( .A(n_575), .Y(n_647) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_576), .B(n_690), .Y(n_707) );
OAI221xp5_ASAP7_75t_L g714 ( .A1(n_577), .A2(n_715), .B1(n_717), .B2(n_719), .C(n_720), .Y(n_714) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
AND2x2_ASAP7_75t_L g652 ( .A(n_579), .B(n_626), .Y(n_652) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_580), .B(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g625 ( .A(n_581), .Y(n_625) );
A2O1A1Ixp33_ASAP7_75t_L g667 ( .A1(n_582), .A2(n_623), .B(n_668), .C(n_670), .Y(n_667) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g634 ( .A(n_584), .B(n_591), .Y(n_634) );
BUFx2_ASAP7_75t_L g644 ( .A(n_584), .Y(n_644) );
INVx1_ASAP7_75t_L g659 ( .A(n_584), .Y(n_659) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
OR2x2_ASAP7_75t_L g665 ( .A(n_587), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g748 ( .A(n_587), .Y(n_748) );
INVx1_ASAP7_75t_L g741 ( .A(n_588), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
AND2x2_ASAP7_75t_L g594 ( .A(n_590), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g698 ( .A(n_590), .B(n_615), .Y(n_698) );
INVx1_ASAP7_75t_L g627 ( .A(n_591), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_598), .B1(n_601), .B2(n_603), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_595), .B(n_711), .Y(n_710) );
INVxp67_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x4_ASAP7_75t_L g663 ( .A(n_596), .B(n_664), .Y(n_663) );
BUFx3_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_SL g626 ( .A(n_597), .B(n_606), .Y(n_626) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g618 ( .A(n_600), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g628 ( .A(n_602), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
OAI221xp5_ASAP7_75t_L g722 ( .A1(n_605), .A2(n_723), .B1(n_725), .B2(n_726), .C(n_727), .Y(n_722) );
INVx1_ASAP7_75t_L g611 ( .A(n_606), .Y(n_611) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_606), .Y(n_677) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_609), .B(n_728), .Y(n_727) );
OAI21xp5_ASAP7_75t_L g617 ( .A1(n_610), .A2(n_615), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_613), .B(n_623), .Y(n_720) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx1_ASAP7_75t_L g689 ( .A(n_614), .Y(n_689) );
AND2x2_ASAP7_75t_L g648 ( .A(n_615), .B(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g737 ( .A(n_615), .Y(n_737) );
INVx1_ASAP7_75t_L g653 ( .A(n_618), .Y(n_653) );
INVx1_ASAP7_75t_L g708 ( .A(n_619), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_624), .B1(n_627), .B2(n_628), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_625), .B(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g693 ( .A(n_626), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g730 ( .A(n_626), .B(n_664), .Y(n_730) );
OR2x2_ASAP7_75t_L g703 ( .A(n_627), .B(n_656), .Y(n_703) );
INVx1_ASAP7_75t_L g642 ( .A(n_628), .Y(n_642) );
INVx1_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_630), .B(n_681), .Y(n_680) );
NOR3xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_650), .C(n_661), .Y(n_631) );
OAI211xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_635), .B(n_639), .C(n_645), .Y(n_632) );
INVxp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_634), .A2(n_705), .B1(n_709), .B2(n_712), .C(n_714), .Y(n_704) );
INVx1_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
AND2x2_ASAP7_75t_L g646 ( .A(n_637), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g700 ( .A(n_637), .B(n_701), .Y(n_700) );
OAI211xp5_ASAP7_75t_L g685 ( .A1(n_638), .A2(n_686), .B(n_688), .C(n_690), .Y(n_685) );
INVx2_ASAP7_75t_L g732 ( .A(n_638), .Y(n_732) );
OAI21xp5_ASAP7_75t_SL g639 ( .A1(n_640), .A2(n_642), .B(n_643), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g711 ( .A(n_644), .B(n_664), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_648), .Y(n_645) );
OAI21xp5_ASAP7_75t_SL g650 ( .A1(n_651), .A2(n_653), .B(n_654), .Y(n_650) );
INVxp67_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OAI21xp5_ASAP7_75t_SL g654 ( .A1(n_655), .A2(n_657), .B(n_660), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_655), .B(n_684), .Y(n_683) );
INVxp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_660), .B(n_747), .Y(n_746) );
OAI21xp33_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_665), .B(n_667), .Y(n_661) );
INVx1_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g688 ( .A(n_664), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AND4x1_ASAP7_75t_L g673 ( .A(n_674), .B(n_704), .C(n_721), .D(n_743), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_675), .B(n_691), .Y(n_674) );
OAI211xp5_ASAP7_75t_SL g675 ( .A1(n_676), .A2(n_680), .B(n_683), .C(n_685), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_679), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_690), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_700), .B(n_702), .Y(n_699) );
INVx1_ASAP7_75t_L g725 ( .A(n_700), .Y(n_725) );
INVx2_ASAP7_75t_SL g713 ( .A(n_701), .Y(n_713) );
OR2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g726 ( .A(n_711), .Y(n_726) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NOR2xp33_ASAP7_75t_SL g721 ( .A(n_722), .B(n_729), .Y(n_721) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
OAI221xp5_ASAP7_75t_SL g729 ( .A1(n_730), .A2(n_731), .B1(n_733), .B2(n_734), .C(n_735), .Y(n_729) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_740), .B1(n_741), .B2(n_742), .Y(n_735) );
NAND2xp5_ASAP7_75t_SL g736 ( .A(n_737), .B(n_738), .Y(n_736) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g754 ( .A(n_750), .Y(n_754) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
endmodule