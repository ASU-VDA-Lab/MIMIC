module fake_jpeg_18567_n_290 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_290);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_8),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g25 ( 
.A(n_23),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_12),
.B(n_10),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_22),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_14),
.Y(n_35)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_27),
.Y(n_55)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_40),
.A2(n_25),
.B1(n_32),
.B2(n_28),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_44),
.A2(n_60),
.B1(n_61),
.B2(n_37),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_35),
.B(n_31),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_31),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_53),
.Y(n_81)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_54),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_17),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_27),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_57),
.B(n_59),
.Y(n_76)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_18),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NAND3xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_17),
.C(n_20),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_57),
.B(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_75),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_48),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_69),
.B(n_70),
.Y(n_83)
);

MAJx2_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_55),
.C(n_31),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_32),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_33),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_44),
.A2(n_42),
.B1(n_43),
.B2(n_37),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_78),
.A2(n_25),
.B1(n_61),
.B2(n_49),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_42),
.B1(n_25),
.B2(n_37),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_39),
.B1(n_58),
.B2(n_53),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_81),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_95),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_84),
.A2(n_89),
.B1(n_24),
.B2(n_68),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_56),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_25),
.B1(n_49),
.B2(n_32),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_50),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_72),
.B1(n_65),
.B2(n_51),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_29),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_56),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_98),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_23),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_96),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_56),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_64),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_64),
.Y(n_104)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_70),
.C(n_73),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_113),
.C(n_96),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_85),
.B(n_76),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_118),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g154 ( 
.A1(n_107),
.A2(n_123),
.B1(n_71),
.B2(n_60),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_98),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_117),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_69),
.Y(n_109)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_90),
.B(n_69),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_96),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_88),
.A2(n_73),
.B1(n_72),
.B2(n_65),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_112),
.A2(n_84),
.B1(n_89),
.B2(n_96),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_66),
.C(n_24),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_56),
.Y(n_114)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_92),
.B1(n_99),
.B2(n_47),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_68),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_120),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_83),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_121),
.Y(n_126)
);

AO22x1_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_60),
.B1(n_51),
.B2(n_29),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_87),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_125),
.A2(n_129),
.B(n_122),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_93),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_140),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_83),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_124),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_131),
.B(n_141),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_88),
.B1(n_97),
.B2(n_100),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_149),
.B1(n_71),
.B2(n_103),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_133),
.B(n_18),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_142),
.C(n_113),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_104),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_139),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_138),
.A2(n_33),
.B1(n_29),
.B2(n_30),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_117),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_120),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_95),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_89),
.C(n_84),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_102),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_148),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_95),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_144),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_145),
.A2(n_116),
.B1(n_107),
.B2(n_122),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_101),
.B(n_99),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_151),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_102),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_112),
.A2(n_71),
.B1(n_17),
.B2(n_11),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_114),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_46),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_77),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_103),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_77),
.Y(n_170)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_174),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_173),
.C(n_127),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_130),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_170),
.Y(n_203)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_163),
.A2(n_138),
.B1(n_150),
.B2(n_139),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_125),
.A2(n_107),
.B(n_123),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_164),
.A2(n_162),
.B(n_155),
.Y(n_185)
);

XOR2x2_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_123),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_165),
.A2(n_179),
.B(n_154),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_107),
.B1(n_11),
.B2(n_18),
.Y(n_166)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_172),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_46),
.C(n_52),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_176),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_126),
.B(n_77),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_177),
.A2(n_180),
.B1(n_11),
.B2(n_19),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_128),
.B(n_52),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_158),
.Y(n_193)
);

NAND3xp33_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_21),
.C(n_20),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_125),
.B(n_46),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_154),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_182),
.A2(n_145),
.B1(n_142),
.B2(n_135),
.Y(n_186)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_186),
.A2(n_205),
.B1(n_168),
.B2(n_156),
.Y(n_207)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_155),
.A2(n_148),
.B1(n_143),
.B2(n_129),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_190),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_198),
.C(n_160),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_129),
.B1(n_146),
.B2(n_154),
.Y(n_190)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_195),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_194),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_140),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_181),
.A2(n_14),
.B1(n_1),
.B2(n_2),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_200),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_52),
.C(n_33),
.Y(n_198)
);

FAx1_ASAP7_75t_SL g200 ( 
.A(n_165),
.B(n_167),
.CI(n_171),
.CON(n_200),
.SN(n_200)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_52),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_180),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_164),
.A2(n_14),
.B1(n_20),
.B2(n_21),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_201),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_159),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_210),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_159),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_189),
.B(n_171),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_218),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_219),
.C(n_30),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_169),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_175),
.C(n_172),
.Y(n_219)
);

FAx1_ASAP7_75t_SL g220 ( 
.A(n_188),
.B(n_190),
.CI(n_200),
.CON(n_220),
.SN(n_220)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_22),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_177),
.Y(n_222)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_222),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_186),
.A2(n_161),
.B1(n_174),
.B2(n_182),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_192),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_187),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_224),
.B(n_196),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_231),
.Y(n_242)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_229),
.B(n_232),
.Y(n_252)
);

AOI322xp5_ASAP7_75t_SL g230 ( 
.A1(n_216),
.A2(n_205),
.A3(n_184),
.B1(n_200),
.B2(n_199),
.C1(n_183),
.C2(n_192),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_230),
.B(n_10),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_215),
.A2(n_204),
.B1(n_195),
.B2(n_21),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_217),
.B(n_52),
.Y(n_232)
);

NOR2xp67_ASAP7_75t_SL g234 ( 
.A(n_211),
.B(n_22),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_239),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_219),
.C(n_221),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_212),
.A2(n_10),
.B1(n_9),
.B2(n_8),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_237),
.A2(n_230),
.B1(n_233),
.B2(n_16),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_210),
.C(n_208),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_206),
.C(n_218),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_245),
.C(n_250),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_228),
.A2(n_213),
.B1(n_209),
.B2(n_214),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_243),
.A2(n_250),
.B1(n_252),
.B2(n_242),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_244),
.B(n_248),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_224),
.C(n_220),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_246),
.A2(n_12),
.B1(n_19),
.B2(n_16),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_247),
.A2(n_12),
.B1(n_8),
.B2(n_10),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_30),
.C(n_26),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_30),
.C(n_26),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_26),
.C(n_13),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_225),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_255),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_226),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_257),
.C(n_259),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_14),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_261),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_241),
.A2(n_19),
.B(n_16),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_262),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_249),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_7),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_241),
.A2(n_26),
.B1(n_15),
.B2(n_7),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_246),
.A2(n_22),
.B(n_6),
.Y(n_262)
);

OAI321xp33_ASAP7_75t_L g267 ( 
.A1(n_260),
.A2(n_15),
.A3(n_6),
.B1(n_9),
.B2(n_8),
.C(n_7),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_267),
.A2(n_266),
.B(n_1),
.Y(n_279)
);

AOI31xp67_ASAP7_75t_L g268 ( 
.A1(n_255),
.A2(n_7),
.A3(n_6),
.B(n_15),
.Y(n_268)
);

AOI322xp5_ASAP7_75t_L g280 ( 
.A1(n_268),
.A2(n_271),
.A3(n_274),
.B1(n_0),
.B2(n_2),
.C1(n_3),
.C2(n_4),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_270),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_264),
.A2(n_15),
.B1(n_6),
.B2(n_2),
.Y(n_270)
);

AOI31xp33_ASAP7_75t_L g271 ( 
.A1(n_254),
.A2(n_23),
.A3(n_1),
.B(n_2),
.Y(n_271)
);

NOR2x1_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_23),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_264),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_277),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_265),
.B(n_259),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_266),
.Y(n_278)
);

AO21x1_ASAP7_75t_L g281 ( 
.A1(n_278),
.A2(n_280),
.B(n_265),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_279),
.A2(n_0),
.B(n_3),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_283),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_282),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_284),
.A2(n_275),
.B(n_276),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_285),
.C(n_4),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_5),
.C(n_3),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_5),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_5),
.B(n_3),
.Y(n_290)
);


endmodule