module fake_jpeg_24061_n_333 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_30),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_46),
.B(n_33),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_49),
.Y(n_63)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_20),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_52),
.B(n_67),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_22),
.B1(n_27),
.B2(n_38),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_54),
.A2(n_78),
.B1(n_31),
.B2(n_36),
.Y(n_95)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_74),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_18),
.B(n_32),
.C(n_35),
.Y(n_58)
);

AO22x1_ASAP7_75t_L g118 ( 
.A1(n_58),
.A2(n_28),
.B1(n_25),
.B2(n_21),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_59),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_38),
.B1(n_26),
.B2(n_23),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_61),
.A2(n_65),
.B1(n_75),
.B2(n_76),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_38),
.B1(n_37),
.B2(n_24),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_19),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_69),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_19),
.Y(n_69)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_41),
.A2(n_19),
.B1(n_36),
.B2(n_31),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_41),
.A2(n_37),
.B1(n_24),
.B2(n_35),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_42),
.A2(n_33),
.B1(n_24),
.B2(n_37),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_42),
.A2(n_31),
.B1(n_36),
.B2(n_28),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_79),
.Y(n_120)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_49),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_34),
.Y(n_122)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_57),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_88),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_94),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_95),
.A2(n_119),
.B1(n_122),
.B2(n_34),
.Y(n_149)
);

INVx3_ASAP7_75t_SL g97 ( 
.A(n_60),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_98),
.Y(n_131)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_104),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_70),
.A2(n_49),
.B1(n_51),
.B2(n_47),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_101),
.A2(n_61),
.B1(n_77),
.B2(n_80),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVxp33_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_63),
.B(n_29),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_107),
.B(n_109),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_58),
.B(n_29),
.Y(n_109)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_71),
.B(n_30),
.Y(n_116)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_118),
.B(n_103),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_78),
.B(n_25),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_75),
.B(n_47),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_79),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_124),
.B(n_137),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_126),
.A2(n_147),
.B1(n_104),
.B2(n_99),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_56),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_133),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_121),
.A2(n_62),
.B(n_45),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_129),
.A2(n_134),
.B(n_1),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_53),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_120),
.A2(n_45),
.B(n_55),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_118),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_96),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_139),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_113),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_39),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_157),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_39),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_3),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_89),
.A2(n_80),
.B1(n_34),
.B2(n_20),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_93),
.A2(n_64),
.B1(n_34),
.B2(n_20),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_144),
.A2(n_152),
.B1(n_91),
.B2(n_2),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_123),
.A2(n_93),
.B1(n_98),
.B2(n_101),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_149),
.B(n_9),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_92),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_159),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_123),
.A2(n_17),
.B1(n_30),
.B2(n_3),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_87),
.B(n_17),
.C(n_30),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_1),
.C(n_2),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_17),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_110),
.Y(n_166)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_131),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_160),
.B(n_164),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_163),
.A2(n_184),
.B1(n_186),
.B2(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_170),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_108),
.Y(n_168)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_124),
.A2(n_100),
.B1(n_112),
.B2(n_97),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_169),
.A2(n_173),
.B1(n_144),
.B2(n_143),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_17),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_105),
.Y(n_171)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_110),
.Y(n_172)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_153),
.A2(n_94),
.B1(n_110),
.B2(n_90),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_136),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_174),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_90),
.Y(n_175)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_148),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_176),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_148),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_179),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_178),
.A2(n_190),
.B1(n_126),
.B2(n_146),
.Y(n_198)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_187),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_151),
.C(n_135),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_155),
.B(n_3),
.Y(n_185)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_128),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_129),
.B(n_4),
.Y(n_188)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_192),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_153),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_159),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_134),
.A2(n_9),
.B(n_10),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_157),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_215),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_198),
.A2(n_205),
.B1(n_213),
.B2(n_221),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_140),
.Y(n_200)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_141),
.B1(n_135),
.B2(n_142),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_208),
.A2(n_222),
.B1(n_178),
.B2(n_189),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_184),
.A2(n_141),
.B1(n_145),
.B2(n_154),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_125),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_214),
.B(n_216),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_156),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_219),
.B(n_223),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_171),
.C(n_170),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_161),
.A2(n_142),
.B1(n_146),
.B2(n_130),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_163),
.A2(n_154),
.B1(n_145),
.B2(n_11),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_173),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_201),
.A2(n_188),
.B1(n_165),
.B2(n_169),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_228),
.A2(n_234),
.B1(n_236),
.B2(n_240),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_209),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_239),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_237),
.C(n_243),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_232),
.A2(n_224),
.B1(n_220),
.B2(n_186),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_233),
.B(n_235),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_201),
.A2(n_223),
.B1(n_207),
.B2(n_205),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_222),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_207),
.A2(n_198),
.B1(n_206),
.B2(n_204),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_175),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_197),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_208),
.A2(n_161),
.B1(n_180),
.B2(n_182),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_200),
.B(n_180),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_243),
.Y(n_249)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_245),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_172),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_211),
.B(n_185),
.Y(n_244)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_244),
.Y(n_251)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_212),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_199),
.Y(n_247)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_247),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_199),
.B(n_180),
.C(n_166),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_218),
.C(n_196),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_250),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_233),
.A2(n_194),
.B(n_224),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_200),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_252),
.B(n_266),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_227),
.A2(n_204),
.B(n_206),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_259),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_258),
.A2(n_264),
.B1(n_225),
.B2(n_227),
.Y(n_272)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_231),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_260),
.B(n_265),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_248),
.C(n_241),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_232),
.A2(n_174),
.B1(n_164),
.B2(n_203),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_226),
.B(n_183),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_234),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_229),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_186),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_193),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_230),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_274),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_250),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_254),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_273),
.B(n_277),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_255),
.A2(n_228),
.B1(n_240),
.B2(n_239),
.Y(n_275)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_276),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_251),
.B(n_238),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_259),
.A2(n_238),
.B1(n_176),
.B2(n_190),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_279),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_263),
.Y(n_281)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_281),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g282 ( 
.A(n_255),
.B(n_9),
.CI(n_10),
.CON(n_282),
.SN(n_282)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_282),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_261),
.A2(n_193),
.B1(n_12),
.B2(n_14),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_283),
.Y(n_297)
);

INVxp67_ASAP7_75t_SL g284 ( 
.A(n_256),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_284),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_286),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_252),
.B(n_10),
.Y(n_286)
);

BUFx12_ASAP7_75t_L g291 ( 
.A(n_284),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_291),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_270),
.A2(n_263),
.B(n_262),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_293),
.A2(n_296),
.B(n_280),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_295),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_SL g296 ( 
.A1(n_281),
.A2(n_279),
.B(n_282),
.C(n_257),
.Y(n_296)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_303),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_296),
.Y(n_304)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_304),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_300),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_306),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_289),
.A2(n_274),
.B(n_253),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_290),
.B(n_269),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_307),
.B(n_278),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_296),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_308),
.A2(n_310),
.B1(n_298),
.B2(n_299),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_289),
.A2(n_269),
.B(n_285),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_309),
.A2(n_297),
.B(n_278),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_294),
.B(n_249),
.Y(n_310)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_311),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_315),
.C(n_317),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_302),
.A2(n_288),
.B1(n_292),
.B2(n_297),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_268),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_287),
.C(n_288),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_316),
.A2(n_302),
.B(n_291),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_321),
.A2(n_315),
.B(n_312),
.Y(n_325)
);

AND2x2_ASAP7_75t_SL g322 ( 
.A(n_317),
.B(n_286),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_323),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_318),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_324),
.B(n_325),
.C(n_320),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_327),
.Y(n_329)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_326),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_313),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_328),
.B(n_266),
.Y(n_331)
);

OAI221xp5_ASAP7_75t_SL g332 ( 
.A1(n_331),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.C(n_16),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_12),
.B(n_16),
.Y(n_333)
);


endmodule