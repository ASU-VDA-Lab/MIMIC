module real_jpeg_32116_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g137 ( 
.A(n_0),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_0),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g267 ( 
.A(n_0),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_0),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_0),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_1),
.B(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_1),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_1),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_1),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_1),
.B(n_306),
.Y(n_305)
);

AND2x2_ASAP7_75t_SL g432 ( 
.A(n_1),
.B(n_433),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_1),
.B(n_459),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_2),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_2),
.B(n_260),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_2),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_2),
.B(n_425),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_2),
.B(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_2),
.B(n_473),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_2),
.B(n_478),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_3),
.B(n_187),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_3),
.Y(n_511)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_4),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_5),
.Y(n_228)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_6),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_6),
.Y(n_159)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_6),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_7),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_7),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_7),
.B(n_48),
.Y(n_47)
);

AND2x4_ASAP7_75t_L g85 ( 
.A(n_7),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_7),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_7),
.B(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_7),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_7),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_8),
.B(n_210),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_8),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_8),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_8),
.B(n_40),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_8),
.B(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_8),
.B(n_455),
.Y(n_454)
);

AND2x2_ASAP7_75t_SL g465 ( 
.A(n_8),
.B(n_325),
.Y(n_465)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_9),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_9),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_9),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_10),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_11),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_11),
.B(n_171),
.Y(n_170)
);

AND2x2_ASAP7_75t_SL g197 ( 
.A(n_11),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_SL g230 ( 
.A(n_11),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_11),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_11),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_11),
.B(n_407),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_11),
.B(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_12),
.Y(n_124)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_12),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_13),
.B(n_65),
.Y(n_64)
);

AND2x6_ASAP7_75t_SL g74 ( 
.A(n_13),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_13),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_13),
.B(n_119),
.Y(n_118)
);

NAND2x1_ASAP7_75t_L g165 ( 
.A(n_13),
.B(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g203 ( 
.A(n_13),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_13),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_13),
.B(n_299),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_14),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_15),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_16),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_16),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_16),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_16),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_16),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_16),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_SL g141 ( 
.A(n_16),
.B(n_142),
.Y(n_141)
);

NAND2x1_ASAP7_75t_L g323 ( 
.A(n_16),
.B(n_265),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_17),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_17),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_17),
.B(n_267),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_17),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_17),
.B(n_325),
.Y(n_324)
);

OAI211xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_188),
.B(n_506),
.C(n_508),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_185),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_20),
.B(n_186),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_182),
.Y(n_20)
);

INVxp33_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_143),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_106),
.B2(n_107),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_24),
.B(n_106),
.Y(n_184)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_25),
.B(n_107),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_79),
.Y(n_25)
);

XNOR2x1_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_53),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_42),
.B1(n_51),
.B2(n_52),
.Y(n_27)
);

INVxp67_ASAP7_75t_SL g51 ( 
.A(n_28),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_R g28 ( 
.A(n_29),
.B(n_34),
.C(n_37),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_29),
.A2(n_34),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_29),
.Y(n_110)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_33),
.Y(n_265)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_34),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_34),
.B(n_165),
.C(n_168),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_34),
.A2(n_111),
.B1(n_168),
.B2(n_334),
.Y(n_333)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_35),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_36),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_36),
.Y(n_243)
);

XOR2x2_ASAP7_75t_L g108 ( 
.A(n_37),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_41),
.Y(n_155)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_42)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_46),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_46),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_46),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_47),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_47),
.A2(n_50),
.B1(n_141),
.B2(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_47),
.A2(n_50),
.B1(n_170),
.B2(n_361),
.Y(n_360)
);

INVx8_ASAP7_75t_L g247 ( 
.A(n_48),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_50),
.B(n_134),
.C(n_141),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_50),
.B(n_164),
.C(n_170),
.Y(n_163)
);

XNOR2x1_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_68),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_59),
.C(n_64),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_R g82 ( 
.A1(n_55),
.A2(n_59),
.B1(n_60),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_97),
.C(n_102),
.Y(n_96)
);

MAJx2_ASAP7_75t_L g223 ( 
.A(n_55),
.B(n_224),
.C(n_230),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_55),
.B(n_224),
.Y(n_236)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_58),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_60),
.B1(n_70),
.B2(n_73),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_59),
.B(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_59),
.B(n_121),
.C(n_271),
.Y(n_302)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_61),
.Y(n_240)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_82),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_74),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_70),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_70),
.A2(n_73),
.B1(n_305),
.B2(n_309),
.Y(n_304)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_73),
.B(n_116),
.C(n_305),
.Y(n_339)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_78),
.Y(n_171)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_78),
.Y(n_273)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.C(n_96),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_81),
.B(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_97),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_84),
.B(n_96),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.C(n_91),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_91),
.B1(n_92),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_88),
.A2(n_116),
.B1(n_304),
.B2(n_310),
.Y(n_303)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_89),
.Y(n_469)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_100),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_101),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_103),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_135),
.C(n_138),
.Y(n_134)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_103),
.B(n_138),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_103),
.B(n_280),
.Y(n_400)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_105),
.Y(n_285)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJx2_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.C(n_133),
.Y(n_107)
);

XNOR2x1_ASAP7_75t_SL g181 ( 
.A(n_108),
.B(n_133),
.Y(n_181)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_113),
.B(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.C(n_130),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_114),
.B(n_117),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.C(n_125),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_125),
.B1(n_126),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_122),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_121),
.A2(n_122),
.B1(n_271),
.B2(n_274),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_124),
.Y(n_404)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_130),
.Y(n_379)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_134),
.B(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_157),
.Y(n_160)
);

XOR2x2_ASAP7_75t_SL g161 ( 
.A(n_135),
.B(n_162),
.Y(n_161)
);

XNOR2x1_ASAP7_75t_L g336 ( 
.A(n_135),
.B(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_135),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_135),
.A2(n_406),
.B1(n_408),
.B2(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_137),
.Y(n_281)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

AOI21x1_ASAP7_75t_L g182 ( 
.A1(n_143),
.A2(n_183),
.B(n_184),
.Y(n_182)
);

MAJx2_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_176),
.C(n_179),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_145),
.B(n_503),
.Y(n_502)
);

MAJx2_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_163),
.C(n_172),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_146),
.B(n_382),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_152),
.C(n_161),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_148),
.B(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_149),
.Y(n_151)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_152),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_156),
.B(n_160),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_153),
.A2(n_154),
.B1(n_157),
.B2(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_157),
.B(n_217),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_157),
.Y(n_249)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_157),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_158),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_159),
.Y(n_434)
);

INVx6_ASAP7_75t_L g457 ( 
.A(n_159),
.Y(n_457)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_160),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_160),
.A2(n_254),
.B1(n_410),
.B2(n_411),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_161),
.B(n_369),
.Y(n_368)
);

XNOR2x1_ASAP7_75t_L g382 ( 
.A(n_163),
.B(n_173),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_164),
.B(n_360),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_165),
.B(n_333),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_167),
.Y(n_232)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_168),
.Y(n_334)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_169),
.Y(n_261)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_170),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVxp67_ASAP7_75t_SL g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_177),
.B(n_180),
.Y(n_503)
);

INVxp67_ASAP7_75t_SL g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_185),
.B(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_188),
.B(n_507),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_497),
.B(n_504),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_389),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_343),
.B1(n_383),
.B2(n_388),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_311),
.B(n_340),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_275),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_193),
.B(n_275),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_234),
.C(n_251),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_194),
.B(n_252),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_214),
.B2(n_233),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_195),
.B(n_215),
.C(n_223),
.Y(n_289)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_201),
.Y(n_196)
);

MAJx2_ASAP7_75t_L g287 ( 
.A(n_197),
.B(n_203),
.C(n_208),
.Y(n_287)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_208),
.B2(n_209),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_222),
.B2(n_223),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_217),
.A2(n_218),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_221),
.Y(n_436)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_229),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_229),
.B(n_429),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_230),
.B(n_236),
.Y(n_235)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_234),
.B(n_395),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.C(n_248),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_235),
.B(n_398),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_237),
.B(n_248),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.C(n_244),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_238),
.B(n_444),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_242),
.B(n_245),
.Y(n_444)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_243),
.Y(n_426)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_249),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_262),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_263),
.C(n_269),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.C(n_258),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_255),
.A2(n_256),
.B1(n_258),
.B2(n_259),
.Y(n_410)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_269),
.Y(n_262)
);

OA21x2_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_266),
.B(n_268),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_266),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_287),
.Y(n_286)
);

MAJx2_ASAP7_75t_L g319 ( 
.A(n_268),
.B(n_279),
.C(n_287),
.Y(n_319)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_271),
.Y(n_274)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_288),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJx2_ASAP7_75t_L g312 ( 
.A(n_277),
.B(n_278),
.C(n_288),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_286),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g327 ( 
.A(n_280),
.B(n_283),
.C(n_284),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_291),
.C(n_303),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_303),
.Y(n_290)
);

XNOR2x2_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_301),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_298),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_293),
.B(n_298),
.C(n_329),
.Y(n_328)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_302),
.Y(n_329)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_304),
.Y(n_310)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_305),
.Y(n_309)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

AOI21x1_ASAP7_75t_L g340 ( 
.A1(n_312),
.A2(n_341),
.B(n_342),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_316),
.B2(n_317),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_314),
.B(n_316),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_314),
.B(n_346),
.C(n_347),
.Y(n_345)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_315),
.B(n_317),
.Y(n_341)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_330),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_318),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_321),
.C(n_352),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_328),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_327),
.Y(n_321)
);

XNOR2x1_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_323),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_324),
.Y(n_363)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

MAJx2_ASAP7_75t_L g362 ( 
.A(n_327),
.B(n_363),
.C(n_364),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_328),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_330),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_335),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_336),
.C(n_339),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_339),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_340),
.B(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_372),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_349),
.Y(n_344)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_345),
.Y(n_386)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_349),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_353),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_351),
.B(n_354),
.C(n_367),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_367),
.B1(n_368),
.B2(n_371),
.Y(n_353)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_354),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_356),
.B1(n_357),
.B2(n_358),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_355),
.B(n_362),
.C(n_366),
.Y(n_376)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_362),
.B1(n_365),
.B2(n_366),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_359),
.Y(n_366)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_362),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_372),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_373),
.Y(n_385)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_374),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_377),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_376),
.B(n_500),
.C(n_501),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_378),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_381),
.Y(n_500)
);

NAND3xp33_ASAP7_75t_L g389 ( 
.A(n_383),
.B(n_390),
.C(n_392),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_384),
.A2(n_385),
.B1(n_386),
.B2(n_387),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_393),
.A2(n_412),
.B(n_496),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_396),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_394),
.B(n_396),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_399),
.C(n_409),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_397),
.B(n_494),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_399),
.B(n_409),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_401),
.C(n_405),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_400),
.A2(n_401),
.B1(n_402),
.B2(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_400),
.Y(n_449)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_404),
.Y(n_430)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_404),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_405),
.B(n_448),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_408),
.Y(n_405)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_406),
.Y(n_439)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_410),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_490),
.B(n_495),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_414),
.A2(n_450),
.B(n_489),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_440),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_415),
.B(n_440),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_431),
.C(n_437),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_416),
.A2(n_417),
.B1(n_485),
.B2(n_487),
.Y(n_484)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_428),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_419),
.A2(n_420),
.B1(n_424),
.B2(n_427),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_419),
.B(n_427),
.C(n_428),
.Y(n_442)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_424),
.Y(n_427)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_431),
.A2(n_437),
.B1(n_438),
.B2(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_431),
.Y(n_486)
);

NAND2x1_ASAP7_75t_SL g431 ( 
.A(n_432),
.B(n_435),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_432),
.B(n_435),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_447),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_442),
.A2(n_443),
.B1(n_445),
.B2(n_446),
.Y(n_441)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_442),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_443),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_443),
.B(n_445),
.C(n_492),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_447),
.Y(n_492)
);

AOI21x1_ASAP7_75t_SL g450 ( 
.A1(n_451),
.A2(n_482),
.B(n_488),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_452),
.A2(n_470),
.B(n_481),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_461),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_453),
.B(n_461),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_458),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_454),
.B(n_458),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_454),
.B(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

BUFx4f_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_463),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_462),
.B(n_465),
.C(n_466),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_464),
.A2(n_465),
.B1(n_466),
.B2(n_467),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_471),
.A2(n_476),
.B(n_480),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_475),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_472),
.B(n_475),
.Y(n_480)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_484),
.Y(n_482)
);

NOR2xp67_ASAP7_75t_SL g488 ( 
.A(n_483),
.B(n_484),
.Y(n_488)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_485),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_493),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_491),
.B(n_493),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_502),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_499),
.B(n_502),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_510),
.Y(n_509)
);

INVx5_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);


endmodule