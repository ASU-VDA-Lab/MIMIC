module fake_jpeg_8046_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_28),
.B1(n_31),
.B2(n_25),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_56),
.B1(n_60),
.B2(n_67),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_20),
.C(n_17),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_17),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_31),
.B1(n_28),
.B2(n_23),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_28),
.B1(n_31),
.B2(n_48),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_46),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_38),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_64),
.B(n_47),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_23),
.B1(n_25),
.B2(n_29),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_66),
.A2(n_36),
.B1(n_43),
.B2(n_32),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_23),
.B1(n_25),
.B2(n_29),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_68),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_42),
.A2(n_16),
.B1(n_18),
.B2(n_22),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_70),
.A2(n_33),
.B1(n_35),
.B2(n_34),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_76),
.Y(n_115)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_79),
.Y(n_127)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_69),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_81),
.B(n_88),
.Y(n_136)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_83),
.A2(n_34),
.B1(n_35),
.B2(n_19),
.Y(n_126)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_73),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_84),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_85),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_41),
.B(n_43),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_87),
.A2(n_91),
.B(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_69),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_90),
.B(n_95),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_20),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

AOI21xp33_ASAP7_75t_L g93 ( 
.A1(n_70),
.A2(n_18),
.B(n_16),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_93),
.A2(n_105),
.B(n_106),
.Y(n_131)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_62),
.B(n_40),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_96),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_97),
.A2(n_102),
.B1(n_103),
.B2(n_114),
.Y(n_119)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_68),
.Y(n_99)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_71),
.A2(n_41),
.B(n_36),
.C(n_32),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_72),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_63),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_58),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_107),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_59),
.B(n_36),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_40),
.C(n_39),
.Y(n_130)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_50),
.B(n_36),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_111),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_112),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_59),
.B1(n_53),
.B2(n_72),
.Y(n_121)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

MAJx2_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_44),
.C(n_39),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_122),
.C(n_130),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_121),
.A2(n_125),
.B1(n_141),
.B2(n_119),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_81),
.A2(n_64),
.B(n_33),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_126),
.A2(n_138),
.B1(n_102),
.B2(n_79),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_95),
.A2(n_86),
.B1(n_88),
.B2(n_74),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_87),
.A2(n_21),
.B(n_24),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_74),
.A2(n_44),
.B1(n_40),
.B2(n_39),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_143),
.A2(n_78),
.B1(n_77),
.B2(n_84),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_155),
.B1(n_164),
.B2(n_167),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_91),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_146),
.B(n_147),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_75),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_127),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_148),
.B(n_151),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_76),
.Y(n_149)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_127),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_153),
.Y(n_190)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_134),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_154),
.A2(n_163),
.B1(n_134),
.B2(n_139),
.Y(n_197)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_144),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_158),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_108),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_157),
.A2(n_173),
.B(n_177),
.Y(n_199)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_159),
.A2(n_170),
.B1(n_175),
.B2(n_176),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_104),
.Y(n_160)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_161),
.B(n_162),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_113),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g164 ( 
.A1(n_119),
.A2(n_84),
.B(n_108),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_136),
.B1(n_143),
.B2(n_118),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_165),
.A2(n_169),
.B1(n_171),
.B2(n_174),
.Y(n_196)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_121),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_104),
.Y(n_168)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_90),
.B1(n_105),
.B2(n_106),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_139),
.A2(n_100),
.B1(n_101),
.B2(n_80),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_122),
.A2(n_103),
.B1(n_114),
.B2(n_101),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_116),
.B(n_104),
.Y(n_172)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_124),
.B(n_15),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_132),
.A2(n_109),
.B1(n_112),
.B2(n_78),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_118),
.A2(n_94),
.B1(n_80),
.B2(n_110),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_140),
.A2(n_98),
.B1(n_110),
.B2(n_89),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_116),
.B(n_40),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_146),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_182),
.C(n_185),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_154),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_184),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_124),
.C(n_135),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_183),
.B(n_188),
.Y(n_232)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_135),
.C(n_140),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_166),
.A2(n_142),
.B1(n_133),
.B2(n_120),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_SL g219 ( 
.A1(n_187),
.A2(n_176),
.B(n_164),
.Y(n_219)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_142),
.C(n_129),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_192),
.C(n_205),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_126),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_194),
.Y(n_212)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_149),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_198),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_197),
.A2(n_128),
.B1(n_123),
.B2(n_111),
.Y(n_233)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_133),
.B(n_129),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_201),
.A2(n_27),
.B(n_24),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_147),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_202),
.B(n_194),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_157),
.B(n_39),
.C(n_44),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_27),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_161),
.C(n_148),
.Y(n_221)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_145),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_159),
.Y(n_218)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_184),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_213),
.B(n_235),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_155),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_216),
.B(n_221),
.C(n_230),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_196),
.A2(n_167),
.B1(n_171),
.B2(n_164),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_217),
.A2(n_223),
.B1(n_224),
.B2(n_187),
.Y(n_245)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_219),
.A2(n_222),
.B1(n_181),
.B2(n_193),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_178),
.A2(n_164),
.B1(n_151),
.B2(n_152),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_L g223 ( 
.A1(n_210),
.A2(n_89),
.B1(n_147),
.B2(n_153),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_196),
.A2(n_158),
.B1(n_156),
.B2(n_137),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_200),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_227),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_137),
.Y(n_226)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_111),
.Y(n_228)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_228),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_203),
.Y(n_229)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_128),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_231),
.B(n_238),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_233),
.A2(n_234),
.B1(n_237),
.B2(n_181),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_198),
.A2(n_34),
.B1(n_123),
.B2(n_30),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_186),
.B(n_14),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_204),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_188),
.A2(n_30),
.B1(n_19),
.B2(n_21),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_207),
.B(n_24),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_224),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_228),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_182),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_254),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_241),
.A2(n_258),
.B1(n_0),
.B2(n_1),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_220),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_252),
.C(n_259),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_245),
.A2(n_248),
.B1(n_251),
.B2(n_232),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_217),
.A2(n_185),
.B1(n_189),
.B2(n_207),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_260),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_250),
.B(n_261),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_218),
.A2(n_192),
.B1(n_208),
.B2(n_195),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_211),
.B(n_205),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_199),
.Y(n_254)
);

AOI22x1_ASAP7_75t_L g258 ( 
.A1(n_222),
.A2(n_201),
.B1(n_199),
.B2(n_180),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_190),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_212),
.B(n_24),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_262),
.A2(n_268),
.B1(n_273),
.B2(n_276),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_258),
.A2(n_256),
.B(n_246),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_252),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_221),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_240),
.Y(n_286)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_266),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_251),
.A2(n_227),
.B1(n_215),
.B2(n_238),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_215),
.C(n_226),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_272),
.C(n_269),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_239),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_271),
.B(n_2),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_248),
.B(n_212),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_272),
.B(n_281),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_245),
.A2(n_225),
.B1(n_223),
.B2(n_214),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_253),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_3),
.Y(n_296)
);

A2O1A1O1Ixp25_ASAP7_75t_L g275 ( 
.A1(n_244),
.A2(n_231),
.B(n_236),
.C(n_24),
.D(n_21),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_13),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_242),
.A2(n_255),
.B1(n_241),
.B2(n_247),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_259),
.B(n_213),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_278),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_244),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_254),
.A2(n_30),
.B1(n_19),
.B2(n_14),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_279),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_273),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_282),
.A2(n_295),
.B1(n_292),
.B2(n_271),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_286),
.C(n_287),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_290),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_257),
.C(n_1),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_SL g288 ( 
.A1(n_280),
.A2(n_14),
.A3(n_13),
.B1(n_11),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_294),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_0),
.C(n_1),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_279),
.C(n_265),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_SL g291 ( 
.A(n_264),
.B(n_13),
.C(n_2),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_291),
.A2(n_3),
.B(n_5),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_293),
.A2(n_274),
.B1(n_275),
.B2(n_268),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_7),
.Y(n_307)
);

XNOR2x1_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_282),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_309),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_297),
.A2(n_262),
.B1(n_276),
.B2(n_267),
.Y(n_300)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_300),
.Y(n_311)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_302),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_305),
.B(n_307),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_308),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_285),
.A2(n_264),
.B1(n_8),
.B2(n_9),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_289),
.A2(n_283),
.B(n_287),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_7),
.C(n_8),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_290),
.C(n_8),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_310),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_304),
.B(n_10),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_318),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_305),
.B(n_10),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_301),
.Y(n_320)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_320),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_314),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_315),
.A2(n_299),
.B1(n_298),
.B2(n_303),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_324),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_315),
.A2(n_303),
.B(n_9),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_7),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_325),
.B(n_326),
.Y(n_327)
);

NAND3xp33_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_9),
.C(n_10),
.Y(n_326)
);

AOI21xp33_ASAP7_75t_L g331 ( 
.A1(n_328),
.A2(n_316),
.B(n_311),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_331),
.B(n_332),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_312),
.C(n_323),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_329),
.B(n_328),
.Y(n_334)
);

NAND2xp33_ASAP7_75t_SL g335 ( 
.A(n_334),
.B(n_327),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_323),
.B(n_9),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_10),
.Y(n_337)
);


endmodule