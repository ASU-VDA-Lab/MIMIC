module fake_jpeg_8479_n_279 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_37),
.Y(n_52)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_40),
.Y(n_64)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_43),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_21),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_35),
.Y(n_69)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_27),
.B1(n_29),
.B2(n_24),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_46),
.A2(n_48),
.B1(n_55),
.B2(n_65),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_45),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_43),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_9),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_35),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_69),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_24),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_57),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_27),
.B1(n_29),
.B2(n_18),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_54),
.A2(n_56),
.B1(n_66),
.B2(n_37),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_29),
.B1(n_26),
.B2(n_32),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_23),
.B1(n_18),
.B2(n_32),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_70),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_0),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_71),
.B(n_19),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_38),
.B(n_26),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_42),
.C(n_36),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_23),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_34),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_26),
.B1(n_18),
.B2(n_34),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_35),
.B1(n_22),
.B2(n_33),
.Y(n_66)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_37),
.A2(n_33),
.B1(n_22),
.B2(n_34),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_72),
.A2(n_76),
.B(n_59),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_73),
.B(n_81),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_36),
.B(n_25),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_78),
.B(n_80),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_46),
.C(n_38),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_20),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_84),
.B(n_90),
.Y(n_132)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_51),
.A2(n_33),
.B1(n_22),
.B2(n_37),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_92),
.B1(n_103),
.B2(n_49),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_57),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_52),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_97),
.A2(n_101),
.B1(n_60),
.B2(n_59),
.Y(n_115)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_106),
.Y(n_123)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

NOR2x1_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_104),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_60),
.A2(n_20),
.B(n_30),
.C(n_3),
.Y(n_103)
);

INVx6_ASAP7_75t_SL g104 ( 
.A(n_67),
.Y(n_104)
);

AO22x2_ASAP7_75t_L g105 ( 
.A1(n_60),
.A2(n_38),
.B1(n_37),
.B2(n_42),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_67),
.B1(n_65),
.B2(n_17),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_50),
.B(n_19),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_109),
.B(n_116),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_111),
.A2(n_125),
.B(n_72),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_115),
.A2(n_82),
.B1(n_77),
.B2(n_87),
.Y(n_154)
);

AND2x6_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_83),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_56),
.B(n_54),
.C(n_61),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_126),
.B1(n_110),
.B2(n_132),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_120),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_76),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_67),
.C(n_70),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_74),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_124),
.A2(n_92),
.B1(n_103),
.B2(n_90),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_30),
.B(n_50),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_79),
.B(n_34),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_85),
.Y(n_142)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_135),
.B(n_138),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_156),
.B1(n_134),
.B2(n_113),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_139),
.Y(n_173)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_140),
.B(n_141),
.Y(n_181)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_148),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_114),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_143),
.B(n_144),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_91),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_122),
.B(n_73),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_146),
.A2(n_134),
.B1(n_93),
.B2(n_108),
.Y(n_170)
);

BUFx24_ASAP7_75t_SL g147 ( 
.A(n_122),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_147),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_73),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_114),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_149),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_150),
.A2(n_162),
.B(n_163),
.Y(n_185)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_130),
.B(n_104),
.Y(n_152)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_155),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_30),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_98),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_116),
.A2(n_75),
.B1(n_93),
.B2(n_99),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_118),
.C(n_111),
.Y(n_164)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

OA21x2_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_108),
.B(n_100),
.Y(n_176)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_0),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_189),
.C(n_166),
.Y(n_205)
);

XNOR2x1_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_126),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_165),
.A2(n_175),
.B(n_186),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_184),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_169),
.A2(n_182),
.B1(n_187),
.B2(n_25),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_174),
.B1(n_138),
.B2(n_141),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_158),
.A2(n_160),
.B1(n_159),
.B2(n_162),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_96),
.B(n_127),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_176),
.A2(n_31),
.B1(n_25),
.B2(n_19),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_98),
.B1(n_102),
.B2(n_127),
.Y(n_182)
);

AND2x2_ASAP7_75t_SL g184 ( 
.A(n_135),
.B(n_31),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_150),
.A2(n_31),
.B(n_86),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_136),
.A2(n_131),
.B1(n_89),
.B2(n_133),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_137),
.B(n_96),
.C(n_31),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_182),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_190),
.B(n_193),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_192),
.A2(n_196),
.B1(n_198),
.B2(n_203),
.Y(n_213)
);

AOI322xp5_ASAP7_75t_SL g193 ( 
.A1(n_165),
.A2(n_140),
.A3(n_148),
.B1(n_144),
.B2(n_146),
.C1(n_157),
.C2(n_142),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_194),
.B(n_199),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_139),
.Y(n_195)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_174),
.A2(n_161),
.B1(n_31),
.B2(n_25),
.Y(n_196)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_167),
.A2(n_25),
.B1(n_19),
.B2(n_0),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_201),
.A2(n_183),
.B1(n_176),
.B2(n_171),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_202),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_170),
.A2(n_25),
.B1(n_19),
.B2(n_0),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_172),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_204),
.B(n_206),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_211),
.C(n_179),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_172),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_208),
.A2(n_209),
.B1(n_181),
.B2(n_177),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_187),
.A2(n_19),
.B1(n_3),
.B2(n_4),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_210),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_189),
.C(n_166),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_212),
.A2(n_219),
.B1(n_224),
.B2(n_225),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_185),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_221),
.C(n_223),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_218),
.B(n_213),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_190),
.A2(n_207),
.B1(n_206),
.B2(n_169),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_185),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_210),
.A2(n_186),
.B1(n_177),
.B2(n_188),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_188),
.B1(n_171),
.B2(n_180),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_215),
.A2(n_196),
.B1(n_168),
.B2(n_183),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_229),
.B(n_236),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_237),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_211),
.C(n_202),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_233),
.C(n_234),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_202),
.C(n_184),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_184),
.C(n_200),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_184),
.C(n_200),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_240),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_217),
.A2(n_175),
.B(n_181),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_212),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_226),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_228),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_198),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_241),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_209),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_213),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_241),
.A2(n_215),
.B1(n_214),
.B2(n_227),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_244),
.A2(n_203),
.B1(n_232),
.B2(n_230),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_219),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_247),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_239),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_234),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_233),
.Y(n_247)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_250),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_253),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_255),
.B(n_258),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_249),
.A2(n_243),
.B(n_244),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_256),
.A2(n_261),
.B(n_5),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_2),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_5),
.Y(n_265)
);

OAI21xp33_ASAP7_75t_L g261 ( 
.A1(n_247),
.A2(n_2),
.B(n_3),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_248),
.Y(n_262)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_262),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_248),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_264),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_260),
.A2(n_251),
.B1(n_252),
.B2(n_178),
.Y(n_264)
);

MAJx2_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_256),
.C(n_6),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_266),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_270)
);

OAI221xp5_ASAP7_75t_L g272 ( 
.A1(n_268),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_267),
.Y(n_273)
);

AOI322xp5_ASAP7_75t_L g276 ( 
.A1(n_272),
.A2(n_273),
.A3(n_274),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_14),
.Y(n_276)
);

AOI322xp5_ASAP7_75t_L g274 ( 
.A1(n_271),
.A2(n_267),
.A3(n_259),
.B1(n_254),
.B2(n_178),
.C1(n_14),
.C2(n_9),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_273),
.A2(n_269),
.B(n_254),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_276),
.C(n_11),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_16),
.C(n_277),
.Y(n_279)
);


endmodule