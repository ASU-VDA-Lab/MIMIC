module fake_jpeg_15398_n_65 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_65);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_65;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_56;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_7),
.B(n_6),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_3),
.B(n_6),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_19),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_20),
.A2(n_17),
.B1(n_24),
.B2(n_25),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_9),
.B(n_0),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_23),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g22 ( 
.A1(n_12),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_11),
.B1(n_15),
.B2(n_17),
.Y(n_28)
);

OR2x2_ASAP7_75t_SL g23 ( 
.A(n_13),
.B(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_10),
.B(n_13),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_17),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_21),
.A2(n_16),
.B1(n_18),
.B2(n_15),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_28),
.B1(n_38),
.B2(n_32),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_14),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_33),
.C(n_34),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_14),
.C(n_15),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_19),
.B(n_22),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_18),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_28),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

OA21x2_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_35),
.B(n_38),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_21),
.A2(n_16),
.B1(n_23),
.B2(n_22),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_44),
.B1(n_46),
.B2(n_29),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_34),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_33),
.C(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_43),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_47),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_SL g57 ( 
.A(n_49),
.B(n_53),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

OAI221xp5_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_41),
.B1(n_40),
.B2(n_46),
.C(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_54),
.B(n_56),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_49),
.B(n_45),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_53),
.A2(n_46),
.B1(n_40),
.B2(n_43),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_48),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_51),
.B(n_31),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_50),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_63),
.B(n_55),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_62),
.B(n_61),
.Y(n_65)
);


endmodule