module fake_jpeg_25461_n_297 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_297);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_245;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_32),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_46),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_18),
.B1(n_25),
.B2(n_14),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_16),
.B1(n_26),
.B2(n_33),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_31),
.B1(n_18),
.B2(n_25),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_50),
.A2(n_52),
.B1(n_55),
.B2(n_58),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_31),
.B1(n_18),
.B2(n_35),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_34),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_18),
.B1(n_15),
.B2(n_24),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_14),
.B1(n_26),
.B2(n_16),
.Y(n_53)
);

OAI22x1_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_27),
.B1(n_34),
.B2(n_29),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_35),
.B1(n_14),
.B2(n_26),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_57),
.Y(n_70)
);

INVxp67_ASAP7_75t_SL g57 ( 
.A(n_45),
.Y(n_57)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_66),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_67),
.B(n_47),
.Y(n_74)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_37),
.B1(n_34),
.B2(n_30),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_82),
.B(n_62),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_36),
.Y(n_77)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_78),
.B(n_79),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_39),
.C(n_43),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_90),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_62),
.B(n_16),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_58),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_83),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_86),
.B1(n_56),
.B2(n_69),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_88),
.A2(n_56),
.B1(n_59),
.B2(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_98),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_95),
.A2(n_105),
.B(n_115),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_99),
.B1(n_114),
.B2(n_87),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_90),
.B1(n_72),
.B2(n_81),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_97),
.A2(n_104),
.B1(n_110),
.B2(n_54),
.Y(n_126)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_78),
.A2(n_50),
.B1(n_67),
.B2(n_64),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_106),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_12),
.C(n_11),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_64),
.B1(n_68),
.B2(n_37),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_73),
.A2(n_0),
.B(n_1),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_29),
.Y(n_127)
);

OA21x2_ASAP7_75t_L g109 ( 
.A1(n_73),
.A2(n_30),
.B(n_29),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_28),
.B(n_17),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_68),
.B1(n_59),
.B2(n_33),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVxp33_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

OAI32xp33_ASAP7_75t_L g113 ( 
.A1(n_76),
.A2(n_36),
.A3(n_19),
.B1(n_21),
.B2(n_13),
.Y(n_113)
);

OAI32xp33_ASAP7_75t_L g122 ( 
.A1(n_113),
.A2(n_89),
.A3(n_91),
.B1(n_87),
.B2(n_30),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_76),
.A2(n_33),
.B1(n_54),
.B2(n_13),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_1),
.B(n_2),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_117),
.B(n_127),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_112),
.A2(n_85),
.B1(n_80),
.B2(n_75),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_136),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_103),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_119),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_89),
.C(n_80),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_143),
.C(n_22),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

AO22x1_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_28),
.B1(n_17),
.B2(n_3),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_123),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_126),
.A2(n_128),
.B1(n_136),
.B2(n_113),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_97),
.A2(n_27),
.B1(n_22),
.B2(n_13),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_130),
.Y(n_169)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_108),
.Y(n_132)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_135),
.Y(n_145)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_95),
.A2(n_22),
.B1(n_27),
.B2(n_17),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_1),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_21),
.Y(n_138)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_135),
.B(n_131),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_98),
.B(n_21),
.Y(n_140)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_103),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_141),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_105),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_142),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_22),
.C(n_28),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_19),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_104),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_SL g146 ( 
.A1(n_130),
.A2(n_133),
.B(n_129),
.C(n_115),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_146),
.A2(n_155),
.B(n_164),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_149),
.B(n_126),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_150),
.A2(n_123),
.B1(n_122),
.B2(n_140),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_166),
.C(n_143),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_156),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_119),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_141),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_163),
.Y(n_183)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_162),
.Y(n_193)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_12),
.Y(n_165)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_11),
.C(n_10),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_168),
.A2(n_128),
.B1(n_142),
.B2(n_116),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_170),
.A2(n_171),
.B(n_173),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_131),
.A2(n_2),
.B(n_3),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_174),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_139),
.A2(n_4),
.B(n_5),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_124),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_176),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_124),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_178),
.B(n_186),
.Y(n_223)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_182),
.Y(n_212)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_185),
.Y(n_217)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_195),
.Y(n_204)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_194),
.A2(n_199),
.B1(n_150),
.B2(n_198),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_144),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_196),
.A2(n_198),
.B1(n_202),
.B2(n_172),
.Y(n_216)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_152),
.B(n_134),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_166),
.C(n_138),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_157),
.B(n_116),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_171),
.Y(n_214)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

XNOR2x1_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_146),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_SL g226 ( 
.A(n_203),
.B(n_209),
.C(n_216),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_160),
.C(n_175),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_211),
.C(n_215),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_160),
.C(n_157),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_213),
.A2(n_194),
.B1(n_179),
.B2(n_186),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_218),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_163),
.C(n_158),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_158),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_219),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_185),
.C(n_182),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_220),
.B(n_222),
.Y(n_236)
);

OA21x2_ASAP7_75t_L g221 ( 
.A1(n_177),
.A2(n_188),
.B(n_197),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_221),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_162),
.C(n_161),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_203),
.A2(n_197),
.B(n_179),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_224),
.A2(n_207),
.B(n_173),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_183),
.Y(n_225)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_225),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_227),
.A2(n_235),
.B1(n_221),
.B2(n_211),
.Y(n_244)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_232),
.Y(n_243)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_221),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_240),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_208),
.A2(n_191),
.B1(n_187),
.B2(n_199),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_154),
.Y(n_239)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_239),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_212),
.Y(n_240)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_230),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_252),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_244),
.A2(n_226),
.B1(n_227),
.B2(n_224),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_204),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_251),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_239),
.Y(n_248)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_248),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_214),
.Y(n_249)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_249),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_204),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_215),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_236),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_254),
.B(n_248),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_229),
.B1(n_223),
.B2(n_231),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_256),
.B(n_264),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_154),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_180),
.Y(n_259)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_259),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_237),
.C(n_235),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_261),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_240),
.C(n_218),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_147),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_262),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_243),
.A2(n_226),
.B(n_147),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_265),
.B(n_252),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_265),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_258),
.B(n_250),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_268),
.B(n_275),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_245),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_271),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_274),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_125),
.B(n_5),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_4),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_263),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_282),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_280),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_257),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_4),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_283),
.A2(n_267),
.B(n_8),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_6),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_284),
.A2(n_272),
.B(n_7),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_288),
.C(n_289),
.Y(n_290)
);

AO21x1_ASAP7_75t_L g288 ( 
.A1(n_281),
.A2(n_267),
.B(n_8),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_279),
.C(n_8),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_279),
.C(n_286),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_292),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_290),
.A2(n_6),
.B(n_8),
.Y(n_293)
);

A2O1A1Ixp33_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_9),
.B(n_293),
.C(n_285),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_9),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_9),
.Y(n_297)
);


endmodule