module fake_ariane_3130_n_5595 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_598, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_631, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_635, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_620, n_228, n_325, n_276, n_93, n_636, n_427, n_108, n_587, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_588, n_638, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_579, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_616, n_617, n_630, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_601, n_565, n_281, n_24, n_7, n_628, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_575, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_451, n_613, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_629, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_67, n_509, n_583, n_306, n_313, n_92, n_430, n_626, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_615, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_624, n_118, n_121, n_618, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_573, n_127, n_531, n_5595);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_616;
input n_617;
input n_630;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_601;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_575;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_451;
input n_613;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_629;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_583;
input n_306;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_615;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_624;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;

output n_5595;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_4030;
wire n_4770;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_2679;
wire n_5402;
wire n_2182;
wire n_5553;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_4962;
wire n_1430;
wire n_2002;
wire n_1238;
wire n_2729;
wire n_4302;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_864;
wire n_5302;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_2790;
wire n_2207;
wire n_3954;
wire n_4982;
wire n_2042;
wire n_1131;
wire n_5479;
wire n_2646;
wire n_737;
wire n_2653;
wire n_4610;
wire n_3115;
wire n_4028;
wire n_5263;
wire n_5565;
wire n_2482;
wire n_1682;
wire n_958;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_5590;
wire n_2621;
wire n_4853;
wire n_1909;
wire n_5229;
wire n_4260;
wire n_903;
wire n_3348;
wire n_3261;
wire n_1761;
wire n_1690;
wire n_2807;
wire n_1018;
wire n_4512;
wire n_4132;
wire n_1364;
wire n_2390;
wire n_4500;
wire n_2322;
wire n_1107;
wire n_2663;
wire n_5481;
wire n_4824;
wire n_5340;
wire n_3545;
wire n_1428;
wire n_1284;
wire n_4741;
wire n_1241;
wire n_4143;
wire n_4273;
wire n_901;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_1519;
wire n_4567;
wire n_786;
wire n_3552;
wire n_2950;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_5589;
wire n_3015;
wire n_3870;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_3482;
wire n_5403;
wire n_823;
wire n_1900;
wire n_4268;
wire n_863;
wire n_3960;
wire n_2433;
wire n_899;
wire n_3975;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_3325;
wire n_661;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_1811;
wire n_3612;
wire n_4505;
wire n_1840;
wire n_5247;
wire n_5464;
wire n_4476;
wire n_844;
wire n_1267;
wire n_2956;
wire n_5210;
wire n_1213;
wire n_2382;
wire n_780;
wire n_5292;
wire n_1918;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_1140;
wire n_3458;
wire n_3511;
wire n_2077;
wire n_1121;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_1216;
wire n_4908;
wire n_3754;
wire n_5060;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_5391;
wire n_5452;
wire n_3359;
wire n_3841;
wire n_5249;
wire n_851;
wire n_3900;
wire n_3413;
wire n_5076;
wire n_3539;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_930;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_5046;
wire n_1386;
wire n_3506;
wire n_4827;
wire n_1842;
wire n_4993;
wire n_3678;
wire n_2791;
wire n_1661;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_966;
wire n_992;
wire n_3549;
wire n_3914;
wire n_5586;
wire n_1692;
wire n_2611;
wire n_5468;
wire n_3029;
wire n_4745;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5056;
wire n_1178;
wire n_2015;
wire n_5204;
wire n_2877;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_2161;
wire n_746;
wire n_1357;
wire n_1787;
wire n_1389;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_4905;
wire n_4508;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_3614;
wire n_959;
wire n_2257;
wire n_1101;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_5179;
wire n_2435;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_5549;
wire n_1087;
wire n_2388;
wire n_2273;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_3700;
wire n_4307;
wire n_2795;
wire n_1841;
wire n_1680;
wire n_2954;
wire n_4438;
wire n_974;
wire n_3814;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_4195;
wire n_5091;
wire n_4866;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_698;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_5454;
wire n_1209;
wire n_4254;
wire n_646;
wire n_3438;
wire n_2625;
wire n_5373;
wire n_1578;
wire n_3147;
wire n_3661;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_1568;
wire n_2919;
wire n_3108;
wire n_2632;
wire n_5557;
wire n_4314;
wire n_2980;
wire n_1728;
wire n_4315;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_4857;
wire n_1651;
wire n_3087;
wire n_4637;
wire n_5523;
wire n_2697;
wire n_1263;
wire n_1817;
wire n_3704;
wire n_670;
wire n_2677;
wire n_4296;
wire n_2483;
wire n_5088;
wire n_1032;
wire n_1592;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_1743;
wire n_720;
wire n_1943;
wire n_5138;
wire n_4588;
wire n_5149;
wire n_1163;
wire n_3054;
wire n_4970;
wire n_5280;
wire n_4153;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_2373;
wire n_3881;
wire n_5089;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_2617;
wire n_808;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_3466;
wire n_2074;
wire n_5031;
wire n_1665;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_2117;
wire n_1053;
wire n_5296;
wire n_5398;
wire n_1906;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_1828;
wire n_1304;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_1349;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_3370;
wire n_874;
wire n_3949;
wire n_2286;
wire n_5192;
wire n_4247;
wire n_707;
wire n_5051;
wire n_5336;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_1015;
wire n_1162;
wire n_4292;
wire n_2118;
wire n_688;
wire n_1490;
wire n_5552;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_1086;
wire n_3025;
wire n_3051;
wire n_986;
wire n_2802;
wire n_1104;
wire n_887;
wire n_2125;
wire n_1156;
wire n_4974;
wire n_5123;
wire n_2861;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_1498;
wire n_1188;
wire n_4856;
wire n_2618;
wire n_4216;
wire n_957;
wire n_1242;
wire n_2707;
wire n_2849;
wire n_1489;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_3713;
wire n_1863;
wire n_5536;
wire n_4798;
wire n_1500;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_1189;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_3214;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5539;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_1957;
wire n_1953;
wire n_1219;
wire n_710;
wire n_3944;
wire n_4729;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_4800;
wire n_1373;
wire n_1540;
wire n_5427;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_5450;
wire n_832;
wire n_744;
wire n_2821;
wire n_3696;
wire n_1331;
wire n_4781;
wire n_1529;
wire n_3531;
wire n_5124;
wire n_655;
wire n_4237;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_1007;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_2448;
wire n_2211;
wire n_951;
wire n_5318;
wire n_5374;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_722;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_5463;
wire n_1338;
wire n_2978;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_704;
wire n_2958;
wire n_1044;
wire n_1714;
wire n_4429;
wire n_5435;
wire n_3340;
wire n_5053;
wire n_5476;
wire n_5483;
wire n_1243;
wire n_5511;
wire n_3486;
wire n_2457;
wire n_2992;
wire n_3197;
wire n_3256;
wire n_1878;
wire n_3646;
wire n_2520;
wire n_811;
wire n_791;
wire n_3864;
wire n_4694;
wire n_1025;
wire n_4664;
wire n_3450;
wire n_687;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_642;
wire n_1406;
wire n_5073;
wire n_4306;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_695;
wire n_2991;
wire n_5419;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_2723;
wire n_1476;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_678;
wire n_651;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_3780;
wire n_1657;
wire n_3753;
wire n_1488;
wire n_4846;
wire n_1330;
wire n_906;
wire n_2295;
wire n_5225;
wire n_4076;
wire n_3142;
wire n_3129;
wire n_3495;
wire n_3843;
wire n_4805;
wire n_2606;
wire n_2386;
wire n_4822;
wire n_1829;
wire n_4635;
wire n_1450;
wire n_5532;
wire n_3740;
wire n_5441;
wire n_2417;
wire n_1815;
wire n_1493;
wire n_2911;
wire n_3313;
wire n_2354;
wire n_4281;
wire n_3945;
wire n_3726;
wire n_4419;
wire n_5405;
wire n_1256;
wire n_5365;
wire n_3560;
wire n_3345;
wire n_3421;
wire n_1448;
wire n_1009;
wire n_3548;
wire n_4906;
wire n_4630;
wire n_4829;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_1995;
wire n_1397;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_4966;
wire n_2250;
wire n_1117;
wire n_3321;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_2506;
wire n_2413;
wire n_4825;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_2626;
wire n_2892;
wire n_2605;
wire n_2804;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_1035;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_2044;
wire n_3886;
wire n_825;
wire n_732;
wire n_2619;
wire n_1192;
wire n_5141;
wire n_3098;
wire n_4503;
wire n_1291;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_3386;
wire n_3921;
wire n_2177;
wire n_2766;
wire n_4196;
wire n_1197;
wire n_2613;
wire n_1517;
wire n_2647;
wire n_5508;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_1671;
wire n_5027;
wire n_2343;
wire n_1048;
wire n_775;
wire n_667;
wire n_3380;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2411;
wire n_4631;
wire n_1504;
wire n_2110;
wire n_5377;
wire n_3822;
wire n_889;
wire n_4355;
wire n_3818;
wire n_3587;
wire n_2608;
wire n_1948;
wire n_4155;
wire n_810;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_3497;
wire n_4542;
wire n_5451;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_5460;
wire n_4685;
wire n_3927;
wire n_2068;
wire n_3595;
wire n_1194;
wire n_4060;
wire n_1647;
wire n_1454;
wire n_2459;
wire n_941;
wire n_3396;
wire n_5517;
wire n_5426;
wire n_4093;
wire n_4123;
wire n_4294;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_5587;
wire n_4722;
wire n_3048;
wire n_3339;
wire n_4164;
wire n_4126;
wire n_5030;
wire n_2963;
wire n_2561;
wire n_1056;
wire n_5584;
wire n_674;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_848;
wire n_5125;
wire n_4922;
wire n_4733;
wire n_1814;
wire n_2441;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_4509;
wire n_4935;
wire n_2073;
wire n_4004;
wire n_5238;
wire n_750;
wire n_834;
wire n_3630;
wire n_1612;
wire n_800;
wire n_1910;
wire n_2189;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_724;
wire n_2931;
wire n_3433;
wire n_5556;
wire n_3597;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_3786;
wire n_875;
wire n_2828;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_4204;
wire n_3553;
wire n_5323;
wire n_3645;
wire n_793;
wire n_4996;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_3550;
wire n_5510;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1805;
wire n_4068;
wire n_5440;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_2443;
wire n_3610;
wire n_5011;
wire n_1554;
wire n_3279;
wire n_5513;
wire n_972;
wire n_4262;
wire n_2923;
wire n_2843;
wire n_3714;
wire n_4832;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_1679;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_3125;
wire n_5128;
wire n_2356;
wire n_4672;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_783;
wire n_4053;
wire n_1127;
wire n_1008;
wire n_3963;
wire n_3091;
wire n_1024;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_936;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_1525;
wire n_4628;
wire n_1775;
wire n_908;
wire n_1036;
wire n_4083;
wire n_1270;
wire n_1272;
wire n_2794;
wire n_2901;
wire n_3940;
wire n_3225;
wire n_3621;
wire n_5529;
wire n_3473;
wire n_3680;
wire n_3565;
wire n_5388;
wire n_5354;
wire n_2453;
wire n_3331;
wire n_1788;
wire n_2138;
wire n_3040;
wire n_4230;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_2000;
wire n_5276;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_917;
wire n_5196;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2215;
wire n_3847;
wire n_4073;
wire n_1261;
wire n_3633;
wire n_857;
wire n_1235;
wire n_2584;
wire n_4001;
wire n_1462;
wire n_1064;
wire n_1446;
wire n_1701;
wire n_3111;
wire n_731;
wire n_1813;
wire n_2997;
wire n_1573;
wire n_3258;
wire n_758;
wire n_3691;
wire n_2252;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_4339;
wire n_4690;
wire n_2987;
wire n_1473;
wire n_1076;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_2522;
wire n_3632;
wire n_1344;
wire n_4064;
wire n_3351;
wire n_5478;
wire n_1141;
wire n_3457;
wire n_5384;
wire n_840;
wire n_2324;
wire n_5283;
wire n_3454;
wire n_2139;
wire n_2521;
wire n_2740;
wire n_1991;
wire n_4066;
wire n_4681;
wire n_3303;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_1113;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_1265;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_1409;
wire n_1684;
wire n_1148;
wire n_1588;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_3018;
wire n_1875;
wire n_2429;
wire n_5286;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_1039;
wire n_5040;
wire n_1150;
wire n_4266;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_1136;
wire n_1190;
wire n_3628;
wire n_4777;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_5399;
wire n_658;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_3872;
wire n_4415;
wire n_5110;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_3441;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_708;
wire n_2545;
wire n_2513;
wire n_4408;
wire n_2115;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_860;
wire n_3555;
wire n_3534;
wire n_4548;
wire n_2670;
wire n_3556;
wire n_896;
wire n_4574;
wire n_2644;
wire n_4557;
wire n_3071;
wire n_1698;
wire n_1337;
wire n_774;
wire n_2148;
wire n_5548;
wire n_1168;
wire n_4663;
wire n_3296;
wire n_3794;
wire n_3762;
wire n_4624;
wire n_656;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_4686;
wire n_2384;
wire n_1705;
wire n_768;
wire n_3707;
wire n_3895;
wire n_1091;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_2058;
wire n_3231;
wire n_1846;
wire n_4161;
wire n_5304;
wire n_5437;
wire n_1581;
wire n_3058;
wire n_757;
wire n_2047;
wire n_946;
wire n_1655;
wire n_3709;
wire n_3398;
wire n_1146;
wire n_5355;
wire n_998;
wire n_3592;
wire n_5321;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_4772;
wire n_1368;
wire n_963;
wire n_4120;
wire n_925;
wire n_2880;
wire n_1313;
wire n_1001;
wire n_3722;
wire n_4716;
wire n_4654;
wire n_1115;
wire n_1339;
wire n_1051;
wire n_5116;
wire n_3771;
wire n_719;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_1010;
wire n_2830;
wire n_5500;
wire n_4622;
wire n_4757;
wire n_1871;
wire n_803;
wire n_4016;
wire n_3334;
wire n_2940;
wire n_3427;
wire n_3162;
wire n_5569;
wire n_4591;
wire n_5515;
wire n_3083;
wire n_4570;
wire n_2491;
wire n_1931;
wire n_5559;
wire n_2259;
wire n_5337;
wire n_849;
wire n_5059;
wire n_4655;
wire n_1820;
wire n_1233;
wire n_4493;
wire n_1808;
wire n_1635;
wire n_1704;
wire n_4896;
wire n_4851;
wire n_2479;
wire n_886;
wire n_1308;
wire n_1451;
wire n_1487;
wire n_675;
wire n_5528;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_2484;
wire n_5358;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_1355;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2334;
wire n_5467;
wire n_1169;
wire n_789;
wire n_3181;
wire n_5493;
wire n_1916;
wire n_4602;
wire n_1713;
wire n_2818;
wire n_1436;
wire n_4900;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1566;
wire n_2837;
wire n_717;
wire n_952;
wire n_2446;
wire n_4116;
wire n_5360;
wire n_2671;
wire n_2702;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_4103;
wire n_2529;
wire n_2374;
wire n_5439;
wire n_1225;
wire n_3154;
wire n_1366;
wire n_3938;
wire n_2278;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_4439;
wire n_870;
wire n_4985;
wire n_3382;
wire n_3930;
wire n_3808;
wire n_5471;
wire n_2248;
wire n_813;
wire n_4660;
wire n_3081;
wire n_5497;
wire n_5519;
wire n_995;
wire n_2579;
wire n_1961;
wire n_1535;
wire n_2960;
wire n_3270;
wire n_871;
wire n_2844;
wire n_1979;
wire n_829;
wire n_4814;
wire n_2221;
wire n_5502;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_3657;
wire n_2634;
wire n_2746;
wire n_645;
wire n_5098;
wire n_721;
wire n_1084;
wire n_1276;
wire n_5145;
wire n_2878;
wire n_3830;
wire n_3252;
wire n_5466;
wire n_1528;
wire n_3315;
wire n_3523;
wire n_3999;
wire n_3420;
wire n_3859;
wire n_868;
wire n_5213;
wire n_3474;
wire n_2458;
wire n_5592;
wire n_3150;
wire n_5491;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1636;
wire n_4597;
wire n_4546;
wire n_5187;
wire n_4031;
wire n_5119;
wire n_1254;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_3571;
wire n_4576;
wire n_3297;
wire n_5148;
wire n_3003;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_5330;
wire n_1560;
wire n_2899;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5526;
wire n_5202;
wire n_3817;
wire n_2722;
wire n_3728;
wire n_5107;
wire n_4680;
wire n_5067;
wire n_1012;
wire n_2061;
wire n_2685;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_1443;
wire n_5264;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_705;
wire n_4593;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_3554;
wire n_2717;
wire n_1391;
wire n_2981;
wire n_1006;
wire n_4995;
wire n_1159;
wire n_4498;
wire n_772;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_676;
wire n_3758;
wire n_5423;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_1872;
wire n_1585;
wire n_3767;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_2216;
wire n_2426;
wire n_652;
wire n_4850;
wire n_1260;
wire n_3716;
wire n_2926;
wire n_4937;
wire n_798;
wire n_5574;
wire n_3391;
wire n_912;
wire n_4786;
wire n_5203;
wire n_4354;
wire n_4235;
wire n_3159;
wire n_2855;
wire n_794;
wire n_2848;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_1292;
wire n_1026;
wire n_3460;
wire n_1610;
wire n_5155;
wire n_2202;
wire n_2952;
wire n_3530;
wire n_2693;
wire n_5408;
wire n_5540;
wire n_3240;
wire n_5066;
wire n_931;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_967;
wire n_5130;
wire n_4175;
wire n_1079;
wire n_5200;
wire n_3393;
wire n_2836;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_2172;
wire n_2601;
wire n_1880;
wire n_2365;
wire n_1399;
wire n_1855;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_5413;
wire n_1903;
wire n_2147;
wire n_4020;
wire n_5150;
wire n_5111;
wire n_2224;
wire n_1226;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_3046;
wire n_2921;
wire n_1240;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_5444;
wire n_3257;
wire n_3730;
wire n_3979;
wire n_5097;
wire n_2695;
wire n_2598;
wire n_3727;
wire n_976;
wire n_4003;
wire n_1832;
wire n_767;
wire n_2302;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_3342;
wire n_2895;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_5550;
wire n_3375;
wire n_2768;
wire n_3760;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_5457;
wire n_5159;
wire n_4022;
wire n_1020;
wire n_2495;
wire n_1058;
wire n_4336;
wire n_5314;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_1279;
wire n_2511;
wire n_3981;
wire n_2681;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_3031;
wire n_2335;
wire n_5482;
wire n_3215;
wire n_1401;
wire n_3138;
wire n_776;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_4494;
wire n_4201;
wire n_5287;
wire n_4719;
wire n_3577;
wire n_4074;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_1217;
wire n_2662;
wire n_4386;
wire n_3917;
wire n_1231;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_5524;
wire n_926;
wire n_2296;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_4225;
wire n_4658;
wire n_4186;
wire n_1501;
wire n_2241;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_1570;
wire n_3377;
wire n_1518;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_855;
wire n_2059;
wire n_4713;
wire n_1287;
wire n_1611;
wire n_3374;
wire n_4870;
wire n_4818;
wire n_4916;
wire n_4323;
wire n_1899;
wire n_5376;
wire n_3508;
wire n_4129;
wire n_5488;
wire n_1105;
wire n_3599;
wire n_4480;
wire n_3734;
wire n_3401;
wire n_983;
wire n_699;
wire n_3542;
wire n_3263;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_1377;
wire n_1614;
wire n_5328;
wire n_3819;
wire n_3222;
wire n_1740;
wire n_4616;
wire n_5016;
wire n_5470;
wire n_1092;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_1963;
wire n_3868;
wire n_729;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_5362;
wire n_2754;
wire n_4580;
wire n_1218;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_877;
wire n_3995;
wire n_3908;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_1089;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_3216;
wire n_3568;
wire n_2555;
wire n_2708;
wire n_735;
wire n_4844;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_845;
wire n_1649;
wire n_2470;
wire n_1297;
wire n_3551;
wire n_1708;
wire n_5037;
wire n_5581;
wire n_4677;
wire n_5189;
wire n_4525;
wire n_3364;
wire n_2643;
wire n_755;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_4369;
wire n_3826;
wire n_2266;
wire n_4324;
wire n_842;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_742;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_769;
wire n_3671;
wire n_2366;
wire n_1753;
wire n_5484;
wire n_1372;
wire n_1895;
wire n_4104;
wire n_982;
wire n_3791;
wire n_915;
wire n_2008;
wire n_4989;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_3151;
wire n_3016;
wire n_2460;
wire n_1319;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_659;
wire n_1332;
wire n_5385;
wire n_1747;
wire n_3990;
wire n_1171;
wire n_4069;
wire n_3582;
wire n_4280;
wire n_1867;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_4811;
wire n_2696;
wire n_5256;
wire n_4779;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_1400;
wire n_3735;
wire n_1527;
wire n_1513;
wire n_3656;
wire n_4524;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_5568;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1257;
wire n_1954;
wire n_3964;
wire n_5364;
wire n_3302;
wire n_2486;
wire n_1897;
wire n_5469;
wire n_2137;
wire n_3685;
wire n_4977;
wire n_2492;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_5021;
wire n_1449;
wire n_2900;
wire n_797;
wire n_2912;
wire n_1405;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_1757;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_3124;
wire n_3811;
wire n_4200;
wire n_2249;
wire n_3411;
wire n_5222;
wire n_3463;
wire n_2785;
wire n_730;
wire n_4938;
wire n_2574;
wire n_1281;
wire n_2364;
wire n_1856;
wire n_1524;
wire n_2928;
wire n_5505;
wire n_1118;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_1293;
wire n_961;
wire n_726;
wire n_5504;
wire n_878;
wire n_4118;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_3157;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_5129;
wire n_806;
wire n_1350;
wire n_4704;
wire n_2720;
wire n_649;
wire n_1561;
wire n_5494;
wire n_2405;
wire n_2700;
wire n_1616;
wire n_2416;
wire n_2064;
wire n_3640;
wire n_5161;
wire n_1557;
wire n_4744;
wire n_5378;
wire n_4706;
wire n_2022;
wire n_3879;
wire n_4343;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_5389;
wire n_4990;
wire n_2986;
wire n_949;
wire n_2454;
wire n_3591;
wire n_2760;
wire n_4919;
wire n_1208;
wire n_3317;
wire n_4835;
wire n_1151;
wire n_4420;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_5266;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_1133;
wire n_883;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_4162;
wire n_5293;
wire n_779;
wire n_4790;
wire n_4173;
wire n_5309;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_1269;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_3654;
wire n_1047;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_1288;
wire n_2173;
wire n_3982;
wire n_3647;
wire n_1143;
wire n_3973;
wire n_4799;
wire n_4534;
wire n_4960;
wire n_1153;
wire n_1103;
wire n_5594;
wire n_3738;
wire n_894;
wire n_1380;
wire n_2020;
wire n_2310;
wire n_3600;
wire n_1023;
wire n_914;
wire n_689;
wire n_5382;
wire n_4327;
wire n_3190;
wire n_3027;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_3733;
wire n_1165;
wire n_3967;
wire n_4370;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_1417;
wire n_3096;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_2234;
wire n_1341;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_1603;
wire n_4478;
wire n_2935;
wire n_4246;
wire n_715;
wire n_1066;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_685;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_4754;
wire n_1534;
wire n_1290;
wire n_4375;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_3117;
wire n_4684;
wire n_743;
wire n_1546;
wire n_3384;
wire n_5279;
wire n_2592;
wire n_3490;
wire n_962;
wire n_5043;
wire n_4241;
wire n_1622;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_918;
wire n_1968;
wire n_639;
wire n_5020;
wire n_673;
wire n_2842;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_5232;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_1193;
wire n_1345;
wire n_5035;
wire n_3037;
wire n_1336;
wire n_1033;
wire n_5453;
wire n_4333;
wire n_5339;
wire n_5443;
wire n_1166;
wire n_2007;
wire n_3363;
wire n_1158;
wire n_1803;
wire n_872;
wire n_3522;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_3481;
wire n_5101;
wire n_2236;
wire n_692;
wire n_4457;
wire n_2150;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_3305;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_3354;
wire n_2204;
wire n_1481;
wire n_2040;
wire n_2151;
wire n_2455;
wire n_827;
wire n_3437;
wire n_2231;
wire n_4212;
wire n_4584;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_4110;
wire n_5182;
wire n_1221;
wire n_4217;
wire n_5277;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_1579;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_923;
wire n_1124;
wire n_1326;
wire n_3969;
wire n_2282;
wire n_4605;
wire n_981;
wire n_3873;
wire n_4649;
wire n_1204;
wire n_2428;
wire n_994;
wire n_1360;
wire n_2858;
wire n_3076;
wire n_3410;
wire n_5415;
wire n_856;
wire n_4999;
wire n_4592;
wire n_1564;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_1411;
wire n_1359;
wire n_3536;
wire n_1721;
wire n_3782;
wire n_1317;
wire n_3594;
wire n_5383;
wire n_2385;
wire n_1980;
wire n_4177;
wire n_2501;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_2028;
wire n_919;
wire n_3114;
wire n_2092;
wire n_3622;
wire n_2817;
wire n_2773;
wire n_2402;
wire n_1458;
wire n_679;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_5512;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_2392;
wire n_3272;
wire n_3122;
wire n_3687;
wire n_2787;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2770;
wire n_4550;
wire n_4347;
wire n_702;
wire n_5193;
wire n_4933;
wire n_968;
wire n_4144;
wire n_5514;
wire n_2375;
wire n_3278;
wire n_5579;
wire n_4167;
wire n_3608;
wire n_4895;
wire n_1282;
wire n_4726;
wire n_5573;
wire n_5143;
wire n_1755;
wire n_5188;
wire n_5049;
wire n_2212;
wire n_5308;
wire n_4434;
wire n_5068;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_816;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_5057;
wire n_5425;
wire n_5273;
wire n_2469;
wire n_1125;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_3068;
wire n_1629;
wire n_1094;
wire n_1510;
wire n_3002;
wire n_1099;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_759;
wire n_4156;
wire n_1727;
wire n_3693;
wire n_3132;
wire n_5002;
wire n_5487;
wire n_5531;
wire n_831;
wire n_3681;
wire n_3970;
wire n_778;
wire n_2351;
wire n_1619;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_1152;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_1236;
wire n_4579;
wire n_4776;
wire n_671;
wire n_2704;
wire n_1334;
wire n_3729;
wire n_4471;
wire n_4392;
wire n_3103;
wire n_2048;
wire n_3028;
wire n_4691;
wire n_3148;
wire n_3775;
wire n_684;
wire n_5461;
wire n_3966;
wire n_4397;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_4165;
wire n_2056;
wire n_2852;
wire n_2515;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1941;
wire n_3637;
wire n_1017;
wire n_734;
wire n_4893;
wire n_2240;
wire n_4258;
wire n_709;
wire n_2917;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_5033;
wire n_1686;
wire n_4232;
wire n_5075;
wire n_2097;
wire n_662;
wire n_3461;
wire n_1410;
wire n_2297;
wire n_939;
wire n_4203;
wire n_5400;
wire n_1325;
wire n_1223;
wire n_5347;
wire n_2957;
wire n_1983;
wire n_4767;
wire n_4569;
wire n_948;
wire n_3820;
wire n_5144;
wire n_3072;
wire n_2961;
wire n_4468;
wire n_5509;
wire n_1923;
wire n_3848;
wire n_3631;
wire n_5169;
wire n_4885;
wire n_1479;
wire n_4698;
wire n_1031;
wire n_3674;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_5349;
wire n_3763;
wire n_933;
wire n_3499;
wire n_5534;
wire n_1821;
wire n_3947;
wire n_3910;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_1186;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_4556;
wire n_2205;
wire n_2183;
wire n_1724;
wire n_3088;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_1126;
wire n_5079;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_895;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_5039;
wire n_1818;
wire n_4265;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_1583;
wire n_4612;
wire n_5375;
wire n_5438;
wire n_1264;
wire n_4958;
wire n_1827;
wire n_4149;
wire n_1752;
wire n_2361;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_5563;
wire n_3075;
wire n_1102;
wire n_2239;
wire n_1296;
wire n_4730;
wire n_4421;
wire n_2464;
wire n_3697;
wire n_882;
wire n_2304;
wire n_2514;
wire n_1299;
wire n_3430;
wire n_2063;
wire n_3489;
wire n_5012;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_4971;
wire n_2095;
wire n_2738;
wire n_2590;
wire n_4661;
wire n_3041;
wire n_2797;
wire n_1421;
wire n_2423;
wire n_2208;
wire n_5422;
wire n_5246;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_1069;
wire n_4305;
wire n_2037;
wire n_2953;
wire n_2823;
wire n_3684;
wire n_5404;
wire n_913;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_5332;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_3268;
wire n_2559;
wire n_1383;
wire n_4259;
wire n_2030;
wire n_850;
wire n_4299;
wire n_2407;
wire n_690;
wire n_5367;
wire n_2243;
wire n_5288;
wire n_2694;
wire n_3742;
wire n_4965;
wire n_1837;
wire n_4178;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_5294;
wire n_5570;
wire n_2731;
wire n_3703;
wire n_5411;
wire n_1246;
wire n_5265;
wire n_2123;
wire n_2238;
wire n_4793;
wire n_4802;
wire n_1196;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_4897;
wire n_1298;
wire n_1745;
wire n_4674;
wire n_4796;
wire n_1088;
wire n_766;
wire n_5184;
wire n_2750;
wire n_2547;
wire n_945;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_3281;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_4589;
wire n_3220;
wire n_4581;
wire n_665;
wire n_4625;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_738;
wire n_5575;
wire n_672;
wire n_4968;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_3856;
wire n_4038;
wire n_5316;
wire n_2735;
wire n_953;
wire n_4214;
wire n_1888;
wire n_5290;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_3419;
wire n_989;
wire n_5048;
wire n_2233;
wire n_5363;
wire n_795;
wire n_4892;
wire n_1936;
wire n_3890;
wire n_821;
wire n_770;
wire n_1514;
wire n_2782;
wire n_3929;
wire n_971;
wire n_4353;
wire n_2201;
wire n_4950;
wire n_1650;
wire n_4176;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_4488;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_4608;
wire n_3948;
wire n_4839;
wire n_1074;
wire n_1765;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_2332;
wire n_2391;
wire n_2060;
wire n_1295;
wire n_3883;
wire n_1013;
wire n_4032;
wire n_2571;
wire n_4929;
wire n_2874;
wire n_4117;
wire n_3049;
wire n_3634;
wire n_5436;
wire n_2341;
wire n_1654;
wire n_3066;
wire n_2045;
wire n_3913;
wire n_5341;
wire n_2575;
wire n_3739;
wire n_1230;
wire n_5140;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_4541;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_5096;
wire n_2043;
wire n_4171;
wire n_4815;
wire n_4665;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_4276;
wire n_1378;
wire n_5268;
wire n_5050;
wire n_5240;
wire n_5503;
wire n_1461;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_1112;
wire n_700;
wire n_4174;
wire n_5131;
wire n_5546;
wire n_5174;
wire n_2145;
wire n_4801;
wire n_680;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_3119;
wire n_4740;
wire n_1108;
wire n_1274;
wire n_4394;
wire n_5544;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_5541;
wire n_916;
wire n_2810;
wire n_1884;
wire n_1555;
wire n_762;
wire n_1253;
wire n_1468;
wire n_4378;
wire n_5166;
wire n_2683;
wire n_4180;
wire n_4459;
wire n_3624;
wire n_1182;
wire n_4594;
wire n_2748;
wire n_4642;
wire n_1376;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_3544;
wire n_5300;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_5381;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_1083;
wire n_5333;
wire n_4914;
wire n_3510;
wire n_4587;
wire n_1139;
wire n_3688;
wire n_5008;
wire n_1312;
wire n_3871;
wire n_892;
wire n_3757;
wire n_1567;
wire n_2219;
wire n_2100;
wire n_3666;
wire n_5538;
wire n_990;
wire n_867;
wire n_3479;
wire n_944;
wire n_5499;
wire n_749;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_4285;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_650;
wire n_3741;
wire n_5582;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_5109;
wire n_712;
wire n_909;
wire n_1392;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_964;
wire n_2220;
wire n_4433;
wire n_2829;
wire n_1914;
wire n_2253;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_1633;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_2434;
wire n_1234;
wire n_3936;
wire n_5564;
wire n_2261;
wire n_3082;
wire n_5162;
wire n_5442;
wire n_2473;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_3867;
wire n_3397;
wire n_1646;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_1237;
wire n_1095;
wire n_3078;
wire n_3971;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_1531;
wire n_2113;
wire n_1387;
wire n_3711;
wire n_5054;
wire n_3171;
wire n_5394;
wire n_4751;
wire n_4242;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_1496;
wire n_2812;
wire n_3300;
wire n_5496;
wire n_3104;
wire n_4122;
wire n_2132;
wire n_4522;
wire n_4952;
wire n_4426;
wire n_4362;
wire n_3267;
wire n_3946;
wire n_2112;
wire n_2640;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_4089;
wire n_3513;
wire n_1173;
wire n_3498;
wire n_5132;
wire n_2350;
wire n_5535;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_4728;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_3863;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_3332;
wire n_2055;
wire n_2998;
wire n_1423;
wire n_4359;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_5176;
wire n_4039;
wire n_1798;
wire n_3057;
wire n_1608;
wire n_677;
wire n_3983;
wire n_703;
wire n_3318;
wire n_3385;
wire n_3773;
wire n_3494;
wire n_1278;
wire n_5074;
wire n_3788;
wire n_3939;
wire n_727;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_2496;
wire n_3260;
wire n_3349;
wire n_4348;
wire n_1602;
wire n_3139;
wire n_3801;
wire n_2338;
wire n_5261;
wire n_1080;
wire n_3636;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_2057;
wire n_1205;
wire n_2716;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_1120;
wire n_1202;
wire n_4084;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_2774;
wire n_2799;
wire n_4393;
wire n_3984;
wire n_1586;
wire n_1431;
wire n_4389;
wire n_1763;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_3737;
wire n_2379;
wire n_3579;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_5244;
wire n_5114;
wire n_4551;
wire n_4521;
wire n_2284;
wire n_3005;
wire n_5420;
wire n_2283;
wire n_5206;
wire n_2526;
wire n_1097;
wire n_1711;
wire n_4387;
wire n_2508;
wire n_3186;
wire n_2594;
wire n_1239;
wire n_5298;
wire n_3417;
wire n_890;
wire n_3626;
wire n_4598;
wire n_4464;
wire n_5106;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_1081;
wire n_2119;
wire n_2493;
wire n_5080;
wire n_4565;
wire n_3392;
wire n_1800;
wire n_5081;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_3512;
wire n_1734;
wire n_1860;
wire n_4552;
wire n_2840;
wire n_4482;
wire n_837;
wire n_812;
wire n_4172;
wire n_4040;
wire n_3024;
wire n_5567;
wire n_5406;
wire n_4328;
wire n_1854;
wire n_666;
wire n_5191;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2893;
wire n_4940;
wire n_785;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_4112;
wire n_2035;
wire n_4928;
wire n_2614;
wire n_5428;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_2128;
wire n_4071;
wire n_4436;
wire n_3586;
wire n_4160;
wire n_1668;
wire n_4137;
wire n_1078;
wire n_5417;
wire n_4545;
wire n_4758;
wire n_1161;
wire n_4840;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_1191;
wire n_4535;
wire n_4385;
wire n_1215;
wire n_3748;
wire n_4731;
wire n_2337;
wire n_1786;
wire n_3732;
wire n_1804;
wire n_4671;
wire n_2272;
wire n_5571;
wire n_4766;
wire n_4558;
wire n_1318;
wire n_1769;
wire n_1632;
wire n_1929;
wire n_4319;
wire n_2929;
wire n_4358;
wire n_1526;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_1997;
wire n_1137;
wire n_1258;
wire n_1733;
wire n_640;
wire n_4651;
wire n_943;
wire n_3167;
wire n_4748;
wire n_1807;
wire n_1123;
wire n_2857;
wire n_1784;
wire n_4618;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_752;
wire n_985;
wire n_5506;
wire n_5475;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_1352;
wire n_5431;
wire n_643;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1822;
wire n_1441;
wire n_682;
wire n_5315;
wire n_2633;
wire n_3708;
wire n_2907;
wire n_1429;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_686;
wire n_1154;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_3718;
wire n_756;
wire n_3390;
wire n_2298;
wire n_1016;
wire n_1149;
wire n_4666;
wire n_4082;
wire n_2320;
wire n_3140;
wire n_979;
wire n_3976;
wire n_2813;
wire n_897;
wire n_2546;
wire n_3381;
wire n_3736;
wire n_4466;
wire n_891;
wire n_885;
wire n_1659;
wire n_3955;
wire n_5366;
wire n_5322;
wire n_1864;
wire n_5414;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_3336;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_714;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_725;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_2198;
wire n_5369;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_1852;
wire n_801;
wire n_4377;
wire n_818;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5593;
wire n_5270;
wire n_3468;
wire n_1877;
wire n_4301;
wire n_5313;
wire n_2133;
wire n_2497;
wire n_879;
wire n_5446;
wire n_4561;
wire n_1541;
wire n_3291;
wire n_1472;
wire n_1050;
wire n_2578;
wire n_1201;
wire n_1185;
wire n_2475;
wire n_4715;
wire n_2715;
wire n_2665;
wire n_4879;
wire n_5044;
wire n_3755;
wire n_1090;
wire n_4536;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_5459;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_4418;
wire n_3341;
wire n_4125;
wire n_5390;
wire n_5351;
wire n_5267;
wire n_1116;
wire n_5024;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_4151;
wire n_2845;
wire n_4412;
wire n_2036;
wire n_843;
wire n_3358;
wire n_2003;
wire n_2533;
wire n_1307;
wire n_4682;
wire n_1128;
wire n_2419;
wire n_2330;
wire n_5078;
wire n_4810;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_1440;
wire n_1370;
wire n_5005;
wire n_1549;
wire n_5207;
wire n_2658;
wire n_3620;
wire n_4601;
wire n_1065;
wire n_4518;
wire n_2767;
wire n_5474;
wire n_3376;
wire n_1362;
wire n_3123;
wire n_5447;
wire n_2692;
wire n_683;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_2862;
wire n_4325;
wire n_1420;
wire n_2645;
wire n_2553;
wire n_4711;
wire n_2749;
wire n_660;
wire n_4413;
wire n_1210;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_1038;
wire n_3723;
wire n_4135;
wire n_5223;
wire n_3880;
wire n_3904;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_3405;
wire n_2313;
wire n_1022;
wire n_5465;
wire n_3532;
wire n_5154;
wire n_2609;
wire n_1767;
wire n_4138;
wire n_1040;
wire n_3131;
wire n_1973;
wire n_1444;
wire n_820;
wire n_2882;
wire n_2303;
wire n_4384;
wire n_4639;
wire n_1664;
wire n_4577;
wire n_2154;
wire n_1986;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_984;
wire n_5087;
wire n_1552;
wire n_2938;
wire n_2498;
wire n_3992;
wire n_1772;
wire n_1311;
wire n_3106;
wire n_2881;
wire n_3092;
wire n_4270;
wire n_697;
wire n_4620;
wire n_5397;
wire n_4924;
wire n_4044;
wire n_2305;
wire n_880;
wire n_5566;
wire n_3304;
wire n_4388;
wire n_3247;
wire n_739;
wire n_1028;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_2809;
wire n_975;
wire n_1645;
wire n_932;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_5492;
wire n_2465;
wire n_5501;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_3178;
wire n_2251;
wire n_3100;
wire n_3721;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_4973;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_2487;
wire n_5473;
wire n_1834;
wire n_1011;
wire n_2534;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_3576;
wire n_5562;
wire n_4858;
wire n_1445;
wire n_5370;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_2387;
wire n_4318;
wire n_5227;
wire n_830;
wire n_987;
wire n_2510;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_2639;
wire n_4738;
wire n_2603;
wire n_5386;
wire n_1167;
wire n_4554;
wire n_4526;
wire n_4105;
wire n_3663;
wire n_969;
wire n_1663;
wire n_2086;
wire n_1926;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3431;
wire n_3355;
wire n_1738;
wire n_3897;
wire n_1735;
wire n_4005;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_2597;
wire n_1077;
wire n_956;
wire n_765;
wire n_4092;
wire n_4875;
wire n_4255;
wire n_2758;
wire n_5036;
wire n_1271;
wire n_2186;
wire n_4647;
wire n_3575;
wire n_2471;
wire n_3042;
wire n_1067;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_900;
wire n_5485;
wire n_5525;
wire n_3004;
wire n_1551;
wire n_4849;
wire n_5271;
wire n_2039;
wire n_1285;
wire n_761;
wire n_733;
wire n_3838;
wire n_4059;
wire n_5194;
wire n_5445;
wire n_2734;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_2420;
wire n_648;
wire n_3273;
wire n_2918;
wire n_835;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_1792;
wire n_5245;
wire n_2062;
wire n_4489;
wire n_822;
wire n_1459;
wire n_2153;
wire n_5329;
wire n_5472;
wire n_839;
wire n_1754;
wire n_4833;
wire n_3394;
wire n_2235;
wire n_1575;
wire n_4564;
wire n_1848;
wire n_1172;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_5072;
wire n_3778;
wire n_4322;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_997;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_3001;
wire n_5260;
wire n_4981;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_5372;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_2422;
wire n_654;
wire n_2933;
wire n_3387;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_1059;
wire n_2736;
wire n_3825;
wire n_4198;
wire n_977;
wire n_2339;
wire n_2532;
wire n_4373;
wire n_1866;
wire n_2664;
wire n_4154;
wire n_4390;
wire n_1782;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_2360;
wire n_4453;
wire n_723;
wire n_1393;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3032;
wire n_4886;
wire n_5172;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1982;
wire n_641;
wire n_5311;
wire n_910;
wire n_5164;
wire n_4964;
wire n_4700;
wire n_4002;
wire n_1114;
wire n_1742;
wire n_4679;
wire n_3815;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_2982;
wire n_1273;
wire n_5495;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_5547;
wire n_4693;
wire n_1043;
wire n_5121;
wire n_4956;
wire n_2869;
wire n_5379;
wire n_4487;
wire n_2674;
wire n_1737;
wire n_1613;
wire n_3026;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_954;
wire n_3112;
wire n_2051;
wire n_3196;
wire n_2673;
wire n_4678;
wire n_664;
wire n_1591;
wire n_5301;
wire n_5126;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_3779;
wire n_1063;
wire n_991;
wire n_2275;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_938;
wire n_1891;
wire n_5348;
wire n_1000;
wire n_4868;
wire n_4072;
wire n_2792;
wire n_4465;
wire n_2596;
wire n_5217;
wire n_3986;
wire n_5558;
wire n_3725;
wire n_4026;
wire n_4245;
wire n_5520;
wire n_2524;
wire n_3894;
wire n_1702;
wire n_4852;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_1232;
wire n_1211;
wire n_996;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_866;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_1644;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_2255;
wire n_5554;
wire n_1252;
wire n_3045;
wire n_773;
wire n_5135;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_5448;
wire n_2573;
wire n_2336;
wire n_5412;
wire n_1662;
wire n_3249;
wire n_3483;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_782;
wire n_2915;
wire n_4869;
wire n_3213;
wire n_5533;
wire n_4047;
wire n_1244;
wire n_1796;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_1574;
wire n_3033;
wire n_893;
wire n_1582;
wire n_1981;
wire n_2824;
wire n_5327;
wire n_4417;
wire n_796;
wire n_1374;
wire n_2089;
wire n_4688;
wire n_4939;
wire n_1486;
wire n_3619;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_691;
wire n_4903;
wire n_2131;
wire n_3853;
wire n_4382;
wire n_2509;
wire n_4085;
wire n_5486;
wire n_2135;
wire n_4475;
wire n_5432;
wire n_1463;
wire n_4626;
wire n_4997;
wire n_5065;
wire n_924;
wire n_781;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_2436;
wire n_3517;
wire n_1706;
wire n_2461;
wire n_3719;
wire n_1214;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_5295;
wire n_1181;
wire n_1999;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_3383;
wire n_1835;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_4600;
wire n_1453;
wire n_3943;
wire n_3145;
wire n_2908;
wire n_4106;
wire n_2156;
wire n_1184;
wire n_754;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_1277;
wire n_1746;
wire n_1062;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_740;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_3283;
wire n_4331;
wire n_4159;
wire n_3451;
wire n_4734;
wire n_2832;
wire n_1688;
wire n_2370;
wire n_1944;
wire n_2914;
wire n_1988;
wire n_1718;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_2539;
wire n_5555;
wire n_2078;
wire n_1145;
wire n_4809;
wire n_787;
wire n_4012;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_1207;
wire n_3606;
wire n_2232;
wire n_1847;
wire n_4320;
wire n_5084;
wire n_5251;
wire n_1314;
wire n_1512;
wire n_884;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_5407;
wire n_2988;
wire n_4560;
wire n_3230;
wire n_3793;
wire n_859;
wire n_5042;
wire n_4768;
wire n_1889;
wire n_693;
wire n_5368;
wire n_929;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_3607;
wire n_1637;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_5310;
wire n_2769;
wire n_1548;
wire n_4987;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_2902;
wire n_4360;
wire n_1544;
wire n_4540;
wire n_2094;
wire n_5588;
wire n_3854;
wire n_1354;
wire n_2349;
wire n_3652;
wire n_3449;
wire n_1021;
wire n_3089;
wire n_4854;
wire n_1595;
wire n_1142;
wire n_5477;
wire n_2727;
wire n_942;
wire n_5234;
wire n_1416;
wire n_1599;
wire n_4747;
wire n_3472;
wire n_2527;
wire n_3126;
wire n_2759;
wire n_5007;
wire n_4881;
wire n_2038;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_2806;
wire n_4502;
wire n_3191;
wire n_1716;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_5253;
wire n_3588;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_5418;
wire n_5019;
wire n_1819;
wire n_3095;
wire n_947;
wire n_3698;
wire n_4513;
wire n_1179;
wire n_696;
wire n_1442;
wire n_4775;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_2499;
wire n_2549;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_3885;
wire n_955;
wire n_4264;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_3839;
wire n_5490;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_5489;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_4794;
wire n_4843;
wire n_669;
wire n_5580;
wire n_5215;
wire n_3937;
wire n_4763;
wire n_1418;
wire n_4170;
wire n_5561;
wire n_2462;
wire n_2155;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_3604;
wire n_5430;
wire n_824;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_3792;
wire n_4267;
wire n_2083;
wire n_815;
wire n_2753;
wire n_1340;
wire n_3021;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_2898;
wire n_1825;
wire n_3567;
wire n_2682;
wire n_5585;
wire n_5112;
wire n_5326;
wire n_1627;
wire n_2903;
wire n_5303;
wire n_3812;
wire n_3127;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_5530;
wire n_965;
wire n_934;
wire n_2213;
wire n_4056;
wire n_4806;
wire n_1674;
wire n_4015;
wire n_2924;
wire n_4445;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_1455;
wire n_2287;
wire n_836;
wire n_3415;
wire n_3464;
wire n_3414;
wire n_4234;
wire n_760;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_3467;
wire n_713;
wire n_3179;
wire n_5522;
wire n_4836;
wire n_3889;
wire n_5262;
wire n_3262;
wire n_5319;
wire n_927;
wire n_3699;
wire n_706;
wire n_2120;
wire n_1419;
wire n_3816;
wire n_3528;
wire n_4207;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_2312;
wire n_1826;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_5335;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_5284;
wire n_4978;
wire n_3246;
wire n_3299;
wire n_980;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_905;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_5516;
wire n_3615;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_3200;
wire n_3642;
wire n_2146;
wire n_4274;
wire n_5583;
wire n_3276;
wire n_5433;
wire n_3682;
wire n_5429;
wire n_4007;
wire n_1456;
wire n_1879;
wire n_2129;
wire n_814;
wire n_5120;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_1134;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_647;
wire n_2932;
wire n_2027;
wire n_3118;
wire n_5560;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_5455;
wire n_1467;
wire n_5209;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_5099;
wire n_681;
wire n_3286;
wire n_2023;
wire n_3974;
wire n_3443;
wire n_2599;
wire n_3988;
wire n_5022;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_1098;
wire n_3009;
wire n_777;
wire n_5219;
wire n_920;
wire n_3951;
wire n_5518;
wire n_3035;
wire n_4261;
wire n_1132;
wire n_1823;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_861;
wire n_1666;
wire n_5103;
wire n_4648;
wire n_2214;
wire n_2256;
wire n_3326;
wire n_2732;
wire n_1883;
wire n_4094;
wire n_2776;
wire n_3224;
wire n_1969;
wire n_2949;
wire n_4269;
wire n_1927;
wire n_1222;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_2449;
wire n_4428;
wire n_745;
wire n_1572;
wire n_4463;
wire n_5357;
wire n_3648;
wire n_1975;
wire n_5421;
wire n_1388;
wire n_1266;
wire n_4396;
wire n_1990;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1075;
wire n_1890;
wire n_4034;
wire n_4228;
wire n_1227;
wire n_3166;
wire n_3649;
wire n_3065;
wire n_5045;
wire n_5237;
wire n_657;
wire n_3924;
wire n_3997;
wire n_3564;
wire n_862;
wire n_2637;
wire n_3795;
wire n_4931;
wire n_2306;
wire n_2071;
wire n_3953;
wire n_4400;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_5434;
wire n_1532;
wire n_1030;
wire n_5181;
wire n_3208;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_852;
wire n_2916;
wire n_1060;
wire n_4424;
wire n_4351;
wire n_4192;
wire n_1748;
wire n_1301;
wire n_3400;
wire n_1466;
wire n_2581;
wire n_1783;
wire n_5146;
wire n_4646;
wire n_4221;
wire n_1037;
wire n_3650;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_4035;
wire n_1480;
wire n_3670;
wire n_2540;
wire n_4190;
wire n_1605;
wire n_3060;
wire n_2984;
wire n_4009;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_5577;
wire n_876;
wire n_5017;
wire n_736;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_4717;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_854;
wire n_2091;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_1658;
wire n_1072;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_2725;
wire n_2667;
wire n_3746;
wire n_4537;
wire n_1046;
wire n_3694;
wire n_771;
wire n_5456;
wire n_3893;
wire n_4847;
wire n_2307;
wire n_3702;
wire n_1984;
wire n_3453;
wire n_1556;
wire n_5345;
wire n_2815;
wire n_4427;
wire n_1824;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_819;
wire n_1971;
wire n_2945;
wire n_3543;
wire n_1324;
wire n_1776;
wire n_3448;
wire n_4279;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_4152;
wire n_5537;
wire n_2698;
wire n_5572;
wire n_4783;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_5409;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_807;
wire n_5142;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_802;
wire n_5401;
wire n_4595;
wire n_960;
wire n_2352;
wire n_5201;
wire n_790;
wire n_5551;
wire n_5416;
wire n_4404;
wire n_2377;
wire n_2652;
wire n_5498;
wire n_5543;
wire n_4054;
wire n_1286;
wire n_4617;
wire n_1685;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_1052;
wire n_4732;
wire n_2076;
wire n_2203;
wire n_1426;
wire n_4969;
wire n_5252;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_4140;
wire n_5171;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_3309;
wire n_2796;
wire n_858;
wire n_5393;
wire n_4817;
wire n_2136;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_2771;
wire n_2403;
wire n_2947;
wire n_928;
wire n_3769;
wire n_1565;
wire n_4437;
wire n_3055;
wire n_4070;
wire n_5346;
wire n_748;
wire n_1045;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_4139;
wire n_4769;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_2713;
wire n_1422;
wire n_1965;
wire n_644;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_2934;
wire n_5104;
wire n_2210;
wire n_4368;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_1049;
wire n_4430;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_1356;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_5578;
wire n_728;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_3255;
wire n_2588;
wire n_935;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_911;
wire n_3509;
wire n_1403;
wire n_5395;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_3456;
wire n_4532;
wire n_3790;
wire n_907;
wire n_847;
wire n_747;
wire n_1135;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_5199;
wire n_4257;
wire n_4282;
wire n_4341;
wire n_1694;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_5480;
wire n_3077;
wire n_4944;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_3533;
wire n_5175;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_3583;
wire n_4316;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_1157;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_1789;
wire n_763;
wire n_2174;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_4703;
wire n_1687;
wire n_4934;
wire n_2638;
wire n_2046;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_1587;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_1427;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_4669;
wire n_5228;
wire n_1100;
wire n_1617;
wire n_2600;
wire n_3436;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_1175;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_1621;
wire n_5186;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_3664;
wire n_4218;
wire n_4687;
wire n_1381;
wire n_3686;
wire n_1183;
wire n_4720;
wire n_2889;
wire n_2141;
wire n_1758;
wire n_1110;
wire n_3470;
wire n_5221;
wire n_1407;
wire n_2865;
wire n_973;
wire n_5591;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_1176;
wire n_3677;
wire n_1054;
wire n_5387;
wire n_3292;
wire n_3989;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_1057;
wire n_4131;
wire n_5449;
wire n_4215;
wire n_978;
wire n_2488;
wire n_1509;
wire n_828;
wire n_4158;
wire n_3079;
wire n_5190;
wire n_3269;
wire n_5325;
wire n_4231;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_653;
wire n_4926;
wire n_2050;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5344;
wire n_2550;
wire n_1536;
wire n_3177;
wire n_4667;
wire n_1471;
wire n_3440;
wire n_3658;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_788;
wire n_2169;
wire n_5133;
wire n_5305;
wire n_2175;
wire n_1625;
wire n_4578;
wire n_3644;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_1922;
wire n_940;
wire n_1537;
wire n_4877;
wire n_2065;
wire n_4470;
wire n_4187;
wire n_1904;
wire n_4998;
wire n_5576;
wire n_2395;
wire n_2868;
wire n_1530;
wire n_4057;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_898;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_5343;
wire n_1093;
wire n_4021;
wire n_3379;
wire n_4379;
wire n_2268;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_668;
wire n_2111;
wire n_3743;
wire n_5542;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_5527;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_2583;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_701;
wire n_1003;
wire n_4472;
wire n_2699;
wire n_3901;
wire n_5180;
wire n_1640;
wire n_2973;
wire n_2710;
wire n_2505;
wire n_4519;
wire n_5025;
wire n_2397;
wire n_3878;
wire n_4197;
wire n_2721;
wire n_1892;
wire n_2615;
wire n_4787;
wire n_1212;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_4371;
wire n_1902;
wire n_2784;
wire n_3898;
wire n_694;
wire n_4749;
wire n_1845;
wire n_921;
wire n_5545;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_5083;
wire n_3253;
wire n_2088;
wire n_1275;
wire n_4238;
wire n_904;
wire n_2005;
wire n_1696;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_3846;
wire n_5122;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_3845;
wire n_3203;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_950;
wire n_711;
wire n_4168;
wire n_1369;
wire n_4298;
wire n_4743;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_3690;
wire n_3229;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_4211;
wire n_3094;
wire n_741;
wire n_5185;
wire n_2964;
wire n_5032;
wire n_865;
wire n_5034;
wire n_3312;
wire n_1041;
wire n_2451;
wire n_2913;
wire n_993;
wire n_1862;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_2839;
wire n_3237;
wire n_4128;
wire n_4036;
wire n_5269;
wire n_3655;
wire n_2955;
wire n_1764;
wire n_4807;
wire n_5115;
wire n_902;
wire n_1723;
wire n_3918;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_4095;
wire n_1310;
wire n_4485;
wire n_3593;
wire n_5163;
wire n_1229;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_1516;
wire n_4890;
wire n_2485;
wire n_4224;
wire n_2563;
wire n_1670;
wire n_1799;
wire n_5507;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_3519;
wire n_2209;
wire n_4042;
wire n_4244;
wire n_1928;
wire n_4708;
wire n_4883;
wire n_4553;
wire n_1634;
wire n_1203;
wire n_1699;
wire n_5226;
wire n_2081;
wire n_1474;
wire n_937;
wire n_1631;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_3772;
wire n_2891;
wire n_4335;
wire n_3128;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_4516;
wire n_5235;
wire n_1129;
wire n_1464;
wire n_2798;
wire n_3217;
wire n_1249;
wire n_3821;
wire n_3201;
wire n_3503;
wire n_1870;
wire n_4467;
wire n_5521;
wire n_2654;
wire n_3935;
wire n_1861;
wire n_1228;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_5410;
wire n_1251;
wire n_1989;
wire n_2689;
wire n_1762;
wire n_3798;
wire n_3080;
wire n_5241;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_3308;
wire n_841;
wire n_3204;
wire n_4134;
wire n_5018;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_5258;

INVx1_ASAP7_75t_L g639 ( 
.A(n_83),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_370),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_452),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_204),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_439),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_472),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_459),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_470),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_483),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_504),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_243),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_617),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_514),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_28),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_364),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_131),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_339),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_619),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_361),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_53),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_276),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_441),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_592),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_399),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_174),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_226),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_544),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_138),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_104),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_46),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_346),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_153),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_261),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_116),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_102),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_219),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_373),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_207),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_126),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_102),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_429),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_43),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_125),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_202),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_380),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_529),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_125),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_558),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_262),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_163),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_73),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_611),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_289),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_218),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_113),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_259),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_285),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_308),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_632),
.Y(n_697)
);

CKINVDCx16_ASAP7_75t_R g698 ( 
.A(n_410),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_599),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_79),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_328),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_457),
.Y(n_702)
);

INVx1_ASAP7_75t_SL g703 ( 
.A(n_566),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_547),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_167),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_87),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_635),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_437),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_474),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_47),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_466),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_8),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_229),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_129),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_76),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_7),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_143),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_638),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_614),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_43),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_397),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_98),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_625),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_268),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_507),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_566),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_34),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_65),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_608),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_17),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_302),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_75),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_479),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_202),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_177),
.Y(n_735)
);

BUFx2_ASAP7_75t_SL g736 ( 
.A(n_109),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_348),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_105),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_309),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_352),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_170),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_307),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_399),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_459),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_55),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_242),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_517),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_447),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_368),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_178),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_215),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_542),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_101),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_373),
.Y(n_754)
);

CKINVDCx16_ASAP7_75t_R g755 ( 
.A(n_12),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_155),
.Y(n_756)
);

BUFx2_ASAP7_75t_SL g757 ( 
.A(n_179),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_47),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_522),
.Y(n_759)
);

CKINVDCx16_ASAP7_75t_R g760 ( 
.A(n_65),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_119),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_11),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_629),
.Y(n_763)
);

INVxp67_ASAP7_75t_L g764 ( 
.A(n_340),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_448),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_156),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_173),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_491),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_484),
.Y(n_769)
);

BUFx10_ASAP7_75t_L g770 ( 
.A(n_605),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_405),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_404),
.Y(n_772)
);

BUFx10_ASAP7_75t_L g773 ( 
.A(n_419),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_93),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_284),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_437),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_5),
.Y(n_777)
);

INVxp67_ASAP7_75t_L g778 ( 
.A(n_213),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_297),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_334),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_343),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_347),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_276),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_626),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_72),
.Y(n_785)
);

BUFx10_ASAP7_75t_L g786 ( 
.A(n_474),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_48),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_231),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_572),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_70),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_83),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_562),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_579),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_360),
.Y(n_794)
);

BUFx10_ASAP7_75t_L g795 ( 
.A(n_201),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_434),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_8),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_57),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_86),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_136),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_303),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_607),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_114),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_455),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_475),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_241),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_367),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_561),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_185),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_613),
.Y(n_810)
);

CKINVDCx20_ASAP7_75t_R g811 ( 
.A(n_624),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_621),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_463),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_40),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_196),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_486),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_630),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_366),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_23),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_575),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_633),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_323),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_319),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_522),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_163),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_304),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_282),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_366),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_557),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_71),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_159),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_434),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_599),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_616),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_71),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_488),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_177),
.Y(n_837)
);

CKINVDCx20_ASAP7_75t_R g838 ( 
.A(n_486),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_631),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_441),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_327),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_24),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_279),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_588),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_248),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_407),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_531),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_467),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_349),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_424),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_596),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_112),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_364),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_196),
.Y(n_854)
);

BUFx10_ASAP7_75t_L g855 ( 
.A(n_610),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_547),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_406),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_497),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_147),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_224),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_111),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_279),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_417),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_557),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_413),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_495),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_444),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_454),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_534),
.Y(n_869)
);

INVx1_ASAP7_75t_SL g870 ( 
.A(n_451),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_200),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_585),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_517),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_420),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_358),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_130),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_275),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_620),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_269),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_259),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_546),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_233),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_33),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_374),
.Y(n_884)
);

INVx2_ASAP7_75t_SL g885 ( 
.A(n_25),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_277),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_380),
.Y(n_887)
);

HB1xp67_ASAP7_75t_L g888 ( 
.A(n_19),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_154),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_244),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_81),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_487),
.Y(n_892)
);

BUFx8_ASAP7_75t_SL g893 ( 
.A(n_450),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_395),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_456),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_138),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_571),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_280),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_447),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_487),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_257),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_148),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_44),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_307),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_321),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_455),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_290),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_421),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_295),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_141),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_356),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_75),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_606),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_545),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_273),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_300),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_171),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_210),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_96),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_530),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_540),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_56),
.Y(n_922)
);

CKINVDCx20_ASAP7_75t_R g923 ( 
.A(n_101),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_355),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_280),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_503),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_591),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_618),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_593),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_386),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_458),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_87),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_450),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_448),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_238),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_402),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_312),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_458),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_107),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_590),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_178),
.Y(n_941)
);

CKINVDCx20_ASAP7_75t_R g942 ( 
.A(n_520),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_179),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_263),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_272),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_483),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_147),
.Y(n_947)
);

CKINVDCx20_ASAP7_75t_R g948 ( 
.A(n_149),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_505),
.Y(n_949)
);

CKINVDCx20_ASAP7_75t_R g950 ( 
.A(n_254),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_258),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_343),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_242),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_347),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_415),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_221),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_318),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_117),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_21),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_174),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_505),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_85),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_113),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_7),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_24),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_159),
.Y(n_966)
);

BUFx10_ASAP7_75t_L g967 ( 
.A(n_285),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_634),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_444),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_593),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_528),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_79),
.Y(n_972)
);

INVx1_ASAP7_75t_SL g973 ( 
.A(n_368),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_78),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_344),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_64),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_130),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_19),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_90),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_585),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_607),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_493),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_628),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_234),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_235),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_144),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_122),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_575),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_636),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_267),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_17),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_622),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_358),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_6),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_5),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_195),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_235),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_497),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_435),
.Y(n_999)
);

CKINVDCx20_ASAP7_75t_R g1000 ( 
.A(n_243),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_605),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_39),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_524),
.Y(n_1003)
);

CKINVDCx14_ASAP7_75t_R g1004 ( 
.A(n_218),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_155),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_176),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_319),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_496),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_435),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_414),
.Y(n_1010)
);

CKINVDCx14_ASAP7_75t_R g1011 ( 
.A(n_99),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_528),
.Y(n_1012)
);

CKINVDCx16_ASAP7_75t_R g1013 ( 
.A(n_340),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_233),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_186),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_145),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_623),
.Y(n_1017)
);

CKINVDCx20_ASAP7_75t_R g1018 ( 
.A(n_109),
.Y(n_1018)
);

BUFx2_ASAP7_75t_L g1019 ( 
.A(n_57),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_390),
.Y(n_1020)
);

BUFx10_ASAP7_75t_L g1021 ( 
.A(n_386),
.Y(n_1021)
);

CKINVDCx20_ASAP7_75t_R g1022 ( 
.A(n_85),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_171),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_562),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_609),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_239),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_197),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_70),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_440),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_466),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_21),
.Y(n_1031)
);

INVxp67_ASAP7_75t_L g1032 ( 
.A(n_349),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_568),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_80),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_342),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_273),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_637),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_417),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_597),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_114),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_304),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_475),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_510),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_627),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_195),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_583),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_211),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_416),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_146),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_303),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_149),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_1),
.Y(n_1052)
);

BUFx10_ASAP7_75t_L g1053 ( 
.A(n_206),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_219),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_305),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_61),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_470),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_49),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_77),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_44),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_188),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_245),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_189),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_537),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_212),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_140),
.Y(n_1066)
);

CKINVDCx16_ASAP7_75t_R g1067 ( 
.A(n_28),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_3),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_272),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_594),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_53),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_299),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_524),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_553),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_338),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_293),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_148),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_248),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_540),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_40),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_390),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_230),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_520),
.Y(n_1083)
);

BUFx8_ASAP7_75t_SL g1084 ( 
.A(n_507),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_384),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_67),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_365),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_451),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_414),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_561),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_266),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_344),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_560),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_275),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_313),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_271),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_491),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_117),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_529),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_568),
.Y(n_1100)
);

CKINVDCx14_ASAP7_75t_R g1101 ( 
.A(n_442),
.Y(n_1101)
);

CKINVDCx14_ASAP7_75t_R g1102 ( 
.A(n_481),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_288),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_161),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_510),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_612),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_333),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_615),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_595),
.Y(n_1109)
);

BUFx10_ASAP7_75t_L g1110 ( 
.A(n_477),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_385),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_73),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_598),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_99),
.Y(n_1114)
);

INVx1_ASAP7_75t_SL g1115 ( 
.A(n_543),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_577),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_66),
.Y(n_1117)
);

BUFx10_ASAP7_75t_L g1118 ( 
.A(n_370),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_337),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_387),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_74),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_374),
.Y(n_1122)
);

INVx1_ASAP7_75t_SL g1123 ( 
.A(n_452),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_388),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_467),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_539),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_119),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_189),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_351),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_124),
.Y(n_1130)
);

CKINVDCx20_ASAP7_75t_R g1131 ( 
.A(n_121),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_604),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_564),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_92),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_197),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_934),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_934),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_934),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_934),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1004),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_713),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_1011),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_713),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_784),
.B(n_1),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_713),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_750),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_1101),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_784),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_656),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_750),
.Y(n_1150)
);

INVx1_ASAP7_75t_SL g1151 ( 
.A(n_893),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_750),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_823),
.Y(n_1153)
);

CKINVDCx20_ASAP7_75t_R g1154 ( 
.A(n_698),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_738),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_823),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_823),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_1102),
.Y(n_1158)
);

INVxp67_ASAP7_75t_SL g1159 ( 
.A(n_836),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_836),
.Y(n_1160)
);

NOR2xp67_ASAP7_75t_L g1161 ( 
.A(n_687),
.B(n_0),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_836),
.Y(n_1162)
);

CKINVDCx20_ASAP7_75t_R g1163 ( 
.A(n_698),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_1084),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_689),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_966),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_966),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_667),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_855),
.Y(n_1169)
);

INVxp67_ASAP7_75t_L g1170 ( 
.A(n_738),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_966),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1026),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1026),
.Y(n_1173)
);

CKINVDCx16_ASAP7_75t_R g1174 ( 
.A(n_755),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_689),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1026),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1074),
.Y(n_1177)
);

CKINVDCx14_ASAP7_75t_R g1178 ( 
.A(n_855),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1074),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_855),
.Y(n_1180)
);

CKINVDCx16_ASAP7_75t_R g1181 ( 
.A(n_755),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1074),
.Y(n_1182)
);

INVxp67_ASAP7_75t_SL g1183 ( 
.A(n_646),
.Y(n_1183)
);

BUFx2_ASAP7_75t_SL g1184 ( 
.A(n_855),
.Y(n_1184)
);

INVxp33_ASAP7_75t_SL g1185 ( 
.A(n_654),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_687),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_687),
.Y(n_1187)
);

INVxp67_ASAP7_75t_L g1188 ( 
.A(n_753),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_650),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_904),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_760),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_904),
.Y(n_1192)
);

NOR2xp67_ASAP7_75t_L g1193 ( 
.A(n_904),
.B(n_0),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_646),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_646),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_664),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_664),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_664),
.Y(n_1198)
);

INVxp33_ASAP7_75t_SL g1199 ( 
.A(n_801),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_686),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_686),
.Y(n_1201)
);

CKINVDCx20_ASAP7_75t_R g1202 ( 
.A(n_760),
.Y(n_1202)
);

CKINVDCx14_ASAP7_75t_R g1203 ( 
.A(n_729),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_689),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_686),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_710),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_710),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_1013),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_710),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_775),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_1013),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1067),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_689),
.Y(n_1213)
);

CKINVDCx20_ASAP7_75t_R g1214 ( 
.A(n_1067),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_775),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_770),
.B(n_2),
.Y(n_1216)
);

INVxp33_ASAP7_75t_SL g1217 ( 
.A(n_888),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_811),
.Y(n_1218)
);

INVxp67_ASAP7_75t_L g1219 ( 
.A(n_753),
.Y(n_1219)
);

INVx1_ASAP7_75t_SL g1220 ( 
.A(n_670),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_775),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_689),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_674),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_689),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_782),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_782),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_782),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_807),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_807),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_807),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_799),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_869),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_640),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_869),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_869),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_908),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_650),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_908),
.Y(n_1238)
);

INVxp67_ASAP7_75t_SL g1239 ( 
.A(n_908),
.Y(n_1239)
);

CKINVDCx16_ASAP7_75t_R g1240 ( 
.A(n_770),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_642),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_912),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_912),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_690),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_643),
.Y(n_1245)
);

INVxp67_ASAP7_75t_SL g1246 ( 
.A(n_912),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_690),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_718),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_718),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_817),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_940),
.Y(n_1251)
);

INVxp33_ASAP7_75t_L g1252 ( 
.A(n_1012),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_799),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_644),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_649),
.Y(n_1255)
);

INVxp33_ASAP7_75t_L g1256 ( 
.A(n_835),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_835),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_656),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_940),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_693),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_940),
.Y(n_1261)
);

CKINVDCx20_ASAP7_75t_R g1262 ( 
.A(n_732),
.Y(n_1262)
);

INVxp67_ASAP7_75t_L g1263 ( 
.A(n_993),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_971),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_971),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_779),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_779),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_652),
.Y(n_1268)
);

INVxp67_ASAP7_75t_SL g1269 ( 
.A(n_971),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_756),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_653),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_984),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_984),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_984),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_650),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_998),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_998),
.Y(n_1277)
);

BUFx10_ASAP7_75t_L g1278 ( 
.A(n_928),
.Y(n_1278)
);

INVxp67_ASAP7_75t_L g1279 ( 
.A(n_993),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_998),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1027),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_657),
.Y(n_1282)
);

CKINVDCx16_ASAP7_75t_R g1283 ( 
.A(n_770),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1027),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_779),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1027),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_658),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1066),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1066),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1066),
.Y(n_1290)
);

INVxp33_ASAP7_75t_L g1291 ( 
.A(n_1019),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1075),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1075),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1075),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1078),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_659),
.Y(n_1296)
);

CKINVDCx20_ASAP7_75t_R g1297 ( 
.A(n_761),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1019),
.Y(n_1298)
);

INVxp67_ASAP7_75t_SL g1299 ( 
.A(n_1078),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1033),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1078),
.Y(n_1301)
);

INVxp67_ASAP7_75t_SL g1302 ( 
.A(n_1092),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_779),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_656),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1092),
.Y(n_1305)
);

INVxp67_ASAP7_75t_L g1306 ( 
.A(n_1033),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1092),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1120),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1120),
.Y(n_1309)
);

CKINVDCx16_ASAP7_75t_R g1310 ( 
.A(n_770),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_661),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_639),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_639),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_641),
.Y(n_1314)
);

CKINVDCx20_ASAP7_75t_R g1315 ( 
.A(n_804),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_641),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_645),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_645),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_647),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_647),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_779),
.Y(n_1321)
);

CKINVDCx20_ASAP7_75t_R g1322 ( 
.A(n_824),
.Y(n_1322)
);

NOR2xp67_ASAP7_75t_L g1323 ( 
.A(n_660),
.B(n_2),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_648),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_648),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_833),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_651),
.Y(n_1327)
);

CKINVDCx20_ASAP7_75t_R g1328 ( 
.A(n_838),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_651),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_662),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_655),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_655),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_665),
.Y(n_1333)
);

CKINVDCx16_ASAP7_75t_R g1334 ( 
.A(n_773),
.Y(n_1334)
);

BUFx2_ASAP7_75t_L g1335 ( 
.A(n_660),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_665),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_663),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_666),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_666),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_668),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_669),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_668),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_673),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_656),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_673),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_675),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_675),
.Y(n_1347)
);

INVxp33_ASAP7_75t_SL g1348 ( 
.A(n_671),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_677),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_779),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_672),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_677),
.Y(n_1352)
);

INVxp33_ASAP7_75t_L g1353 ( 
.A(n_678),
.Y(n_1353)
);

INVxp67_ASAP7_75t_L g1354 ( 
.A(n_736),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_792),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_678),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_676),
.Y(n_1357)
);

INVxp67_ASAP7_75t_SL g1358 ( 
.A(n_792),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_679),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_680),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_681),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_682),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_679),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_684),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_853),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_684),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_694),
.Y(n_1367)
);

CKINVDCx20_ASAP7_75t_R g1368 ( 
.A(n_874),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_694),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_705),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_705),
.Y(n_1371)
);

CKINVDCx20_ASAP7_75t_R g1372 ( 
.A(n_889),
.Y(n_1372)
);

INVx4_ASAP7_75t_R g1373 ( 
.A(n_812),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_706),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_706),
.Y(n_1375)
);

INVxp33_ASAP7_75t_SL g1376 ( 
.A(n_683),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_714),
.Y(n_1377)
);

NOR2xp67_ASAP7_75t_L g1378 ( 
.A(n_780),
.B(n_885),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_685),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_714),
.Y(n_1380)
);

CKINVDCx14_ASAP7_75t_R g1381 ( 
.A(n_773),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_688),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_715),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_715),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_792),
.Y(n_1385)
);

INVxp33_ASAP7_75t_L g1386 ( 
.A(n_716),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_716),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_727),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_727),
.Y(n_1389)
);

CKINVDCx20_ASAP7_75t_R g1390 ( 
.A(n_897),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_688),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_733),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_656),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_733),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_742),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_742),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_745),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_745),
.Y(n_1398)
);

INVxp33_ASAP7_75t_SL g1399 ( 
.A(n_691),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_746),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_764),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_792),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_923),
.Y(n_1403)
);

INVxp67_ASAP7_75t_SL g1404 ( 
.A(n_792),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_780),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_746),
.Y(n_1406)
);

CKINVDCx20_ASAP7_75t_R g1407 ( 
.A(n_942),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_752),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_792),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_752),
.Y(n_1410)
);

INVxp67_ASAP7_75t_SL g1411 ( 
.A(n_949),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_762),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_762),
.Y(n_1413)
);

CKINVDCx20_ASAP7_75t_R g1414 ( 
.A(n_948),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_764),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_692),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_767),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_767),
.Y(n_1418)
);

INVx2_ASAP7_75t_SL g1419 ( 
.A(n_773),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_771),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_695),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_696),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_771),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_785),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_785),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_788),
.Y(n_1426)
);

CKINVDCx20_ASAP7_75t_R g1427 ( 
.A(n_950),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_778),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_788),
.Y(n_1429)
);

CKINVDCx16_ASAP7_75t_R g1430 ( 
.A(n_773),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_791),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_949),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_949),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_949),
.Y(n_1434)
);

INVxp33_ASAP7_75t_SL g1435 ( 
.A(n_699),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_949),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_700),
.Y(n_1437)
);

CKINVDCx14_ASAP7_75t_R g1438 ( 
.A(n_786),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_885),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_791),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_794),
.Y(n_1441)
);

INVx1_ASAP7_75t_SL g1442 ( 
.A(n_1000),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_949),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_794),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_797),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_797),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_800),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_977),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_800),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_802),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_1014),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_701),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_702),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_802),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_814),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_814),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_1018),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_815),
.Y(n_1458)
);

INVxp67_ASAP7_75t_SL g1459 ( 
.A(n_977),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_778),
.Y(n_1460)
);

INVxp67_ASAP7_75t_L g1461 ( 
.A(n_736),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_815),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_825),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_704),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_708),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_977),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_825),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_826),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_656),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_826),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_831),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_709),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_831),
.Y(n_1473)
);

CKINVDCx16_ASAP7_75t_R g1474 ( 
.A(n_786),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_832),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_711),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_712),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_977),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_977),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_977),
.Y(n_1480)
);

CKINVDCx16_ASAP7_75t_R g1481 ( 
.A(n_786),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_832),
.Y(n_1482)
);

INVxp67_ASAP7_75t_L g1483 ( 
.A(n_757),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1060),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_837),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_717),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_837),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_845),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_845),
.Y(n_1489)
);

BUFx6f_ASAP7_75t_L g1490 ( 
.A(n_1060),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_720),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_721),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_851),
.Y(n_1493)
);

INVxp33_ASAP7_75t_SL g1494 ( 
.A(n_722),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_724),
.Y(n_1495)
);

INVxp33_ASAP7_75t_L g1496 ( 
.A(n_851),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_858),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1036),
.Y(n_1498)
);

INVxp67_ASAP7_75t_L g1499 ( 
.A(n_757),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_725),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_858),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_726),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_728),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_860),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_860),
.Y(n_1505)
);

INVxp67_ASAP7_75t_L g1506 ( 
.A(n_866),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_866),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_868),
.Y(n_1508)
);

INVxp33_ASAP7_75t_SL g1509 ( 
.A(n_731),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1060),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_868),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_875),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_875),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_877),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_877),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_882),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_734),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_735),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_882),
.Y(n_1519)
);

BUFx10_ASAP7_75t_L g1520 ( 
.A(n_1060),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_891),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1060),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1032),
.Y(n_1523)
);

INVxp33_ASAP7_75t_SL g1524 ( 
.A(n_737),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1060),
.Y(n_1525)
);

CKINVDCx20_ASAP7_75t_R g1526 ( 
.A(n_1022),
.Y(n_1526)
);

CKINVDCx14_ASAP7_75t_R g1527 ( 
.A(n_786),
.Y(n_1527)
);

CKINVDCx20_ASAP7_75t_R g1528 ( 
.A(n_1065),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_891),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_892),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_892),
.Y(n_1531)
);

CKINVDCx20_ASAP7_75t_R g1532 ( 
.A(n_1131),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_895),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1032),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_895),
.Y(n_1535)
);

INVxp67_ASAP7_75t_L g1536 ( 
.A(n_896),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_896),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_902),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_902),
.Y(n_1539)
);

BUFx6f_ASAP7_75t_L g1540 ( 
.A(n_1109),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_913),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_913),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_915),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_915),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_916),
.Y(n_1545)
);

CKINVDCx14_ASAP7_75t_R g1546 ( 
.A(n_795),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_916),
.Y(n_1547)
);

INVxp33_ASAP7_75t_SL g1548 ( 
.A(n_739),
.Y(n_1548)
);

INVxp67_ASAP7_75t_L g1549 ( 
.A(n_918),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_918),
.Y(n_1550)
);

CKINVDCx20_ASAP7_75t_R g1551 ( 
.A(n_795),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1109),
.Y(n_1552)
);

CKINVDCx20_ASAP7_75t_R g1553 ( 
.A(n_795),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_920),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_740),
.Y(n_1555)
);

INVxp67_ASAP7_75t_SL g1556 ( 
.A(n_1109),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_920),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_922),
.Y(n_1558)
);

INVxp67_ASAP7_75t_SL g1559 ( 
.A(n_1109),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_817),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_922),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1137),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1218),
.Y(n_1563)
);

CKINVDCx20_ASAP7_75t_R g1564 ( 
.A(n_1223),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1138),
.Y(n_1565)
);

CKINVDCx20_ASAP7_75t_R g1566 ( 
.A(n_1223),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1165),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1184),
.B(n_821),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1139),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1183),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_L g1571 ( 
.A(n_1480),
.Y(n_1571)
);

CKINVDCx20_ASAP7_75t_R g1572 ( 
.A(n_1260),
.Y(n_1572)
);

CKINVDCx20_ASAP7_75t_R g1573 ( 
.A(n_1260),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1174),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1181),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1520),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1178),
.B(n_821),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_1218),
.Y(n_1578)
);

CKINVDCx20_ASAP7_75t_R g1579 ( 
.A(n_1262),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1239),
.Y(n_1580)
);

INVxp67_ASAP7_75t_L g1581 ( 
.A(n_1184),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1246),
.Y(n_1582)
);

INVxp67_ASAP7_75t_L g1583 ( 
.A(n_1168),
.Y(n_1583)
);

INVxp67_ASAP7_75t_L g1584 ( 
.A(n_1220),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_1203),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1269),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1299),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1208),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1302),
.Y(n_1589)
);

CKINVDCx20_ASAP7_75t_R g1590 ( 
.A(n_1262),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1136),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1136),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1186),
.Y(n_1593)
);

INVxp67_ASAP7_75t_SL g1594 ( 
.A(n_1189),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1164),
.Y(n_1595)
);

INVxp67_ASAP7_75t_SL g1596 ( 
.A(n_1189),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1164),
.Y(n_1597)
);

CKINVDCx20_ASAP7_75t_R g1598 ( 
.A(n_1270),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1442),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1159),
.B(n_834),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_1381),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1208),
.Y(n_1602)
);

INVxp67_ASAP7_75t_SL g1603 ( 
.A(n_1237),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_1438),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1169),
.B(n_834),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_1527),
.Y(n_1606)
);

CKINVDCx20_ASAP7_75t_R g1607 ( 
.A(n_1270),
.Y(n_1607)
);

CKINVDCx16_ASAP7_75t_R g1608 ( 
.A(n_1240),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1546),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1237),
.B(n_839),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1187),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1169),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_1180),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1211),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_1180),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1211),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1140),
.Y(n_1617)
);

INVxp67_ASAP7_75t_L g1618 ( 
.A(n_1382),
.Y(n_1618)
);

INVxp67_ASAP7_75t_L g1619 ( 
.A(n_1391),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1140),
.Y(n_1620)
);

CKINVDCx16_ASAP7_75t_R g1621 ( 
.A(n_1283),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1190),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1192),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1275),
.B(n_839),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1275),
.B(n_983),
.Y(n_1625)
);

CKINVDCx20_ASAP7_75t_R g1626 ( 
.A(n_1297),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1141),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_1142),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1143),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1142),
.B(n_983),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1145),
.Y(n_1631)
);

CKINVDCx20_ASAP7_75t_R g1632 ( 
.A(n_1297),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_1147),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1146),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1150),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1152),
.Y(n_1636)
);

CKINVDCx20_ASAP7_75t_R g1637 ( 
.A(n_1315),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1147),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1165),
.Y(n_1639)
);

CKINVDCx20_ASAP7_75t_R g1640 ( 
.A(n_1315),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_1233),
.Y(n_1641)
);

CKINVDCx20_ASAP7_75t_R g1642 ( 
.A(n_1322),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1233),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1256),
.B(n_1291),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1212),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1153),
.Y(n_1646)
);

INVxp33_ASAP7_75t_L g1647 ( 
.A(n_1252),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1241),
.Y(n_1648)
);

INVxp67_ASAP7_75t_SL g1649 ( 
.A(n_1358),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1156),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1157),
.Y(n_1651)
);

BUFx2_ASAP7_75t_L g1652 ( 
.A(n_1212),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1241),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_1245),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_1245),
.Y(n_1655)
);

BUFx6f_ASAP7_75t_L g1656 ( 
.A(n_1480),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1160),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1162),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1166),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1167),
.Y(n_1660)
);

CKINVDCx20_ASAP7_75t_R g1661 ( 
.A(n_1322),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1254),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1254),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_1255),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1171),
.Y(n_1665)
);

CKINVDCx20_ASAP7_75t_R g1666 ( 
.A(n_1326),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1255),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_1268),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1419),
.B(n_992),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_1268),
.Y(n_1670)
);

CKINVDCx20_ASAP7_75t_R g1671 ( 
.A(n_1326),
.Y(n_1671)
);

INVxp33_ASAP7_75t_SL g1672 ( 
.A(n_1158),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1172),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1173),
.Y(n_1674)
);

INVxp67_ASAP7_75t_L g1675 ( 
.A(n_1401),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1271),
.Y(n_1676)
);

CKINVDCx20_ASAP7_75t_R g1677 ( 
.A(n_1328),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1271),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_1282),
.Y(n_1679)
);

CKINVDCx20_ASAP7_75t_R g1680 ( 
.A(n_1328),
.Y(n_1680)
);

CKINVDCx20_ASAP7_75t_R g1681 ( 
.A(n_1365),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_1282),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_1287),
.Y(n_1683)
);

CKINVDCx20_ASAP7_75t_R g1684 ( 
.A(n_1365),
.Y(n_1684)
);

NOR2xp67_ASAP7_75t_L g1685 ( 
.A(n_1419),
.B(n_812),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1176),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1231),
.B(n_703),
.Y(n_1687)
);

INVxp67_ASAP7_75t_L g1688 ( 
.A(n_1415),
.Y(n_1688)
);

INVxp33_ASAP7_75t_SL g1689 ( 
.A(n_1158),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1177),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_1287),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1296),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1179),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_1296),
.Y(n_1694)
);

BUFx2_ASAP7_75t_L g1695 ( 
.A(n_1154),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1348),
.B(n_992),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1182),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1311),
.Y(n_1698)
);

INVxp67_ASAP7_75t_SL g1699 ( 
.A(n_1404),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1311),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1165),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1411),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1443),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1459),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1556),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_1330),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1559),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1244),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1348),
.B(n_763),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1244),
.Y(n_1710)
);

INVxp67_ASAP7_75t_L g1711 ( 
.A(n_1428),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_1330),
.Y(n_1712)
);

CKINVDCx16_ASAP7_75t_R g1713 ( 
.A(n_1310),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1337),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1247),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1247),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_1337),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1341),
.Y(n_1718)
);

BUFx3_ASAP7_75t_L g1719 ( 
.A(n_1520),
.Y(n_1719)
);

CKINVDCx20_ASAP7_75t_R g1720 ( 
.A(n_1368),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1341),
.Y(n_1721)
);

CKINVDCx20_ASAP7_75t_R g1722 ( 
.A(n_1368),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1148),
.B(n_763),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_1351),
.Y(n_1724)
);

INVxp67_ASAP7_75t_SL g1725 ( 
.A(n_1354),
.Y(n_1725)
);

CKINVDCx20_ASAP7_75t_R g1726 ( 
.A(n_1372),
.Y(n_1726)
);

BUFx3_ASAP7_75t_L g1727 ( 
.A(n_1520),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1248),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1443),
.Y(n_1729)
);

CKINVDCx20_ASAP7_75t_R g1730 ( 
.A(n_1372),
.Y(n_1730)
);

NOR2xp67_ASAP7_75t_L g1731 ( 
.A(n_1351),
.B(n_697),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1148),
.B(n_763),
.Y(n_1732)
);

INVxp67_ASAP7_75t_SL g1733 ( 
.A(n_1461),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1248),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1443),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_1357),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1249),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1249),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1357),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1360),
.Y(n_1740)
);

CKINVDCx16_ASAP7_75t_R g1741 ( 
.A(n_1334),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_1360),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_1361),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1250),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1361),
.Y(n_1745)
);

CKINVDCx20_ASAP7_75t_R g1746 ( 
.A(n_1390),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1231),
.B(n_1155),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1250),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1560),
.Y(n_1749)
);

CKINVDCx16_ASAP7_75t_R g1750 ( 
.A(n_1430),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1560),
.Y(n_1751)
);

NOR2xp67_ASAP7_75t_L g1752 ( 
.A(n_1362),
.B(n_707),
.Y(n_1752)
);

CKINVDCx14_ASAP7_75t_R g1753 ( 
.A(n_1551),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1362),
.Y(n_1754)
);

CKINVDCx16_ASAP7_75t_R g1755 ( 
.A(n_1474),
.Y(n_1755)
);

INVxp67_ASAP7_75t_SL g1756 ( 
.A(n_1483),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_1379),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_1379),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_1416),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1312),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_1416),
.Y(n_1761)
);

CKINVDCx20_ASAP7_75t_R g1762 ( 
.A(n_1390),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1313),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1421),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1314),
.Y(n_1765)
);

CKINVDCx20_ASAP7_75t_R g1766 ( 
.A(n_1403),
.Y(n_1766)
);

NOR2xp67_ASAP7_75t_L g1767 ( 
.A(n_1421),
.B(n_719),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1316),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1317),
.Y(n_1769)
);

CKINVDCx16_ASAP7_75t_R g1770 ( 
.A(n_1481),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_1422),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1318),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1319),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1320),
.Y(n_1774)
);

CKINVDCx16_ASAP7_75t_R g1775 ( 
.A(n_1551),
.Y(n_1775)
);

HB1xp67_ASAP7_75t_L g1776 ( 
.A(n_1422),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_1437),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1376),
.B(n_723),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_1437),
.Y(n_1779)
);

CKINVDCx20_ASAP7_75t_R g1780 ( 
.A(n_1403),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_1452),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1499),
.B(n_1378),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1324),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_1452),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1325),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1335),
.B(n_810),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1327),
.Y(n_1787)
);

INVxp33_ASAP7_75t_L g1788 ( 
.A(n_1253),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_1453),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1522),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1329),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_1453),
.Y(n_1792)
);

CKINVDCx20_ASAP7_75t_R g1793 ( 
.A(n_1407),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1331),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1376),
.B(n_878),
.Y(n_1795)
);

NOR2xp67_ASAP7_75t_L g1796 ( 
.A(n_1464),
.B(n_968),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_1464),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_1465),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1332),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1333),
.Y(n_1800)
);

CKINVDCx20_ASAP7_75t_R g1801 ( 
.A(n_1407),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1336),
.Y(n_1802)
);

CKINVDCx20_ASAP7_75t_R g1803 ( 
.A(n_1414),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1338),
.Y(n_1804)
);

NOR2xp67_ASAP7_75t_L g1805 ( 
.A(n_1465),
.B(n_1472),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1339),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_1472),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_1476),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_1476),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_1477),
.Y(n_1810)
);

CKINVDCx20_ASAP7_75t_R g1811 ( 
.A(n_1414),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1340),
.Y(n_1812)
);

HB1xp67_ASAP7_75t_L g1813 ( 
.A(n_1477),
.Y(n_1813)
);

INVxp33_ASAP7_75t_SL g1814 ( 
.A(n_1486),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1522),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1342),
.Y(n_1816)
);

INVxp67_ASAP7_75t_SL g1817 ( 
.A(n_1522),
.Y(n_1817)
);

NOR2xp67_ASAP7_75t_L g1818 ( 
.A(n_1486),
.B(n_989),
.Y(n_1818)
);

BUFx2_ASAP7_75t_L g1819 ( 
.A(n_1154),
.Y(n_1819)
);

CKINVDCx20_ASAP7_75t_R g1820 ( 
.A(n_1427),
.Y(n_1820)
);

CKINVDCx16_ASAP7_75t_R g1821 ( 
.A(n_1553),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1343),
.Y(n_1822)
);

CKINVDCx14_ASAP7_75t_R g1823 ( 
.A(n_1553),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_1491),
.Y(n_1824)
);

CKINVDCx5p33_ASAP7_75t_R g1825 ( 
.A(n_1491),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1345),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_1492),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1346),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1347),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1349),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1492),
.Y(n_1831)
);

CKINVDCx5p33_ASAP7_75t_R g1832 ( 
.A(n_1495),
.Y(n_1832)
);

CKINVDCx20_ASAP7_75t_R g1833 ( 
.A(n_1427),
.Y(n_1833)
);

CKINVDCx20_ASAP7_75t_R g1834 ( 
.A(n_1451),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1352),
.Y(n_1835)
);

CKINVDCx5p33_ASAP7_75t_R g1836 ( 
.A(n_1495),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_1500),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1356),
.Y(n_1838)
);

CKINVDCx20_ASAP7_75t_R g1839 ( 
.A(n_1451),
.Y(n_1839)
);

CKINVDCx20_ASAP7_75t_R g1840 ( 
.A(n_1457),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_1500),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1359),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_1502),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1502),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_1503),
.Y(n_1845)
);

CKINVDCx20_ASAP7_75t_R g1846 ( 
.A(n_1457),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_1503),
.Y(n_1847)
);

CKINVDCx20_ASAP7_75t_R g1848 ( 
.A(n_1526),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1363),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1364),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_1517),
.Y(n_1851)
);

CKINVDCx16_ASAP7_75t_R g1852 ( 
.A(n_1163),
.Y(n_1852)
);

INVxp33_ASAP7_75t_L g1853 ( 
.A(n_1257),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_1517),
.Y(n_1854)
);

INVxp33_ASAP7_75t_L g1855 ( 
.A(n_1298),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1366),
.Y(n_1856)
);

BUFx2_ASAP7_75t_L g1857 ( 
.A(n_1163),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1367),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_1518),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_1518),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1369),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1370),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1371),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_1555),
.Y(n_1864)
);

INVx1_ASAP7_75t_SL g1865 ( 
.A(n_1191),
.Y(n_1865)
);

CKINVDCx5p33_ASAP7_75t_R g1866 ( 
.A(n_1555),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1480),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1374),
.Y(n_1868)
);

NOR2xp67_ASAP7_75t_L g1869 ( 
.A(n_1506),
.B(n_1017),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_L g1870 ( 
.A(n_1399),
.B(n_1435),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_1151),
.Y(n_1871)
);

CKINVDCx20_ASAP7_75t_R g1872 ( 
.A(n_1526),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1375),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1377),
.Y(n_1874)
);

INVxp67_ASAP7_75t_L g1875 ( 
.A(n_1460),
.Y(n_1875)
);

CKINVDCx5p33_ASAP7_75t_R g1876 ( 
.A(n_1399),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1480),
.Y(n_1877)
);

OR2x2_ASAP7_75t_L g1878 ( 
.A(n_1300),
.B(n_703),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1380),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1383),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1384),
.Y(n_1881)
);

BUFx6f_ASAP7_75t_L g1882 ( 
.A(n_1480),
.Y(n_1882)
);

INVxp67_ASAP7_75t_SL g1883 ( 
.A(n_1484),
.Y(n_1883)
);

NOR2xp67_ASAP7_75t_L g1884 ( 
.A(n_1536),
.B(n_1538),
.Y(n_1884)
);

INVxp67_ASAP7_75t_L g1885 ( 
.A(n_1523),
.Y(n_1885)
);

CKINVDCx20_ASAP7_75t_R g1886 ( 
.A(n_1528),
.Y(n_1886)
);

INVxp67_ASAP7_75t_L g1887 ( 
.A(n_1534),
.Y(n_1887)
);

INVxp67_ASAP7_75t_L g1888 ( 
.A(n_1278),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1387),
.Y(n_1889)
);

CKINVDCx20_ASAP7_75t_R g1890 ( 
.A(n_1528),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1484),
.Y(n_1891)
);

HB1xp67_ASAP7_75t_L g1892 ( 
.A(n_1191),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1388),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_1435),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_1494),
.Y(n_1895)
);

INVxp67_ASAP7_75t_L g1896 ( 
.A(n_1278),
.Y(n_1896)
);

INVxp67_ASAP7_75t_L g1897 ( 
.A(n_1278),
.Y(n_1897)
);

INVxp33_ASAP7_75t_L g1898 ( 
.A(n_1353),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1389),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1392),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1335),
.B(n_1025),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1394),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1395),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_L g1904 ( 
.A(n_1494),
.B(n_1037),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1396),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_1509),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1397),
.Y(n_1907)
);

BUFx3_ASAP7_75t_L g1908 ( 
.A(n_1484),
.Y(n_1908)
);

INVxp33_ASAP7_75t_SL g1909 ( 
.A(n_1144),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1398),
.Y(n_1910)
);

HB1xp67_ASAP7_75t_L g1911 ( 
.A(n_1202),
.Y(n_1911)
);

INVxp67_ASAP7_75t_SL g1912 ( 
.A(n_1484),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1400),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_1509),
.Y(n_1914)
);

HB1xp67_ASAP7_75t_L g1915 ( 
.A(n_1202),
.Y(n_1915)
);

INVxp33_ASAP7_75t_L g1916 ( 
.A(n_1386),
.Y(n_1916)
);

CKINVDCx20_ASAP7_75t_R g1917 ( 
.A(n_1532),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_1524),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1406),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1649),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1567),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1699),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1708),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_SL g1924 ( 
.A(n_1909),
.B(n_1524),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1710),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1715),
.Y(n_1926)
);

INVx3_ASAP7_75t_L g1927 ( 
.A(n_1908),
.Y(n_1927)
);

OAI21x1_ASAP7_75t_L g1928 ( 
.A1(n_1610),
.A2(n_1204),
.B(n_1175),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1567),
.Y(n_1929)
);

INVxp67_ASAP7_75t_L g1930 ( 
.A(n_1644),
.Y(n_1930)
);

INVx3_ASAP7_75t_L g1931 ( 
.A(n_1908),
.Y(n_1931)
);

CKINVDCx5p33_ASAP7_75t_R g1932 ( 
.A(n_1871),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1639),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1716),
.Y(n_1934)
);

INVx3_ASAP7_75t_L g1935 ( 
.A(n_1639),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1568),
.B(n_1548),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_1595),
.Y(n_1937)
);

INVx3_ASAP7_75t_L g1938 ( 
.A(n_1701),
.Y(n_1938)
);

BUFx2_ASAP7_75t_L g1939 ( 
.A(n_1583),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1709),
.B(n_1548),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1701),
.Y(n_1941)
);

XNOR2xp5_ASAP7_75t_L g1942 ( 
.A(n_1564),
.B(n_1532),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1703),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1703),
.Y(n_1944)
);

BUFx6f_ASAP7_75t_L g1945 ( 
.A(n_1571),
.Y(n_1945)
);

AND2x4_ASAP7_75t_L g1946 ( 
.A(n_1594),
.B(n_1216),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1898),
.B(n_1496),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1728),
.Y(n_1948)
);

INVx3_ASAP7_75t_L g1949 ( 
.A(n_1729),
.Y(n_1949)
);

OAI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1909),
.A2(n_1199),
.B1(n_1217),
.B2(n_1185),
.Y(n_1950)
);

BUFx6f_ASAP7_75t_L g1951 ( 
.A(n_1571),
.Y(n_1951)
);

AND2x4_ASAP7_75t_L g1952 ( 
.A(n_1596),
.B(n_1549),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_1597),
.Y(n_1953)
);

AND2x4_ASAP7_75t_L g1954 ( 
.A(n_1603),
.B(n_1161),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1729),
.Y(n_1955)
);

AND2x4_ASAP7_75t_L g1956 ( 
.A(n_1685),
.B(n_1193),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1735),
.Y(n_1957)
);

BUFx6f_ASAP7_75t_L g1958 ( 
.A(n_1571),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1605),
.B(n_1405),
.Y(n_1959)
);

BUFx3_ASAP7_75t_L g1960 ( 
.A(n_1719),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1734),
.Y(n_1961)
);

CKINVDCx20_ASAP7_75t_R g1962 ( 
.A(n_1564),
.Y(n_1962)
);

BUFx6f_ASAP7_75t_L g1963 ( 
.A(n_1571),
.Y(n_1963)
);

BUFx3_ASAP7_75t_L g1964 ( 
.A(n_1719),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1737),
.Y(n_1965)
);

INVx3_ASAP7_75t_L g1966 ( 
.A(n_1735),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_R g1967 ( 
.A(n_1601),
.B(n_1214),
.Y(n_1967)
);

BUFx6f_ASAP7_75t_L g1968 ( 
.A(n_1571),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1738),
.Y(n_1969)
);

HB1xp67_ASAP7_75t_L g1970 ( 
.A(n_1916),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1790),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1744),
.Y(n_1972)
);

AND2x4_ASAP7_75t_L g1973 ( 
.A(n_1570),
.B(n_1323),
.Y(n_1973)
);

CKINVDCx6p67_ASAP7_75t_R g1974 ( 
.A(n_1608),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1884),
.B(n_1405),
.Y(n_1975)
);

INVx3_ASAP7_75t_L g1976 ( 
.A(n_1790),
.Y(n_1976)
);

INVxp33_ASAP7_75t_SL g1977 ( 
.A(n_1612),
.Y(n_1977)
);

INVx3_ASAP7_75t_L g1978 ( 
.A(n_1815),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1815),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_1601),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1748),
.Y(n_1981)
);

BUFx6f_ASAP7_75t_L g1982 ( 
.A(n_1656),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1749),
.Y(n_1983)
);

BUFx6f_ASAP7_75t_L g1984 ( 
.A(n_1656),
.Y(n_1984)
);

CKINVDCx5p33_ASAP7_75t_R g1985 ( 
.A(n_1604),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1751),
.Y(n_1986)
);

INVx4_ASAP7_75t_L g1987 ( 
.A(n_1576),
.Y(n_1987)
);

OAI22xp5_ASAP7_75t_SL g1988 ( 
.A1(n_1566),
.A2(n_1214),
.B1(n_1917),
.B2(n_1573),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1867),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1593),
.Y(n_1990)
);

BUFx6f_ASAP7_75t_L g1991 ( 
.A(n_1656),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1611),
.Y(n_1992)
);

CKINVDCx20_ASAP7_75t_R g1993 ( 
.A(n_1566),
.Y(n_1993)
);

CKINVDCx11_ASAP7_75t_R g1994 ( 
.A(n_1572),
.Y(n_1994)
);

CKINVDCx20_ASAP7_75t_R g1995 ( 
.A(n_1572),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1647),
.B(n_1562),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1867),
.Y(n_1997)
);

BUFx3_ASAP7_75t_L g1998 ( 
.A(n_1727),
.Y(n_1998)
);

INVx3_ASAP7_75t_L g1999 ( 
.A(n_1656),
.Y(n_1999)
);

INVx3_ASAP7_75t_L g2000 ( 
.A(n_1656),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1622),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1623),
.Y(n_2002)
);

CKINVDCx20_ASAP7_75t_R g2003 ( 
.A(n_1573),
.Y(n_2003)
);

BUFx6f_ASAP7_75t_L g2004 ( 
.A(n_1882),
.Y(n_2004)
);

AND2x4_ASAP7_75t_L g2005 ( 
.A(n_1580),
.B(n_1439),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1877),
.Y(n_2006)
);

NAND2x1_ASAP7_75t_L g2007 ( 
.A(n_1576),
.B(n_1373),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_SL g2008 ( 
.A(n_1696),
.B(n_1109),
.Y(n_2008)
);

CKINVDCx8_ASAP7_75t_R g2009 ( 
.A(n_1621),
.Y(n_2009)
);

XNOR2xp5_ASAP7_75t_L g2010 ( 
.A(n_1579),
.B(n_1590),
.Y(n_2010)
);

CKINVDCx5p33_ASAP7_75t_R g2011 ( 
.A(n_1604),
.Y(n_2011)
);

CKINVDCx20_ASAP7_75t_R g2012 ( 
.A(n_1579),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1760),
.Y(n_2013)
);

INVx3_ASAP7_75t_L g2014 ( 
.A(n_1882),
.Y(n_2014)
);

INVxp67_ASAP7_75t_SL g2015 ( 
.A(n_1576),
.Y(n_2015)
);

CKINVDCx20_ASAP7_75t_R g2016 ( 
.A(n_1590),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1565),
.B(n_1439),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1763),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1765),
.Y(n_2019)
);

BUFx3_ASAP7_75t_L g2020 ( 
.A(n_1727),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1768),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1769),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1877),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1772),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1773),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1702),
.B(n_1704),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_R g2027 ( 
.A(n_1606),
.B(n_1308),
.Y(n_2027)
);

CKINVDCx5p33_ASAP7_75t_R g2028 ( 
.A(n_1606),
.Y(n_2028)
);

INVx3_ASAP7_75t_L g2029 ( 
.A(n_1882),
.Y(n_2029)
);

CKINVDCx20_ASAP7_75t_R g2030 ( 
.A(n_1598),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1774),
.Y(n_2031)
);

CKINVDCx11_ASAP7_75t_R g2032 ( 
.A(n_1598),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1783),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1785),
.Y(n_2034)
);

BUFx6f_ASAP7_75t_L g2035 ( 
.A(n_1882),
.Y(n_2035)
);

INVx3_ASAP7_75t_L g2036 ( 
.A(n_1882),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1891),
.Y(n_2037)
);

CKINVDCx5p33_ASAP7_75t_R g2038 ( 
.A(n_1609),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1569),
.B(n_1498),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1891),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1787),
.Y(n_2041)
);

BUFx6f_ASAP7_75t_L g2042 ( 
.A(n_1591),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1791),
.Y(n_2043)
);

NAND2xp33_ASAP7_75t_SL g2044 ( 
.A(n_1612),
.B(n_1036),
.Y(n_2044)
);

NOR2xp33_ASAP7_75t_L g2045 ( 
.A(n_1581),
.B(n_1185),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1705),
.B(n_1498),
.Y(n_2046)
);

AOI22xp5_ASAP7_75t_L g2047 ( 
.A1(n_1778),
.A2(n_1217),
.B1(n_1199),
.B2(n_1188),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1707),
.B(n_1194),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1794),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1592),
.Y(n_2050)
);

INVx3_ASAP7_75t_L g2051 ( 
.A(n_1627),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1799),
.Y(n_2052)
);

CKINVDCx20_ASAP7_75t_R g2053 ( 
.A(n_1607),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1800),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1629),
.Y(n_2055)
);

HB1xp67_ASAP7_75t_L g2056 ( 
.A(n_1574),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1631),
.Y(n_2057)
);

AND2x4_ASAP7_75t_L g2058 ( 
.A(n_1582),
.B(n_1545),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1634),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1802),
.Y(n_2060)
);

INVx3_ASAP7_75t_L g2061 ( 
.A(n_1635),
.Y(n_2061)
);

OAI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_1870),
.A2(n_1219),
.B1(n_1263),
.B2(n_1170),
.Y(n_2062)
);

BUFx6f_ASAP7_75t_L g2063 ( 
.A(n_1636),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1804),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_1609),
.Y(n_2065)
);

BUFx3_ASAP7_75t_L g2066 ( 
.A(n_1646),
.Y(n_2066)
);

BUFx6f_ASAP7_75t_L g2067 ( 
.A(n_1650),
.Y(n_2067)
);

BUFx10_ASAP7_75t_L g2068 ( 
.A(n_1795),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_SL g2069 ( 
.A(n_1904),
.B(n_1109),
.Y(n_2069)
);

AND2x4_ASAP7_75t_L g2070 ( 
.A(n_1586),
.B(n_1587),
.Y(n_2070)
);

BUFx6f_ASAP7_75t_L g2071 ( 
.A(n_1651),
.Y(n_2071)
);

BUFx6f_ASAP7_75t_L g2072 ( 
.A(n_1657),
.Y(n_2072)
);

BUFx6f_ASAP7_75t_L g2073 ( 
.A(n_1658),
.Y(n_2073)
);

OR2x2_ASAP7_75t_L g2074 ( 
.A(n_1687),
.B(n_1279),
.Y(n_2074)
);

NOR2xp33_ASAP7_75t_R g2075 ( 
.A(n_1641),
.B(n_1309),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1723),
.B(n_1408),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1659),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1660),
.Y(n_2078)
);

CKINVDCx8_ASAP7_75t_R g2079 ( 
.A(n_1713),
.Y(n_2079)
);

INVx3_ASAP7_75t_L g2080 ( 
.A(n_1665),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_SL g2081 ( 
.A(n_1805),
.B(n_1044),
.Y(n_2081)
);

HB1xp67_ASAP7_75t_L g2082 ( 
.A(n_1575),
.Y(n_2082)
);

CKINVDCx5p33_ASAP7_75t_R g2083 ( 
.A(n_1563),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_1673),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_1732),
.B(n_1806),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1812),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1725),
.B(n_1195),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1816),
.Y(n_2088)
);

CKINVDCx20_ASAP7_75t_R g2089 ( 
.A(n_1607),
.Y(n_2089)
);

NOR2xp33_ASAP7_75t_R g2090 ( 
.A(n_1643),
.B(n_1106),
.Y(n_2090)
);

INVx3_ASAP7_75t_L g2091 ( 
.A(n_1674),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_1822),
.B(n_1410),
.Y(n_2092)
);

OAI21x1_ASAP7_75t_L g2093 ( 
.A1(n_1624),
.A2(n_1204),
.B(n_1175),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1733),
.B(n_1196),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1826),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_1828),
.B(n_1412),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1829),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1830),
.Y(n_2098)
);

CKINVDCx5p33_ASAP7_75t_R g2099 ( 
.A(n_1578),
.Y(n_2099)
);

CKINVDCx20_ASAP7_75t_R g2100 ( 
.A(n_1626),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1835),
.Y(n_2101)
);

OAI22xp5_ASAP7_75t_L g2102 ( 
.A1(n_1613),
.A2(n_1306),
.B1(n_790),
.B2(n_870),
.Y(n_2102)
);

BUFx6f_ASAP7_75t_L g2103 ( 
.A(n_1686),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_SL g2104 ( 
.A(n_1613),
.B(n_1108),
.Y(n_2104)
);

BUFx3_ASAP7_75t_L g2105 ( 
.A(n_1690),
.Y(n_2105)
);

BUFx3_ASAP7_75t_L g2106 ( 
.A(n_1693),
.Y(n_2106)
);

HB1xp67_ASAP7_75t_L g2107 ( 
.A(n_1584),
.Y(n_2107)
);

INVx3_ASAP7_75t_L g2108 ( 
.A(n_1697),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_1838),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_1756),
.B(n_1197),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1842),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1817),
.B(n_1577),
.Y(n_2112)
);

OAI22xp5_ASAP7_75t_L g2113 ( 
.A1(n_1615),
.A2(n_790),
.B1(n_870),
.B2(n_730),
.Y(n_2113)
);

HB1xp67_ASAP7_75t_L g2114 ( 
.A(n_1892),
.Y(n_2114)
);

HB1xp67_ASAP7_75t_L g2115 ( 
.A(n_1911),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1849),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1850),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_1856),
.B(n_1858),
.Y(n_2118)
);

BUFx6f_ASAP7_75t_L g2119 ( 
.A(n_1861),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1862),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1863),
.Y(n_2121)
);

CKINVDCx5p33_ASAP7_75t_R g2122 ( 
.A(n_1615),
.Y(n_2122)
);

BUFx3_ASAP7_75t_L g2123 ( 
.A(n_1868),
.Y(n_2123)
);

INVx3_ASAP7_75t_L g2124 ( 
.A(n_1873),
.Y(n_2124)
);

BUFx2_ASAP7_75t_L g2125 ( 
.A(n_1712),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1874),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1879),
.Y(n_2127)
);

NOR2xp33_ASAP7_75t_L g2128 ( 
.A(n_1589),
.B(n_1413),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1880),
.Y(n_2129)
);

CKINVDCx16_ASAP7_75t_R g2130 ( 
.A(n_1741),
.Y(n_2130)
);

AND2x4_ASAP7_75t_L g2131 ( 
.A(n_1600),
.B(n_1558),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_1881),
.B(n_1417),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1889),
.Y(n_2133)
);

NOR2xp67_ASAP7_75t_L g2134 ( 
.A(n_1888),
.B(n_1418),
.Y(n_2134)
);

AOI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_1630),
.A2(n_901),
.B1(n_973),
.B2(n_730),
.Y(n_2135)
);

NOR2xp33_ASAP7_75t_L g2136 ( 
.A(n_1786),
.B(n_1420),
.Y(n_2136)
);

BUFx6f_ASAP7_75t_L g2137 ( 
.A(n_1919),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1893),
.Y(n_2138)
);

CKINVDCx20_ASAP7_75t_R g2139 ( 
.A(n_1626),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1899),
.Y(n_2140)
);

INVx3_ASAP7_75t_L g2141 ( 
.A(n_1900),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1669),
.B(n_1198),
.Y(n_2142)
);

BUFx6f_ASAP7_75t_L g2143 ( 
.A(n_1902),
.Y(n_2143)
);

OAI22xp5_ASAP7_75t_SL g2144 ( 
.A1(n_1632),
.A2(n_1917),
.B1(n_1640),
.B2(n_1642),
.Y(n_2144)
);

AND2x4_ASAP7_75t_L g2145 ( 
.A(n_1903),
.B(n_1539),
.Y(n_2145)
);

CKINVDCx5p33_ASAP7_75t_R g2146 ( 
.A(n_1712),
.Y(n_2146)
);

INVx3_ASAP7_75t_L g2147 ( 
.A(n_1905),
.Y(n_2147)
);

AND2x4_ASAP7_75t_L g2148 ( 
.A(n_1907),
.B(n_1541),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1910),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1901),
.B(n_1200),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1913),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_1618),
.B(n_1423),
.Y(n_2152)
);

CKINVDCx5p33_ASAP7_75t_R g2153 ( 
.A(n_1717),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_1619),
.B(n_1424),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1625),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1883),
.Y(n_2156)
);

XNOR2x2_ASAP7_75t_R g2157 ( 
.A(n_1753),
.B(n_4),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1912),
.Y(n_2158)
);

OAI22x1_ASAP7_75t_L g2159 ( 
.A1(n_1675),
.A2(n_973),
.B1(n_1045),
.B2(n_901),
.Y(n_2159)
);

AND2x4_ASAP7_75t_L g2160 ( 
.A(n_1782),
.B(n_1550),
.Y(n_2160)
);

BUFx6f_ASAP7_75t_L g2161 ( 
.A(n_1648),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1869),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1731),
.Y(n_2163)
);

AND2x4_ASAP7_75t_L g2164 ( 
.A(n_1752),
.B(n_1554),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_1688),
.B(n_1425),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1767),
.Y(n_2166)
);

HB1xp67_ASAP7_75t_L g2167 ( 
.A(n_1915),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1711),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_1796),
.B(n_1818),
.Y(n_2169)
);

CKINVDCx5p33_ASAP7_75t_R g2170 ( 
.A(n_1717),
.Y(n_2170)
);

CKINVDCx5p33_ASAP7_75t_R g2171 ( 
.A(n_1807),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1875),
.Y(n_2172)
);

INVx2_ASAP7_75t_SL g2173 ( 
.A(n_1878),
.Y(n_2173)
);

BUFx2_ASAP7_75t_L g2174 ( 
.A(n_1807),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1678),
.Y(n_2175)
);

INVx6_ASAP7_75t_L g2176 ( 
.A(n_1750),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_1896),
.B(n_1201),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_1885),
.Y(n_2178)
);

BUFx6f_ASAP7_75t_L g2179 ( 
.A(n_1653),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1887),
.Y(n_2180)
);

OAI22xp33_ASAP7_75t_L g2181 ( 
.A1(n_1808),
.A2(n_1062),
.B1(n_1079),
.B2(n_1045),
.Y(n_2181)
);

AND2x6_ASAP7_75t_L g2182 ( 
.A(n_1865),
.B(n_931),
.Y(n_2182)
);

BUFx6f_ASAP7_75t_L g2183 ( 
.A(n_1654),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1692),
.Y(n_2184)
);

NOR2xp33_ASAP7_75t_L g2185 ( 
.A(n_1897),
.B(n_1426),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1747),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1714),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1718),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1721),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1739),
.Y(n_2190)
);

INVx3_ASAP7_75t_L g2191 ( 
.A(n_1655),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1740),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_1662),
.B(n_1663),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_1754),
.Y(n_2194)
);

AND2x2_ASAP7_75t_SL g2195 ( 
.A(n_1755),
.B(n_931),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1764),
.Y(n_2196)
);

CKINVDCx5p33_ASAP7_75t_R g2197 ( 
.A(n_1808),
.Y(n_2197)
);

BUFx6f_ASAP7_75t_L g2198 ( 
.A(n_1664),
.Y(n_2198)
);

INVx1_ASAP7_75t_SL g2199 ( 
.A(n_1599),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_1776),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1813),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1831),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_1667),
.B(n_1205),
.Y(n_2203)
);

HB1xp67_ASAP7_75t_L g2204 ( 
.A(n_1695),
.Y(n_2204)
);

HB1xp67_ASAP7_75t_L g2205 ( 
.A(n_1819),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1668),
.Y(n_2206)
);

INVx3_ASAP7_75t_L g2207 ( 
.A(n_1670),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1588),
.Y(n_2208)
);

BUFx2_ASAP7_75t_L g2209 ( 
.A(n_1809),
.Y(n_2209)
);

AND3x2_ASAP7_75t_L g2210 ( 
.A(n_1602),
.B(n_933),
.C(n_932),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1616),
.Y(n_2211)
);

OA21x2_ASAP7_75t_L g2212 ( 
.A1(n_1617),
.A2(n_1552),
.B(n_1222),
.Y(n_2212)
);

CKINVDCx5p33_ASAP7_75t_R g2213 ( 
.A(n_1809),
.Y(n_2213)
);

INVx4_ASAP7_75t_L g2214 ( 
.A(n_1676),
.Y(n_2214)
);

CKINVDCx5p33_ASAP7_75t_R g2215 ( 
.A(n_1810),
.Y(n_2215)
);

NOR2xp33_ASAP7_75t_L g2216 ( 
.A(n_1814),
.B(n_1429),
.Y(n_2216)
);

AOI22xp5_ASAP7_75t_L g2217 ( 
.A1(n_1814),
.A2(n_1079),
.B1(n_1115),
.B2(n_1062),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1679),
.Y(n_2218)
);

BUFx6f_ASAP7_75t_L g2219 ( 
.A(n_1682),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_1683),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_1691),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1694),
.Y(n_2222)
);

INVx3_ASAP7_75t_L g2223 ( 
.A(n_1698),
.Y(n_2223)
);

CKINVDCx20_ASAP7_75t_R g2224 ( 
.A(n_1632),
.Y(n_2224)
);

AND2x6_ASAP7_75t_L g2225 ( 
.A(n_1672),
.B(n_932),
.Y(n_2225)
);

BUFx6f_ASAP7_75t_L g2226 ( 
.A(n_1700),
.Y(n_2226)
);

HB1xp67_ASAP7_75t_L g2227 ( 
.A(n_1857),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_1788),
.B(n_1431),
.Y(n_2228)
);

AOI22xp5_ASAP7_75t_L g2229 ( 
.A1(n_1810),
.A2(n_1123),
.B1(n_1115),
.B2(n_743),
.Y(n_2229)
);

OAI22xp5_ASAP7_75t_SL g2230 ( 
.A1(n_1637),
.A2(n_1123),
.B1(n_769),
.B2(n_789),
.Y(n_2230)
);

INVx3_ASAP7_75t_L g2231 ( 
.A(n_1706),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1724),
.Y(n_2232)
);

BUFx2_ASAP7_75t_L g2233 ( 
.A(n_1824),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_1736),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1742),
.Y(n_2235)
);

AND2x4_ASAP7_75t_L g2236 ( 
.A(n_1614),
.B(n_1557),
.Y(n_2236)
);

INVx4_ASAP7_75t_L g2237 ( 
.A(n_1743),
.Y(n_2237)
);

INVx3_ASAP7_75t_L g2238 ( 
.A(n_1745),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1757),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1758),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_1759),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_1853),
.B(n_1440),
.Y(n_2242)
);

INVx3_ASAP7_75t_L g2243 ( 
.A(n_1761),
.Y(n_2243)
);

AND2x4_ASAP7_75t_L g2244 ( 
.A(n_1645),
.B(n_1561),
.Y(n_2244)
);

BUFx6f_ASAP7_75t_L g2245 ( 
.A(n_1771),
.Y(n_2245)
);

INVxp33_ASAP7_75t_SL g2246 ( 
.A(n_1824),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_1777),
.Y(n_2247)
);

CKINVDCx16_ASAP7_75t_R g2248 ( 
.A(n_1770),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1779),
.Y(n_2249)
);

AND2x4_ASAP7_75t_L g2250 ( 
.A(n_1652),
.B(n_1441),
.Y(n_2250)
);

CKINVDCx5p33_ASAP7_75t_R g2251 ( 
.A(n_1825),
.Y(n_2251)
);

BUFx6f_ASAP7_75t_L g2252 ( 
.A(n_1781),
.Y(n_2252)
);

CKINVDCx20_ASAP7_75t_R g2253 ( 
.A(n_1637),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_1784),
.Y(n_2254)
);

CKINVDCx5p33_ASAP7_75t_R g2255 ( 
.A(n_1825),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1789),
.Y(n_2256)
);

HB1xp67_ASAP7_75t_L g2257 ( 
.A(n_1827),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1792),
.Y(n_2258)
);

OAI22xp5_ASAP7_75t_L g2259 ( 
.A1(n_1672),
.A2(n_772),
.B1(n_813),
.B2(n_749),
.Y(n_2259)
);

AOI22xp5_ASAP7_75t_L g2260 ( 
.A1(n_1827),
.A2(n_744),
.B1(n_747),
.B2(n_741),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1797),
.Y(n_2261)
);

NOR2x1_ASAP7_75t_L g2262 ( 
.A(n_1689),
.B(n_1533),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_1798),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_1847),
.Y(n_2264)
);

AND2x4_ASAP7_75t_L g2265 ( 
.A(n_1832),
.B(n_1535),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_1851),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1854),
.Y(n_2267)
);

AND2x2_ASAP7_75t_L g2268 ( 
.A(n_1855),
.B(n_1444),
.Y(n_2268)
);

CKINVDCx6p67_ASAP7_75t_R g2269 ( 
.A(n_1852),
.Y(n_2269)
);

AOI22xp5_ASAP7_75t_L g2270 ( 
.A1(n_1832),
.A2(n_751),
.B1(n_754),
.B2(n_748),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1859),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_1860),
.Y(n_2272)
);

CKINVDCx8_ASAP7_75t_R g2273 ( 
.A(n_1775),
.Y(n_2273)
);

BUFx6f_ASAP7_75t_L g2274 ( 
.A(n_1864),
.Y(n_2274)
);

CKINVDCx20_ASAP7_75t_R g2275 ( 
.A(n_1640),
.Y(n_2275)
);

INVxp67_ASAP7_75t_L g2276 ( 
.A(n_1836),
.Y(n_2276)
);

AND2x4_ASAP7_75t_L g2277 ( 
.A(n_1836),
.B(n_1544),
.Y(n_2277)
);

AND2x4_ASAP7_75t_L g2278 ( 
.A(n_1837),
.B(n_1547),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1866),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_1837),
.B(n_1206),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1841),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_1841),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1843),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_1843),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_1844),
.Y(n_2285)
);

INVx3_ASAP7_75t_L g2286 ( 
.A(n_1844),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_1845),
.B(n_1445),
.Y(n_2287)
);

AOI22xp5_ASAP7_75t_L g2288 ( 
.A1(n_1845),
.A2(n_759),
.B1(n_765),
.B2(n_758),
.Y(n_2288)
);

BUFx2_ASAP7_75t_L g2289 ( 
.A(n_1617),
.Y(n_2289)
);

AND2x4_ASAP7_75t_L g2290 ( 
.A(n_1620),
.B(n_1446),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_1876),
.B(n_1207),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_1620),
.Y(n_2292)
);

AND2x6_ASAP7_75t_L g2293 ( 
.A(n_1689),
.B(n_933),
.Y(n_2293)
);

HB1xp67_ASAP7_75t_L g2294 ( 
.A(n_1628),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1628),
.Y(n_2295)
);

NAND2x1_ASAP7_75t_L g2296 ( 
.A(n_1633),
.B(n_1213),
.Y(n_2296)
);

INVx3_ASAP7_75t_L g2297 ( 
.A(n_1633),
.Y(n_2297)
);

AND2x4_ASAP7_75t_L g2298 ( 
.A(n_1638),
.B(n_1529),
.Y(n_2298)
);

HB1xp67_ASAP7_75t_L g2299 ( 
.A(n_1638),
.Y(n_2299)
);

CKINVDCx5p33_ASAP7_75t_R g2300 ( 
.A(n_1585),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_1918),
.B(n_1447),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_1894),
.Y(n_2302)
);

BUFx6f_ASAP7_75t_L g2303 ( 
.A(n_1895),
.Y(n_2303)
);

BUFx6f_ASAP7_75t_L g2304 ( 
.A(n_1906),
.Y(n_2304)
);

CKINVDCx5p33_ASAP7_75t_R g2305 ( 
.A(n_1914),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_1918),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_1821),
.Y(n_2307)
);

CKINVDCx5p33_ASAP7_75t_R g2308 ( 
.A(n_1823),
.Y(n_2308)
);

NOR2xp33_ASAP7_75t_L g2309 ( 
.A(n_1642),
.B(n_1449),
.Y(n_2309)
);

BUFx6f_ASAP7_75t_L g2310 ( 
.A(n_1661),
.Y(n_2310)
);

NOR2xp33_ASAP7_75t_L g2311 ( 
.A(n_1661),
.B(n_1450),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_1666),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_SL g2313 ( 
.A(n_1666),
.B(n_1085),
.Y(n_2313)
);

OAI22xp5_ASAP7_75t_SL g2314 ( 
.A1(n_1671),
.A2(n_803),
.B1(n_820),
.B2(n_777),
.Y(n_2314)
);

INVx3_ASAP7_75t_L g2315 ( 
.A(n_1671),
.Y(n_2315)
);

INVxp67_ASAP7_75t_L g2316 ( 
.A(n_1677),
.Y(n_2316)
);

CKINVDCx20_ASAP7_75t_R g2317 ( 
.A(n_1677),
.Y(n_2317)
);

INVx3_ASAP7_75t_L g2318 ( 
.A(n_1680),
.Y(n_2318)
);

INVx3_ASAP7_75t_L g2319 ( 
.A(n_1680),
.Y(n_2319)
);

NOR2xp33_ASAP7_75t_R g2320 ( 
.A(n_1681),
.B(n_1454),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2118),
.Y(n_2321)
);

AOI22xp5_ASAP7_75t_L g2322 ( 
.A1(n_2225),
.A2(n_1085),
.B1(n_768),
.B2(n_774),
.Y(n_2322)
);

HB1xp67_ASAP7_75t_L g2323 ( 
.A(n_1970),
.Y(n_2323)
);

BUFx6f_ASAP7_75t_L g2324 ( 
.A(n_1945),
.Y(n_2324)
);

BUFx2_ASAP7_75t_L g2325 ( 
.A(n_2320),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_1947),
.B(n_1455),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_1921),
.Y(n_2327)
);

INVxp67_ASAP7_75t_L g2328 ( 
.A(n_1939),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2136),
.B(n_938),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_1921),
.Y(n_2330)
);

INVx1_ASAP7_75t_SL g2331 ( 
.A(n_1947),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_1929),
.Y(n_2332)
);

NOR2xp33_ASAP7_75t_L g2333 ( 
.A(n_1936),
.B(n_766),
.Y(n_2333)
);

BUFx6f_ASAP7_75t_L g2334 ( 
.A(n_1945),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2118),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2055),
.Y(n_2336)
);

OAI22xp33_ASAP7_75t_L g2337 ( 
.A1(n_2047),
.A2(n_943),
.B1(n_951),
.B2(n_938),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2055),
.Y(n_2338)
);

BUFx6f_ASAP7_75t_L g2339 ( 
.A(n_1945),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2155),
.B(n_943),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_1929),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2057),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_SL g2343 ( 
.A(n_1987),
.B(n_795),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_1933),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2057),
.Y(n_2345)
);

OAI22xp5_ASAP7_75t_SL g2346 ( 
.A1(n_1962),
.A2(n_1684),
.B1(n_1720),
.B2(n_1681),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2059),
.Y(n_2347)
);

AND2x4_ASAP7_75t_L g2348 ( 
.A(n_1946),
.B(n_2164),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2059),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_1933),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2077),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_1941),
.Y(n_2352)
);

OAI22xp5_ASAP7_75t_SL g2353 ( 
.A1(n_1962),
.A2(n_1720),
.B1(n_1722),
.B2(n_1684),
.Y(n_2353)
);

INVxp67_ASAP7_75t_L g2354 ( 
.A(n_2107),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2077),
.Y(n_2355)
);

AO22x1_ASAP7_75t_SL g2356 ( 
.A1(n_2157),
.A2(n_1726),
.B1(n_1730),
.B2(n_1722),
.Y(n_2356)
);

HB1xp67_ASAP7_75t_L g2357 ( 
.A(n_2204),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2216),
.B(n_951),
.Y(n_2358)
);

INVx3_ASAP7_75t_L g2359 ( 
.A(n_2042),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2078),
.Y(n_2360)
);

NAND2xp33_ASAP7_75t_SL g2361 ( 
.A(n_2214),
.B(n_953),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2078),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2084),
.Y(n_2363)
);

HB1xp67_ASAP7_75t_L g2364 ( 
.A(n_2205),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_2228),
.B(n_1456),
.Y(n_2365)
);

HB1xp67_ASAP7_75t_L g2366 ( 
.A(n_2227),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_1941),
.Y(n_2367)
);

INVx3_ASAP7_75t_L g2368 ( 
.A(n_2042),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_1943),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2084),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2131),
.B(n_953),
.Y(n_2371)
);

NAND2x1p5_ASAP7_75t_L g2372 ( 
.A(n_1960),
.B(n_1209),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2228),
.B(n_1458),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2109),
.Y(n_2374)
);

BUFx6f_ASAP7_75t_L g2375 ( 
.A(n_1945),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_1943),
.Y(n_2376)
);

NOR2xp33_ASAP7_75t_SL g2377 ( 
.A(n_1932),
.B(n_2199),
.Y(n_2377)
);

BUFx6f_ASAP7_75t_SL g2378 ( 
.A(n_2161),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2109),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_1944),
.Y(n_2380)
);

AOI22xp5_ASAP7_75t_L g2381 ( 
.A1(n_2225),
.A2(n_781),
.B1(n_783),
.B2(n_776),
.Y(n_2381)
);

AND2x4_ASAP7_75t_L g2382 ( 
.A(n_1946),
.B(n_2164),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2138),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2131),
.B(n_954),
.Y(n_2384)
);

AOI22xp5_ASAP7_75t_L g2385 ( 
.A1(n_2225),
.A2(n_793),
.B1(n_796),
.B2(n_787),
.Y(n_2385)
);

AND2x4_ASAP7_75t_L g2386 ( 
.A(n_1946),
.B(n_2164),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_1944),
.Y(n_2387)
);

OAI22xp5_ASAP7_75t_SL g2388 ( 
.A1(n_1993),
.A2(n_1730),
.B1(n_1746),
.B2(n_1726),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2138),
.Y(n_2389)
);

BUFx6f_ASAP7_75t_L g2390 ( 
.A(n_1951),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_1923),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_SL g2392 ( 
.A(n_1987),
.B(n_2265),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2131),
.B(n_954),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_1925),
.Y(n_2394)
);

HB1xp67_ASAP7_75t_L g2395 ( 
.A(n_2056),
.Y(n_2395)
);

INVx4_ASAP7_75t_L g2396 ( 
.A(n_2119),
.Y(n_2396)
);

BUFx6f_ASAP7_75t_L g2397 ( 
.A(n_1951),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_1926),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_1955),
.Y(n_2399)
);

BUFx6f_ASAP7_75t_L g2400 ( 
.A(n_1951),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_1955),
.Y(n_2401)
);

BUFx2_ASAP7_75t_L g2402 ( 
.A(n_1932),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_1934),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_SL g2404 ( 
.A(n_1987),
.B(n_2265),
.Y(n_2404)
);

HB1xp67_ASAP7_75t_L g2405 ( 
.A(n_2082),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_SL g2406 ( 
.A(n_2265),
.B(n_967),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_1948),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_2242),
.B(n_1462),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_SL g2409 ( 
.A(n_2277),
.B(n_967),
.Y(n_2409)
);

BUFx2_ASAP7_75t_L g2410 ( 
.A(n_1993),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_1961),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_1965),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_SL g2413 ( 
.A(n_2277),
.B(n_967),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_1957),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_1969),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_SL g2416 ( 
.A(n_2277),
.B(n_967),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_1957),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_1972),
.Y(n_2418)
);

AND2x4_ASAP7_75t_L g2419 ( 
.A(n_2286),
.B(n_1463),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_1971),
.Y(n_2420)
);

NOR2xp33_ASAP7_75t_L g2421 ( 
.A(n_1940),
.B(n_798),
.Y(n_2421)
);

OAI22xp5_ASAP7_75t_L g2422 ( 
.A1(n_1959),
.A2(n_806),
.B1(n_808),
.B2(n_805),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_1971),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_1979),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_1981),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_1983),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_1979),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_1935),
.Y(n_2428)
);

INVx3_ASAP7_75t_L g2429 ( 
.A(n_2042),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_SL g2430 ( 
.A(n_2278),
.B(n_1021),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_1986),
.Y(n_2431)
);

BUFx2_ASAP7_75t_L g2432 ( 
.A(n_2312),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_1990),
.Y(n_2433)
);

NOR2xp33_ASAP7_75t_L g2434 ( 
.A(n_2112),
.B(n_809),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_1992),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_SL g2436 ( 
.A(n_2278),
.B(n_1021),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_1935),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_1935),
.Y(n_2438)
);

NAND2x1p5_ASAP7_75t_L g2439 ( 
.A(n_1960),
.B(n_1210),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_1938),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_1938),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_1938),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2001),
.Y(n_2443)
);

BUFx6f_ASAP7_75t_L g2444 ( 
.A(n_1951),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2002),
.Y(n_2445)
);

INVx5_ASAP7_75t_L g2446 ( 
.A(n_1991),
.Y(n_2446)
);

BUFx2_ASAP7_75t_L g2447 ( 
.A(n_2312),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_1949),
.Y(n_2448)
);

AND2x4_ASAP7_75t_L g2449 ( 
.A(n_2286),
.B(n_1467),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_1949),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2085),
.B(n_959),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_SL g2452 ( 
.A(n_2278),
.B(n_1021),
.Y(n_2452)
);

NAND2xp33_ASAP7_75t_SL g2453 ( 
.A(n_2214),
.B(n_959),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2085),
.B(n_2076),
.Y(n_2454)
);

HB1xp67_ASAP7_75t_L g2455 ( 
.A(n_2236),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_SL g2456 ( 
.A(n_2290),
.B(n_1021),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2013),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_1949),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2018),
.Y(n_2459)
);

AOI22xp5_ASAP7_75t_L g2460 ( 
.A1(n_2225),
.A2(n_818),
.B1(n_819),
.B2(n_816),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2076),
.B(n_960),
.Y(n_2461)
);

CKINVDCx5p33_ASAP7_75t_R g2462 ( 
.A(n_1937),
.Y(n_2462)
);

NOR2xp33_ASAP7_75t_SL g2463 ( 
.A(n_2009),
.B(n_1746),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_1966),
.Y(n_2464)
);

BUFx8_ASAP7_75t_L g2465 ( 
.A(n_2289),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_SL g2466 ( 
.A(n_2290),
.B(n_1053),
.Y(n_2466)
);

INVx1_ASAP7_75t_SL g2467 ( 
.A(n_1995),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2242),
.B(n_1468),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_1966),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2019),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2021),
.Y(n_2471)
);

OAI22xp5_ASAP7_75t_L g2472 ( 
.A1(n_1924),
.A2(n_827),
.B1(n_828),
.B2(n_822),
.Y(n_2472)
);

AND2x4_ASAP7_75t_L g2473 ( 
.A(n_2286),
.B(n_1470),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_1966),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2022),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2024),
.Y(n_2476)
);

NAND2xp33_ASAP7_75t_SL g2477 ( 
.A(n_2214),
.B(n_960),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2025),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_1976),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_SL g2480 ( 
.A(n_2290),
.B(n_1053),
.Y(n_2480)
);

BUFx2_ASAP7_75t_L g2481 ( 
.A(n_1995),
.Y(n_2481)
);

NAND2x1_ASAP7_75t_L g2482 ( 
.A(n_1976),
.B(n_1213),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_1976),
.Y(n_2483)
);

AND2x2_ASAP7_75t_L g2484 ( 
.A(n_2268),
.B(n_1471),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_1978),
.Y(n_2485)
);

INVx3_ASAP7_75t_L g2486 ( 
.A(n_2042),
.Y(n_2486)
);

INVx1_ASAP7_75t_SL g2487 ( 
.A(n_2003),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_1978),
.Y(n_2488)
);

OAI22xp5_ASAP7_75t_SL g2489 ( 
.A1(n_2003),
.A2(n_1766),
.B1(n_1780),
.B2(n_1762),
.Y(n_2489)
);

AND3x1_ASAP7_75t_L g2490 ( 
.A(n_2306),
.B(n_962),
.C(n_961),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_SL g2491 ( 
.A(n_2298),
.B(n_2282),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_SL g2492 ( 
.A(n_2298),
.B(n_1053),
.Y(n_2492)
);

AND2x4_ASAP7_75t_L g2493 ( 
.A(n_1964),
.B(n_1473),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2031),
.Y(n_2494)
);

BUFx6f_ASAP7_75t_L g2495 ( 
.A(n_1958),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2033),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2124),
.B(n_961),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_SL g2498 ( 
.A(n_2298),
.B(n_1053),
.Y(n_2498)
);

BUFx8_ASAP7_75t_L g2499 ( 
.A(n_2125),
.Y(n_2499)
);

INVx3_ASAP7_75t_L g2500 ( 
.A(n_1927),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_1978),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_SL g2502 ( 
.A(n_2282),
.B(n_1110),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_1989),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_1989),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2034),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2041),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_1997),
.Y(n_2507)
);

NOR2x1_ASAP7_75t_L g2508 ( 
.A(n_2262),
.B(n_1475),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_1997),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2043),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2049),
.Y(n_2511)
);

NAND2xp33_ASAP7_75t_SL g2512 ( 
.A(n_2237),
.B(n_962),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2052),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2054),
.Y(n_2514)
);

OAI22xp5_ASAP7_75t_SL g2515 ( 
.A1(n_2012),
.A2(n_1766),
.B1(n_1780),
.B2(n_1762),
.Y(n_2515)
);

BUFx6f_ASAP7_75t_L g2516 ( 
.A(n_1958),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2060),
.Y(n_2517)
);

AOI22xp5_ASAP7_75t_L g2518 ( 
.A1(n_2225),
.A2(n_830),
.B1(n_840),
.B2(n_829),
.Y(n_2518)
);

INVxp67_ASAP7_75t_L g2519 ( 
.A(n_2309),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2124),
.B(n_975),
.Y(n_2520)
);

BUFx2_ASAP7_75t_L g2521 ( 
.A(n_2012),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2064),
.Y(n_2522)
);

INVx3_ASAP7_75t_L g2523 ( 
.A(n_1927),
.Y(n_2523)
);

INVx3_ASAP7_75t_L g2524 ( 
.A(n_1927),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_2124),
.B(n_975),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2006),
.Y(n_2526)
);

INVx1_ASAP7_75t_SL g2527 ( 
.A(n_2016),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2006),
.Y(n_2528)
);

BUFx2_ASAP7_75t_L g2529 ( 
.A(n_2316),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2086),
.Y(n_2530)
);

INVx3_ASAP7_75t_L g2531 ( 
.A(n_1931),
.Y(n_2531)
);

AND3x1_ASAP7_75t_L g2532 ( 
.A(n_2306),
.B(n_2285),
.C(n_2284),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2088),
.Y(n_2533)
);

AND2x2_ASAP7_75t_L g2534 ( 
.A(n_2268),
.B(n_1482),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2095),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2141),
.B(n_981),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_2141),
.B(n_981),
.Y(n_2537)
);

OAI22xp5_ASAP7_75t_SL g2538 ( 
.A1(n_2016),
.A2(n_1801),
.B1(n_1803),
.B2(n_1793),
.Y(n_2538)
);

INVx3_ASAP7_75t_L g2539 ( 
.A(n_1931),
.Y(n_2539)
);

NAND2xp33_ASAP7_75t_SL g2540 ( 
.A(n_2237),
.B(n_982),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2097),
.Y(n_2541)
);

BUFx6f_ASAP7_75t_L g2542 ( 
.A(n_1958),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2023),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2141),
.B(n_982),
.Y(n_2544)
);

CKINVDCx5p33_ASAP7_75t_R g2545 ( 
.A(n_1937),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_SL g2546 ( 
.A(n_2284),
.B(n_1110),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2098),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2101),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2023),
.Y(n_2549)
);

OAI22xp5_ASAP7_75t_L g2550 ( 
.A1(n_1924),
.A2(n_842),
.B1(n_843),
.B2(n_841),
.Y(n_2550)
);

NOR2xp33_ASAP7_75t_SL g2551 ( 
.A(n_2009),
.B(n_1793),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2111),
.Y(n_2552)
);

AND2x6_ASAP7_75t_L g2553 ( 
.A(n_2236),
.B(n_985),
.Y(n_2553)
);

BUFx6f_ASAP7_75t_L g2554 ( 
.A(n_1958),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2037),
.Y(n_2555)
);

BUFx6f_ASAP7_75t_L g2556 ( 
.A(n_1963),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2116),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2117),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2120),
.Y(n_2559)
);

AOI22xp5_ASAP7_75t_L g2560 ( 
.A1(n_2225),
.A2(n_846),
.B1(n_847),
.B2(n_844),
.Y(n_2560)
);

AOI22xp5_ASAP7_75t_L g2561 ( 
.A1(n_2293),
.A2(n_849),
.B1(n_850),
.B2(n_848),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2121),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2037),
.Y(n_2563)
);

AND2x4_ASAP7_75t_L g2564 ( 
.A(n_1964),
.B(n_1485),
.Y(n_2564)
);

AND2x4_ASAP7_75t_L g2565 ( 
.A(n_1998),
.B(n_1487),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2126),
.Y(n_2566)
);

BUFx6f_ASAP7_75t_L g2567 ( 
.A(n_1963),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2127),
.Y(n_2568)
);

OAI22xp5_ASAP7_75t_L g2569 ( 
.A1(n_2045),
.A2(n_854),
.B1(n_856),
.B2(n_852),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2129),
.Y(n_2570)
);

INVx3_ASAP7_75t_L g2571 ( 
.A(n_1931),
.Y(n_2571)
);

BUFx6f_ASAP7_75t_L g2572 ( 
.A(n_1963),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_SL g2573 ( 
.A(n_2285),
.B(n_1110),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2133),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2140),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2149),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2151),
.Y(n_2577)
);

BUFx6f_ASAP7_75t_L g2578 ( 
.A(n_1963),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2040),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2147),
.Y(n_2580)
);

INVxp67_ASAP7_75t_L g2581 ( 
.A(n_2311),
.Y(n_2581)
);

BUFx6f_ASAP7_75t_L g2582 ( 
.A(n_1968),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2147),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2147),
.Y(n_2584)
);

AOI22xp5_ASAP7_75t_L g2585 ( 
.A1(n_2293),
.A2(n_859),
.B1(n_861),
.B2(n_857),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2050),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2050),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2040),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_SL g2589 ( 
.A(n_2161),
.B(n_1110),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2123),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2123),
.Y(n_2591)
);

INVx2_ASAP7_75t_L g2592 ( 
.A(n_2051),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2051),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2051),
.Y(n_2594)
);

BUFx6f_ASAP7_75t_L g2595 ( 
.A(n_1968),
.Y(n_2595)
);

HB1xp67_ASAP7_75t_L g2596 ( 
.A(n_2236),
.Y(n_2596)
);

AOI22xp5_ASAP7_75t_L g2597 ( 
.A1(n_2293),
.A2(n_863),
.B1(n_864),
.B2(n_862),
.Y(n_2597)
);

NOR2x1_ASAP7_75t_L g2598 ( 
.A(n_2237),
.B(n_1488),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2061),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2061),
.Y(n_2600)
);

INVx3_ASAP7_75t_L g2601 ( 
.A(n_1999),
.Y(n_2601)
);

INVx1_ASAP7_75t_SL g2602 ( 
.A(n_2030),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2061),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2080),
.Y(n_2604)
);

OAI22xp5_ASAP7_75t_SL g2605 ( 
.A1(n_2030),
.A2(n_1803),
.B1(n_1811),
.B2(n_1801),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2080),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2080),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_SL g2608 ( 
.A(n_2161),
.B(n_1118),
.Y(n_2608)
);

BUFx6f_ASAP7_75t_SL g2609 ( 
.A(n_2161),
.Y(n_2609)
);

AND2x2_ASAP7_75t_L g2610 ( 
.A(n_2173),
.B(n_1489),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2091),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2091),
.Y(n_2612)
);

INVxp67_ASAP7_75t_L g2613 ( 
.A(n_2173),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_2091),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2108),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_1920),
.B(n_985),
.Y(n_2616)
);

BUFx8_ASAP7_75t_L g2617 ( 
.A(n_2174),
.Y(n_2617)
);

NAND2xp33_ASAP7_75t_SL g2618 ( 
.A(n_2179),
.B(n_986),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2108),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2108),
.Y(n_2620)
);

BUFx6f_ASAP7_75t_L g2621 ( 
.A(n_1968),
.Y(n_2621)
);

CKINVDCx20_ASAP7_75t_R g2622 ( 
.A(n_2053),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_1928),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_1928),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2093),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2092),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2092),
.Y(n_2627)
);

AOI22xp5_ASAP7_75t_L g2628 ( 
.A1(n_2293),
.A2(n_867),
.B1(n_871),
.B2(n_865),
.Y(n_2628)
);

NAND3xp33_ASAP7_75t_L g2629 ( 
.A(n_1950),
.B(n_873),
.C(n_872),
.Y(n_2629)
);

INVx1_ASAP7_75t_SL g2630 ( 
.A(n_2053),
.Y(n_2630)
);

INVx3_ASAP7_75t_L g2631 ( 
.A(n_1999),
.Y(n_2631)
);

INVx3_ASAP7_75t_L g2632 ( 
.A(n_1999),
.Y(n_2632)
);

NAND2xp33_ASAP7_75t_SL g2633 ( 
.A(n_2179),
.B(n_986),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2096),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2096),
.Y(n_2635)
);

AND2x4_ASAP7_75t_L g2636 ( 
.A(n_1998),
.B(n_1493),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2132),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_SL g2638 ( 
.A(n_2179),
.B(n_1118),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_2093),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2132),
.Y(n_2640)
);

INVx3_ASAP7_75t_L g2641 ( 
.A(n_2000),
.Y(n_2641)
);

HB1xp67_ASAP7_75t_L g2642 ( 
.A(n_2244),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2119),
.Y(n_2643)
);

AND2x2_ASAP7_75t_L g2644 ( 
.A(n_2287),
.B(n_1497),
.Y(n_2644)
);

AND2x2_ASAP7_75t_L g2645 ( 
.A(n_2287),
.B(n_1501),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_2119),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2048),
.Y(n_2647)
);

BUFx6f_ASAP7_75t_L g2648 ( 
.A(n_1968),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_2119),
.Y(n_2649)
);

AOI22xp33_ASAP7_75t_SL g2650 ( 
.A1(n_2195),
.A2(n_1811),
.B1(n_1833),
.B2(n_1820),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_1922),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2137),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2070),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_1952),
.B(n_988),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2070),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2137),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2070),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2026),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2137),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2137),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2143),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_SL g2662 ( 
.A(n_2179),
.B(n_1118),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2143),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2143),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2143),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2066),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_SL g2667 ( 
.A(n_2183),
.B(n_1118),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2066),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_SL g2669 ( 
.A(n_2183),
.B(n_876),
.Y(n_2669)
);

INVxp67_ASAP7_75t_L g2670 ( 
.A(n_2209),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_2000),
.Y(n_2671)
);

NAND2xp33_ASAP7_75t_SL g2672 ( 
.A(n_2183),
.B(n_2198),
.Y(n_2672)
);

BUFx6f_ASAP7_75t_L g2673 ( 
.A(n_1982),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2105),
.Y(n_2674)
);

HB1xp67_ASAP7_75t_L g2675 ( 
.A(n_2244),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2105),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2106),
.Y(n_2677)
);

CKINVDCx5p33_ASAP7_75t_R g2678 ( 
.A(n_1953),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2106),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2156),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2158),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2145),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_SL g2683 ( 
.A(n_2183),
.B(n_879),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_2000),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2145),
.Y(n_2685)
);

AND2x6_ASAP7_75t_L g2686 ( 
.A(n_2244),
.B(n_988),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2145),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2014),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2148),
.Y(n_2689)
);

INVx3_ASAP7_75t_L g2690 ( 
.A(n_2014),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2148),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2148),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2058),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2058),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2058),
.Y(n_2695)
);

NAND2xp33_ASAP7_75t_SL g2696 ( 
.A(n_2198),
.B(n_991),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_SL g2697 ( 
.A(n_2198),
.B(n_880),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2152),
.B(n_2154),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2014),
.Y(n_2699)
);

INVx3_ASAP7_75t_L g2700 ( 
.A(n_2029),
.Y(n_2700)
);

OAI22xp5_ASAP7_75t_SL g2701 ( 
.A1(n_2089),
.A2(n_1833),
.B1(n_1834),
.B2(n_1820),
.Y(n_2701)
);

OAI22xp5_ASAP7_75t_L g2702 ( 
.A1(n_2015),
.A2(n_883),
.B1(n_884),
.B2(n_881),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_1952),
.B(n_991),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2063),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2063),
.Y(n_2705)
);

INVx3_ASAP7_75t_L g2706 ( 
.A(n_2029),
.Y(n_2706)
);

BUFx3_ASAP7_75t_L g2707 ( 
.A(n_2176),
.Y(n_2707)
);

BUFx6f_ASAP7_75t_L g2708 ( 
.A(n_1982),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2029),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2063),
.Y(n_2710)
);

INVx2_ASAP7_75t_L g2711 ( 
.A(n_2036),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2036),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2063),
.Y(n_2713)
);

OA21x2_ASAP7_75t_L g2714 ( 
.A1(n_2069),
.A2(n_1224),
.B(n_1222),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2036),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2067),
.Y(n_2716)
);

NAND2xp33_ASAP7_75t_SL g2717 ( 
.A(n_2198),
.B(n_996),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2212),
.Y(n_2718)
);

HB1xp67_ASAP7_75t_L g2719 ( 
.A(n_2250),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2067),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2067),
.Y(n_2721)
);

HB1xp67_ASAP7_75t_L g2722 ( 
.A(n_2250),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2067),
.Y(n_2723)
);

INVx3_ASAP7_75t_L g2724 ( 
.A(n_2212),
.Y(n_2724)
);

CKINVDCx8_ASAP7_75t_R g2725 ( 
.A(n_2130),
.Y(n_2725)
);

OAI22xp5_ASAP7_75t_SL g2726 ( 
.A1(n_2089),
.A2(n_1839),
.B1(n_1840),
.B2(n_1834),
.Y(n_2726)
);

AND2x2_ASAP7_75t_L g2727 ( 
.A(n_2152),
.B(n_2154),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_2212),
.Y(n_2728)
);

INVx2_ASAP7_75t_L g2729 ( 
.A(n_2071),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2071),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2071),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2071),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2072),
.Y(n_2733)
);

AND2x2_ASAP7_75t_L g2734 ( 
.A(n_2165),
.B(n_1504),
.Y(n_2734)
);

BUFx6f_ASAP7_75t_SL g2735 ( 
.A(n_2219),
.Y(n_2735)
);

NOR2xp33_ASAP7_75t_L g2736 ( 
.A(n_2519),
.B(n_2581),
.Y(n_2736)
);

BUFx6f_ASAP7_75t_L g2737 ( 
.A(n_2707),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_2327),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2327),
.Y(n_2739)
);

BUFx10_ASAP7_75t_L g2740 ( 
.A(n_2378),
.Y(n_2740)
);

AOI22xp33_ASAP7_75t_L g2741 ( 
.A1(n_2454),
.A2(n_2293),
.B1(n_2159),
.B2(n_2182),
.Y(n_2741)
);

INVx1_ASAP7_75t_SL g2742 ( 
.A(n_2467),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2653),
.Y(n_2743)
);

BUFx10_ASAP7_75t_L g2744 ( 
.A(n_2378),
.Y(n_2744)
);

NOR2x1p5_ASAP7_75t_L g2745 ( 
.A(n_2462),
.B(n_1974),
.Y(n_2745)
);

BUFx6f_ASAP7_75t_L g2746 ( 
.A(n_2707),
.Y(n_2746)
);

BUFx3_ASAP7_75t_L g2747 ( 
.A(n_2725),
.Y(n_2747)
);

INVx4_ASAP7_75t_L g2748 ( 
.A(n_2378),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2330),
.Y(n_2749)
);

NOR2xp33_ASAP7_75t_L g2750 ( 
.A(n_2348),
.B(n_1977),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2658),
.B(n_2647),
.Y(n_2751)
);

NOR2xp33_ASAP7_75t_L g2752 ( 
.A(n_2348),
.B(n_1977),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2698),
.B(n_2727),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2655),
.Y(n_2754)
);

INVx4_ASAP7_75t_L g2755 ( 
.A(n_2609),
.Y(n_2755)
);

INVx3_ASAP7_75t_L g2756 ( 
.A(n_2396),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2657),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2433),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2435),
.Y(n_2759)
);

AND2x4_ASAP7_75t_L g2760 ( 
.A(n_2348),
.B(n_2219),
.Y(n_2760)
);

INVx2_ASAP7_75t_L g2761 ( 
.A(n_2330),
.Y(n_2761)
);

NOR2xp33_ASAP7_75t_L g2762 ( 
.A(n_2382),
.B(n_2246),
.Y(n_2762)
);

AND2x4_ASAP7_75t_L g2763 ( 
.A(n_2382),
.B(n_2219),
.Y(n_2763)
);

OR2x6_ASAP7_75t_L g2764 ( 
.A(n_2356),
.B(n_2176),
.Y(n_2764)
);

AOI22xp33_ASAP7_75t_L g2765 ( 
.A1(n_2382),
.A2(n_2293),
.B1(n_2159),
.B2(n_2182),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2443),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2698),
.B(n_2160),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_SL g2768 ( 
.A(n_2377),
.B(n_2219),
.Y(n_2768)
);

INVx2_ASAP7_75t_L g2769 ( 
.A(n_2332),
.Y(n_2769)
);

INVxp67_ASAP7_75t_L g2770 ( 
.A(n_2357),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2332),
.Y(n_2771)
);

AND2x2_ASAP7_75t_L g2772 ( 
.A(n_2727),
.B(n_2301),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2445),
.Y(n_2773)
);

NOR2xp33_ASAP7_75t_L g2774 ( 
.A(n_2386),
.B(n_2246),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2644),
.B(n_2160),
.Y(n_2775)
);

AND2x2_ASAP7_75t_L g2776 ( 
.A(n_2455),
.B(n_2301),
.Y(n_2776)
);

AND2x4_ASAP7_75t_L g2777 ( 
.A(n_2386),
.B(n_2226),
.Y(n_2777)
);

XOR2x2_ASAP7_75t_L g2778 ( 
.A(n_2346),
.B(n_1942),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2457),
.Y(n_2779)
);

BUFx3_ASAP7_75t_L g2780 ( 
.A(n_2725),
.Y(n_2780)
);

BUFx6f_ASAP7_75t_L g2781 ( 
.A(n_2324),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2459),
.Y(n_2782)
);

NOR2xp33_ASAP7_75t_L g2783 ( 
.A(n_2386),
.B(n_2297),
.Y(n_2783)
);

BUFx3_ASAP7_75t_L g2784 ( 
.A(n_2465),
.Y(n_2784)
);

INVx4_ASAP7_75t_L g2785 ( 
.A(n_2609),
.Y(n_2785)
);

NOR2xp33_ASAP7_75t_L g2786 ( 
.A(n_2331),
.B(n_2491),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2470),
.Y(n_2787)
);

AND2x6_ASAP7_75t_L g2788 ( 
.A(n_2718),
.B(n_2728),
.Y(n_2788)
);

INVx4_ASAP7_75t_L g2789 ( 
.A(n_2609),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2644),
.B(n_2160),
.Y(n_2790)
);

OA22x2_ASAP7_75t_L g2791 ( 
.A1(n_2596),
.A2(n_2135),
.B1(n_2217),
.B2(n_2229),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_2645),
.B(n_1952),
.Y(n_2792)
);

INVx4_ASAP7_75t_L g2793 ( 
.A(n_2735),
.Y(n_2793)
);

AND2x6_ASAP7_75t_L g2794 ( 
.A(n_2693),
.B(n_2226),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2471),
.Y(n_2795)
);

INVx4_ASAP7_75t_L g2796 ( 
.A(n_2735),
.Y(n_2796)
);

INVx4_ASAP7_75t_L g2797 ( 
.A(n_2735),
.Y(n_2797)
);

NOR2xp33_ASAP7_75t_L g2798 ( 
.A(n_2491),
.B(n_2297),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2645),
.B(n_2150),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2475),
.Y(n_2800)
);

INVx2_ASAP7_75t_L g2801 ( 
.A(n_2341),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_L g2802 ( 
.A(n_2592),
.B(n_1975),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2476),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2478),
.Y(n_2804)
);

NOR2xp33_ASAP7_75t_L g2805 ( 
.A(n_2333),
.B(n_2297),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2494),
.Y(n_2806)
);

CKINVDCx14_ASAP7_75t_R g2807 ( 
.A(n_2353),
.Y(n_2807)
);

INVx3_ASAP7_75t_L g2808 ( 
.A(n_2396),
.Y(n_2808)
);

NOR2x1p5_ASAP7_75t_L g2809 ( 
.A(n_2462),
.B(n_1974),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2496),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2592),
.B(n_1975),
.Y(n_2811)
);

INVx1_ASAP7_75t_SL g2812 ( 
.A(n_2487),
.Y(n_2812)
);

OR2x2_ASAP7_75t_L g2813 ( 
.A(n_2527),
.B(n_2074),
.Y(n_2813)
);

NOR2xp33_ASAP7_75t_L g2814 ( 
.A(n_2333),
.B(n_2068),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2505),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2600),
.B(n_2068),
.Y(n_2816)
);

NOR2xp33_ASAP7_75t_L g2817 ( 
.A(n_2421),
.B(n_2068),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2506),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2510),
.Y(n_2819)
);

CKINVDCx16_ASAP7_75t_R g2820 ( 
.A(n_2622),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2511),
.Y(n_2821)
);

AND2x4_ASAP7_75t_L g2822 ( 
.A(n_2694),
.B(n_2226),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2341),
.Y(n_2823)
);

NOR2xp33_ASAP7_75t_L g2824 ( 
.A(n_2421),
.B(n_2191),
.Y(n_2824)
);

NOR2xp33_ASAP7_75t_L g2825 ( 
.A(n_2392),
.B(n_2191),
.Y(n_2825)
);

INVx2_ASAP7_75t_L g2826 ( 
.A(n_2344),
.Y(n_2826)
);

NOR2xp33_ASAP7_75t_L g2827 ( 
.A(n_2392),
.B(n_2404),
.Y(n_2827)
);

BUFx6f_ASAP7_75t_L g2828 ( 
.A(n_2324),
.Y(n_2828)
);

BUFx2_ASAP7_75t_L g2829 ( 
.A(n_2622),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2600),
.B(n_2165),
.Y(n_2830)
);

INVx4_ASAP7_75t_L g2831 ( 
.A(n_2545),
.Y(n_2831)
);

NOR2xp33_ASAP7_75t_L g2832 ( 
.A(n_2404),
.B(n_2191),
.Y(n_2832)
);

INVx3_ASAP7_75t_L g2833 ( 
.A(n_2396),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2513),
.Y(n_2834)
);

AND2x2_ASAP7_75t_L g2835 ( 
.A(n_2642),
.B(n_2233),
.Y(n_2835)
);

AND2x4_ASAP7_75t_L g2836 ( 
.A(n_2695),
.B(n_2226),
.Y(n_2836)
);

NOR2xp33_ASAP7_75t_L g2837 ( 
.A(n_2675),
.B(n_2207),
.Y(n_2837)
);

BUFx6f_ASAP7_75t_L g2838 ( 
.A(n_2324),
.Y(n_2838)
);

INVx4_ASAP7_75t_L g2839 ( 
.A(n_2545),
.Y(n_2839)
);

INVx2_ASAP7_75t_SL g2840 ( 
.A(n_2325),
.Y(n_2840)
);

CKINVDCx6p67_ASAP7_75t_R g2841 ( 
.A(n_2402),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2606),
.B(n_2128),
.Y(n_2842)
);

CKINVDCx20_ASAP7_75t_R g2843 ( 
.A(n_2678),
.Y(n_2843)
);

INVx2_ASAP7_75t_SL g2844 ( 
.A(n_2325),
.Y(n_2844)
);

INVx5_ASAP7_75t_L g2845 ( 
.A(n_2324),
.Y(n_2845)
);

INVx2_ASAP7_75t_SL g2846 ( 
.A(n_2465),
.Y(n_2846)
);

AND2x2_ASAP7_75t_L g2847 ( 
.A(n_2719),
.B(n_2250),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2606),
.B(n_1954),
.Y(n_2848)
);

AND2x4_ASAP7_75t_L g2849 ( 
.A(n_2682),
.B(n_2245),
.Y(n_2849)
);

AOI22xp5_ASAP7_75t_L g2850 ( 
.A1(n_2553),
.A2(n_2122),
.B1(n_2153),
.B2(n_2146),
.Y(n_2850)
);

BUFx2_ASAP7_75t_L g2851 ( 
.A(n_2328),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_SL g2852 ( 
.A(n_2672),
.B(n_2245),
.Y(n_2852)
);

BUFx10_ASAP7_75t_L g2853 ( 
.A(n_2678),
.Y(n_2853)
);

INVx2_ASAP7_75t_L g2854 ( 
.A(n_2344),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2514),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2517),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2350),
.Y(n_2857)
);

AND2x4_ASAP7_75t_L g2858 ( 
.A(n_2685),
.B(n_2245),
.Y(n_2858)
);

NAND2x1p5_ASAP7_75t_L g2859 ( 
.A(n_2446),
.B(n_2245),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2522),
.Y(n_2860)
);

BUFx4f_ASAP7_75t_L g2861 ( 
.A(n_2553),
.Y(n_2861)
);

INVx2_ASAP7_75t_L g2862 ( 
.A(n_2350),
.Y(n_2862)
);

INVx2_ASAP7_75t_L g2863 ( 
.A(n_2352),
.Y(n_2863)
);

BUFx6f_ASAP7_75t_L g2864 ( 
.A(n_2334),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2530),
.Y(n_2865)
);

INVx2_ASAP7_75t_SL g2866 ( 
.A(n_2465),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2352),
.Y(n_2867)
);

AOI22xp33_ASAP7_75t_L g2868 ( 
.A1(n_2553),
.A2(n_2182),
.B1(n_2230),
.B2(n_2195),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2533),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2535),
.Y(n_2870)
);

AND2x2_ASAP7_75t_L g2871 ( 
.A(n_2722),
.B(n_2146),
.Y(n_2871)
);

AND2x2_ASAP7_75t_L g2872 ( 
.A(n_2610),
.B(n_2153),
.Y(n_2872)
);

CKINVDCx16_ASAP7_75t_R g2873 ( 
.A(n_2388),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2541),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2547),
.Y(n_2875)
);

AND2x6_ASAP7_75t_L g2876 ( 
.A(n_2687),
.B(n_2252),
.Y(n_2876)
);

BUFx6f_ASAP7_75t_L g2877 ( 
.A(n_2334),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2548),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2552),
.Y(n_2879)
);

CKINVDCx20_ASAP7_75t_R g2880 ( 
.A(n_2499),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2367),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2557),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2558),
.Y(n_2883)
);

INVx4_ASAP7_75t_L g2884 ( 
.A(n_2446),
.Y(n_2884)
);

AND2x4_ASAP7_75t_L g2885 ( 
.A(n_2689),
.B(n_2252),
.Y(n_2885)
);

BUFx6f_ASAP7_75t_L g2886 ( 
.A(n_2334),
.Y(n_2886)
);

BUFx3_ASAP7_75t_L g2887 ( 
.A(n_2499),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2559),
.Y(n_2888)
);

CKINVDCx5p33_ASAP7_75t_R g2889 ( 
.A(n_2499),
.Y(n_2889)
);

INVx3_ASAP7_75t_L g2890 ( 
.A(n_2334),
.Y(n_2890)
);

AOI22xp5_ASAP7_75t_L g2891 ( 
.A1(n_2553),
.A2(n_2122),
.B1(n_2171),
.B2(n_2170),
.Y(n_2891)
);

AND2x6_ASAP7_75t_L g2892 ( 
.A(n_2691),
.B(n_2692),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2562),
.Y(n_2893)
);

CKINVDCx5p33_ASAP7_75t_R g2894 ( 
.A(n_2617),
.Y(n_2894)
);

NAND3xp33_ASAP7_75t_L g2895 ( 
.A(n_2434),
.B(n_2280),
.C(n_2203),
.Y(n_2895)
);

INVx1_ASAP7_75t_SL g2896 ( 
.A(n_2602),
.Y(n_2896)
);

CKINVDCx5p33_ASAP7_75t_R g2897 ( 
.A(n_2617),
.Y(n_2897)
);

INVxp67_ASAP7_75t_L g2898 ( 
.A(n_2364),
.Y(n_2898)
);

BUFx6f_ASAP7_75t_L g2899 ( 
.A(n_2339),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2607),
.B(n_2614),
.Y(n_2900)
);

OR2x6_ASAP7_75t_SL g2901 ( 
.A(n_2629),
.B(n_2170),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2367),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2566),
.Y(n_2903)
);

INVx4_ASAP7_75t_L g2904 ( 
.A(n_2446),
.Y(n_2904)
);

OAI22xp33_ASAP7_75t_L g2905 ( 
.A1(n_2358),
.A2(n_2113),
.B1(n_2102),
.B2(n_2074),
.Y(n_2905)
);

AND2x2_ASAP7_75t_L g2906 ( 
.A(n_2610),
.B(n_2171),
.Y(n_2906)
);

INVx2_ASAP7_75t_L g2907 ( 
.A(n_2369),
.Y(n_2907)
);

NOR2xp33_ASAP7_75t_L g2908 ( 
.A(n_2434),
.B(n_2207),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2568),
.Y(n_2909)
);

NAND2x1p5_ASAP7_75t_L g2910 ( 
.A(n_2446),
.B(n_2252),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2369),
.Y(n_2911)
);

CKINVDCx5p33_ASAP7_75t_R g2912 ( 
.A(n_2617),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_SL g2913 ( 
.A(n_2672),
.B(n_2252),
.Y(n_2913)
);

NOR2xp33_ASAP7_75t_L g2914 ( 
.A(n_2613),
.B(n_2207),
.Y(n_2914)
);

AO21x1_ASAP7_75t_L g2915 ( 
.A1(n_2329),
.A2(n_2069),
.B(n_2008),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_SL g2916 ( 
.A(n_2419),
.B(n_2263),
.Y(n_2916)
);

NAND3x1_ASAP7_75t_L g2917 ( 
.A(n_2489),
.B(n_2318),
.C(n_2315),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2570),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2574),
.Y(n_2919)
);

AND2x6_ASAP7_75t_L g2920 ( 
.A(n_2718),
.B(n_2263),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_L g2921 ( 
.A(n_2607),
.B(n_1954),
.Y(n_2921)
);

INVx2_ASAP7_75t_SL g2922 ( 
.A(n_2323),
.Y(n_2922)
);

INVx4_ASAP7_75t_L g2923 ( 
.A(n_2446),
.Y(n_2923)
);

AND2x2_ASAP7_75t_L g2924 ( 
.A(n_2365),
.B(n_2197),
.Y(n_2924)
);

AND2x6_ASAP7_75t_L g2925 ( 
.A(n_2728),
.B(n_2263),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2575),
.Y(n_2926)
);

INVx2_ASAP7_75t_L g2927 ( 
.A(n_2376),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2614),
.B(n_1954),
.Y(n_2928)
);

AND2x4_ASAP7_75t_L g2929 ( 
.A(n_2419),
.B(n_2263),
.Y(n_2929)
);

INVx1_ASAP7_75t_SL g2930 ( 
.A(n_2630),
.Y(n_2930)
);

INVx3_ASAP7_75t_L g2931 ( 
.A(n_2339),
.Y(n_2931)
);

INVxp67_ASAP7_75t_SL g2932 ( 
.A(n_2724),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2376),
.Y(n_2933)
);

OAI21xp33_ASAP7_75t_L g2934 ( 
.A1(n_2381),
.A2(n_2062),
.B(n_2197),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2576),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_SL g2936 ( 
.A(n_2419),
.B(n_2274),
.Y(n_2936)
);

AND2x4_ASAP7_75t_L g2937 ( 
.A(n_2449),
.B(n_2274),
.Y(n_2937)
);

INVx3_ASAP7_75t_L g2938 ( 
.A(n_2339),
.Y(n_2938)
);

AND2x2_ASAP7_75t_L g2939 ( 
.A(n_2365),
.B(n_2213),
.Y(n_2939)
);

INVx2_ASAP7_75t_SL g2940 ( 
.A(n_2410),
.Y(n_2940)
);

BUFx10_ASAP7_75t_L g2941 ( 
.A(n_2449),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2577),
.Y(n_2942)
);

AND2x4_ASAP7_75t_L g2943 ( 
.A(n_2449),
.B(n_2274),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2651),
.Y(n_2944)
);

BUFx2_ASAP7_75t_L g2945 ( 
.A(n_2366),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2391),
.Y(n_2946)
);

INVx2_ASAP7_75t_L g2947 ( 
.A(n_2380),
.Y(n_2947)
);

NOR2xp33_ASAP7_75t_L g2948 ( 
.A(n_2406),
.B(n_2223),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_L g2949 ( 
.A(n_2580),
.B(n_2223),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2380),
.Y(n_2950)
);

AND2x6_ASAP7_75t_L g2951 ( 
.A(n_2643),
.B(n_2274),
.Y(n_2951)
);

NAND2x1p5_ASAP7_75t_L g2952 ( 
.A(n_2359),
.B(n_2303),
.Y(n_2952)
);

INVx2_ASAP7_75t_L g2953 ( 
.A(n_2387),
.Y(n_2953)
);

INVx3_ASAP7_75t_L g2954 ( 
.A(n_2339),
.Y(n_2954)
);

BUFx6f_ASAP7_75t_L g2955 ( 
.A(n_2375),
.Y(n_2955)
);

BUFx6f_ASAP7_75t_L g2956 ( 
.A(n_2375),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_SL g2957 ( 
.A(n_2473),
.B(n_2223),
.Y(n_2957)
);

AND2x6_ASAP7_75t_L g2958 ( 
.A(n_2643),
.B(n_2231),
.Y(n_2958)
);

BUFx2_ASAP7_75t_L g2959 ( 
.A(n_2481),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_SL g2960 ( 
.A(n_2473),
.B(n_2231),
.Y(n_2960)
);

NAND2x1_ASAP7_75t_L g2961 ( 
.A(n_2500),
.B(n_1991),
.Y(n_2961)
);

NOR2xp33_ASAP7_75t_L g2962 ( 
.A(n_2406),
.B(n_2231),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2394),
.Y(n_2963)
);

AOI22xp33_ASAP7_75t_L g2964 ( 
.A1(n_2553),
.A2(n_2182),
.B1(n_2181),
.B2(n_2314),
.Y(n_2964)
);

OR2x2_ASAP7_75t_L g2965 ( 
.A(n_2395),
.B(n_2010),
.Y(n_2965)
);

INVx2_ASAP7_75t_L g2966 ( 
.A(n_2387),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2398),
.Y(n_2967)
);

BUFx3_ASAP7_75t_L g2968 ( 
.A(n_2521),
.Y(n_2968)
);

BUFx2_ASAP7_75t_L g2969 ( 
.A(n_2405),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2403),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_SL g2971 ( 
.A(n_2473),
.B(n_2238),
.Y(n_2971)
);

AND2x4_ASAP7_75t_L g2972 ( 
.A(n_2321),
.B(n_2238),
.Y(n_2972)
);

OR2x2_ASAP7_75t_L g2973 ( 
.A(n_2515),
.B(n_2010),
.Y(n_2973)
);

AO22x2_ASAP7_75t_L g2974 ( 
.A1(n_2650),
.A2(n_2313),
.B1(n_2318),
.B2(n_2315),
.Y(n_2974)
);

AND2x2_ASAP7_75t_L g2975 ( 
.A(n_2373),
.B(n_2213),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2407),
.Y(n_2976)
);

INVx2_ASAP7_75t_L g2977 ( 
.A(n_2399),
.Y(n_2977)
);

NOR2xp33_ASAP7_75t_L g2978 ( 
.A(n_2409),
.B(n_2238),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2411),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2583),
.B(n_2243),
.Y(n_2980)
);

INVx3_ASAP7_75t_L g2981 ( 
.A(n_2375),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2412),
.Y(n_2982)
);

INVx2_ASAP7_75t_L g2983 ( 
.A(n_2399),
.Y(n_2983)
);

INVx4_ASAP7_75t_L g2984 ( 
.A(n_2553),
.Y(n_2984)
);

OR2x2_ASAP7_75t_L g2985 ( 
.A(n_2538),
.B(n_2248),
.Y(n_2985)
);

NOR2xp33_ASAP7_75t_L g2986 ( 
.A(n_2409),
.B(n_2243),
.Y(n_2986)
);

BUFx6f_ASAP7_75t_L g2987 ( 
.A(n_2375),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2415),
.Y(n_2988)
);

INVx3_ASAP7_75t_L g2989 ( 
.A(n_2390),
.Y(n_2989)
);

INVxp67_ASAP7_75t_SL g2990 ( 
.A(n_2724),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2418),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_SL g2992 ( 
.A(n_2532),
.B(n_2243),
.Y(n_2992)
);

INVx3_ASAP7_75t_L g2993 ( 
.A(n_2390),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2401),
.Y(n_2994)
);

BUFx3_ASAP7_75t_L g2995 ( 
.A(n_2432),
.Y(n_2995)
);

INVx5_ASAP7_75t_L g2996 ( 
.A(n_2390),
.Y(n_2996)
);

AND2x2_ASAP7_75t_L g2997 ( 
.A(n_2373),
.B(n_2215),
.Y(n_2997)
);

AND2x6_ASAP7_75t_L g2998 ( 
.A(n_2646),
.B(n_2303),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2425),
.Y(n_2999)
);

INVx3_ASAP7_75t_L g3000 ( 
.A(n_2390),
.Y(n_3000)
);

INVx6_ASAP7_75t_L g3001 ( 
.A(n_2493),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2401),
.Y(n_3002)
);

BUFx10_ASAP7_75t_L g3003 ( 
.A(n_2493),
.Y(n_3003)
);

OR2x2_ASAP7_75t_L g3004 ( 
.A(n_2605),
.B(n_1942),
.Y(n_3004)
);

AOI22xp33_ASAP7_75t_L g3005 ( 
.A1(n_2686),
.A2(n_2182),
.B1(n_2186),
.B2(n_2008),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_L g3006 ( 
.A(n_2584),
.B(n_2142),
.Y(n_3006)
);

HB1xp67_ASAP7_75t_L g3007 ( 
.A(n_2529),
.Y(n_3007)
);

AND2x4_ASAP7_75t_L g3008 ( 
.A(n_2335),
.B(n_2206),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2426),
.Y(n_3009)
);

NOR2xp33_ASAP7_75t_L g3010 ( 
.A(n_2413),
.B(n_2188),
.Y(n_3010)
);

INVx1_ASAP7_75t_SL g3011 ( 
.A(n_2529),
.Y(n_3011)
);

HB1xp67_ASAP7_75t_L g3012 ( 
.A(n_2432),
.Y(n_3012)
);

BUFx6f_ASAP7_75t_L g3013 ( 
.A(n_2397),
.Y(n_3013)
);

HB1xp67_ASAP7_75t_L g3014 ( 
.A(n_2447),
.Y(n_3014)
);

BUFx6f_ASAP7_75t_L g3015 ( 
.A(n_2397),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2414),
.Y(n_3016)
);

OR2x2_ASAP7_75t_L g3017 ( 
.A(n_2701),
.B(n_2186),
.Y(n_3017)
);

BUFx3_ASAP7_75t_L g3018 ( 
.A(n_2447),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2431),
.Y(n_3019)
);

BUFx10_ASAP7_75t_L g3020 ( 
.A(n_2493),
.Y(n_3020)
);

NOR2xp33_ASAP7_75t_L g3021 ( 
.A(n_2413),
.B(n_2188),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_L g3022 ( 
.A(n_2593),
.B(n_2594),
.Y(n_3022)
);

AND2x6_ASAP7_75t_L g3023 ( 
.A(n_2646),
.B(n_2303),
.Y(n_3023)
);

INVx1_ASAP7_75t_SL g3024 ( 
.A(n_2726),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2336),
.Y(n_3025)
);

BUFx6f_ASAP7_75t_SL g3026 ( 
.A(n_2686),
.Y(n_3026)
);

INVx3_ASAP7_75t_L g3027 ( 
.A(n_2397),
.Y(n_3027)
);

INVx2_ASAP7_75t_L g3028 ( 
.A(n_2414),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2338),
.Y(n_3029)
);

INVx3_ASAP7_75t_L g3030 ( 
.A(n_2397),
.Y(n_3030)
);

AND2x4_ASAP7_75t_L g3031 ( 
.A(n_2564),
.B(n_2565),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2342),
.Y(n_3032)
);

BUFx2_ASAP7_75t_L g3033 ( 
.A(n_2670),
.Y(n_3033)
);

AND2x4_ASAP7_75t_L g3034 ( 
.A(n_2564),
.B(n_2206),
.Y(n_3034)
);

BUFx6f_ASAP7_75t_L g3035 ( 
.A(n_2400),
.Y(n_3035)
);

NOR2xp33_ASAP7_75t_L g3036 ( 
.A(n_2416),
.B(n_2194),
.Y(n_3036)
);

BUFx10_ASAP7_75t_L g3037 ( 
.A(n_2564),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_SL g3038 ( 
.A(n_2361),
.B(n_2220),
.Y(n_3038)
);

AND2x2_ASAP7_75t_L g3039 ( 
.A(n_2408),
.B(n_2215),
.Y(n_3039)
);

INVx2_ASAP7_75t_SL g3040 ( 
.A(n_2408),
.Y(n_3040)
);

BUFx2_ASAP7_75t_L g3041 ( 
.A(n_2354),
.Y(n_3041)
);

AND2x2_ASAP7_75t_L g3042 ( 
.A(n_2468),
.B(n_2251),
.Y(n_3042)
);

CKINVDCx5p33_ASAP7_75t_R g3043 ( 
.A(n_2422),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2345),
.Y(n_3044)
);

INVxp33_ASAP7_75t_SL g3045 ( 
.A(n_2463),
.Y(n_3045)
);

AND2x4_ASAP7_75t_L g3046 ( 
.A(n_2565),
.B(n_2220),
.Y(n_3046)
);

CKINVDCx20_ASAP7_75t_R g3047 ( 
.A(n_2361),
.Y(n_3047)
);

BUFx3_ASAP7_75t_L g3048 ( 
.A(n_2326),
.Y(n_3048)
);

BUFx2_ASAP7_75t_L g3049 ( 
.A(n_2686),
.Y(n_3049)
);

NOR2xp33_ASAP7_75t_L g3050 ( 
.A(n_2416),
.B(n_2194),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2599),
.B(n_2005),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2347),
.Y(n_3052)
);

NAND3x1_ASAP7_75t_L g3053 ( 
.A(n_2598),
.B(n_2318),
.C(n_2315),
.Y(n_3053)
);

BUFx6f_ASAP7_75t_L g3054 ( 
.A(n_2400),
.Y(n_3054)
);

OAI22xp5_ASAP7_75t_L g3055 ( 
.A1(n_2322),
.A2(n_2255),
.B1(n_2251),
.B2(n_2281),
.Y(n_3055)
);

BUFx6f_ASAP7_75t_L g3056 ( 
.A(n_2400),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2349),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_SL g3058 ( 
.A(n_2453),
.B(n_2221),
.Y(n_3058)
);

CKINVDCx5p33_ASAP7_75t_R g3059 ( 
.A(n_2453),
.Y(n_3059)
);

BUFx3_ASAP7_75t_L g3060 ( 
.A(n_2326),
.Y(n_3060)
);

AND2x2_ASAP7_75t_SL g3061 ( 
.A(n_2551),
.B(n_2310),
.Y(n_3061)
);

INVx4_ASAP7_75t_L g3062 ( 
.A(n_2686),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2351),
.Y(n_3063)
);

INVx3_ASAP7_75t_L g3064 ( 
.A(n_2400),
.Y(n_3064)
);

NOR2xp33_ASAP7_75t_L g3065 ( 
.A(n_2430),
.B(n_2200),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2355),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2360),
.Y(n_3067)
);

CKINVDCx5p33_ASAP7_75t_R g3068 ( 
.A(n_2477),
.Y(n_3068)
);

INVx5_ASAP7_75t_L g3069 ( 
.A(n_2444),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2362),
.Y(n_3070)
);

CKINVDCx20_ASAP7_75t_R g3071 ( 
.A(n_2477),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2603),
.B(n_2604),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_2417),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2363),
.Y(n_3074)
);

INVx4_ASAP7_75t_SL g3075 ( 
.A(n_2686),
.Y(n_3075)
);

INVx5_ASAP7_75t_L g3076 ( 
.A(n_2444),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_2417),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2370),
.Y(n_3078)
);

NAND2xp33_ASAP7_75t_L g3079 ( 
.A(n_2611),
.B(n_2303),
.Y(n_3079)
);

AOI22xp5_ASAP7_75t_L g3080 ( 
.A1(n_2686),
.A2(n_2255),
.B1(n_2283),
.B2(n_2276),
.Y(n_3080)
);

OR2x2_ASAP7_75t_L g3081 ( 
.A(n_2468),
.B(n_2319),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2374),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2379),
.Y(n_3083)
);

AND2x6_ASAP7_75t_L g3084 ( 
.A(n_2649),
.B(n_2304),
.Y(n_3084)
);

BUFx3_ASAP7_75t_L g3085 ( 
.A(n_2565),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2383),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_SL g3087 ( 
.A(n_2512),
.B(n_2221),
.Y(n_3087)
);

NOR2x1p5_ASAP7_75t_L g3088 ( 
.A(n_2654),
.B(n_2269),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2389),
.Y(n_3089)
);

OAI22xp33_ASAP7_75t_L g3090 ( 
.A1(n_2626),
.A2(n_2201),
.B1(n_2200),
.B2(n_2232),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_SL g3091 ( 
.A(n_2512),
.B(n_2232),
.Y(n_3091)
);

INVx4_ASAP7_75t_SL g3092 ( 
.A(n_2444),
.Y(n_3092)
);

BUFx4f_ASAP7_75t_L g3093 ( 
.A(n_2372),
.Y(n_3093)
);

BUFx6f_ASAP7_75t_L g3094 ( 
.A(n_2444),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2680),
.Y(n_3095)
);

AO21x2_ASAP7_75t_L g3096 ( 
.A1(n_2623),
.A2(n_2081),
.B(n_2169),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2681),
.Y(n_3097)
);

NAND2xp33_ASAP7_75t_L g3098 ( 
.A(n_2612),
.B(n_2304),
.Y(n_3098)
);

NOR3xp33_ASAP7_75t_L g3099 ( 
.A(n_2540),
.B(n_2193),
.C(n_2099),
.Y(n_3099)
);

INVx6_ASAP7_75t_L g3100 ( 
.A(n_2636),
.Y(n_3100)
);

INVx1_ASAP7_75t_SL g3101 ( 
.A(n_2734),
.Y(n_3101)
);

INVx2_ASAP7_75t_L g3102 ( 
.A(n_2420),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2586),
.Y(n_3103)
);

CKINVDCx20_ASAP7_75t_R g3104 ( 
.A(n_2540),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_L g3105 ( 
.A(n_2615),
.B(n_2619),
.Y(n_3105)
);

BUFx6f_ASAP7_75t_L g3106 ( 
.A(n_2495),
.Y(n_3106)
);

NAND3xp33_ASAP7_75t_L g3107 ( 
.A(n_2385),
.B(n_2185),
.C(n_2291),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2587),
.Y(n_3108)
);

OR2x2_ASAP7_75t_L g3109 ( 
.A(n_2484),
.B(n_2319),
.Y(n_3109)
);

NAND3x1_ASAP7_75t_L g3110 ( 
.A(n_2460),
.B(n_2319),
.C(n_2157),
.Y(n_3110)
);

INVx4_ASAP7_75t_L g3111 ( 
.A(n_2495),
.Y(n_3111)
);

NOR2xp33_ASAP7_75t_L g3112 ( 
.A(n_2430),
.B(n_2201),
.Y(n_3112)
);

INVx3_ASAP7_75t_L g3113 ( 
.A(n_2495),
.Y(n_3113)
);

BUFx6f_ASAP7_75t_L g3114 ( 
.A(n_2495),
.Y(n_3114)
);

INVx1_ASAP7_75t_SL g3115 ( 
.A(n_2734),
.Y(n_3115)
);

AND2x2_ASAP7_75t_L g3116 ( 
.A(n_2484),
.B(n_2168),
.Y(n_3116)
);

INVx3_ASAP7_75t_L g3117 ( 
.A(n_2516),
.Y(n_3117)
);

INVx2_ASAP7_75t_L g3118 ( 
.A(n_2420),
.Y(n_3118)
);

BUFx2_ASAP7_75t_L g3119 ( 
.A(n_2636),
.Y(n_3119)
);

INVxp67_ASAP7_75t_SL g3120 ( 
.A(n_2724),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2627),
.Y(n_3121)
);

BUFx4f_ASAP7_75t_L g3122 ( 
.A(n_2372),
.Y(n_3122)
);

INVx2_ASAP7_75t_L g3123 ( 
.A(n_2423),
.Y(n_3123)
);

BUFx6f_ASAP7_75t_L g3124 ( 
.A(n_2516),
.Y(n_3124)
);

OAI22xp5_ASAP7_75t_L g3125 ( 
.A1(n_2634),
.A2(n_2234),
.B1(n_2247),
.B2(n_2241),
.Y(n_3125)
);

INVx1_ASAP7_75t_SL g3126 ( 
.A(n_2534),
.Y(n_3126)
);

AND2x4_ASAP7_75t_L g3127 ( 
.A(n_2636),
.B(n_2234),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_SL g3128 ( 
.A(n_2590),
.B(n_2241),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2620),
.B(n_2005),
.Y(n_3129)
);

NOR2xp33_ASAP7_75t_L g3130 ( 
.A(n_2436),
.B(n_2247),
.Y(n_3130)
);

OR2x6_ASAP7_75t_L g3131 ( 
.A(n_2439),
.B(n_2176),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2635),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2637),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2640),
.Y(n_3134)
);

NOR2xp33_ASAP7_75t_L g3135 ( 
.A(n_2436),
.B(n_2254),
.Y(n_3135)
);

OAI22xp5_ASAP7_75t_L g3136 ( 
.A1(n_2518),
.A2(n_2254),
.B1(n_2264),
.B2(n_2258),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2423),
.Y(n_3137)
);

BUFx6f_ASAP7_75t_L g3138 ( 
.A(n_2516),
.Y(n_3138)
);

INVx2_ASAP7_75t_L g3139 ( 
.A(n_2424),
.Y(n_3139)
);

NOR2xp33_ASAP7_75t_L g3140 ( 
.A(n_2452),
.B(n_2258),
.Y(n_3140)
);

AND2x2_ASAP7_75t_L g3141 ( 
.A(n_2872),
.B(n_2906),
.Y(n_3141)
);

NOR2xp33_ASAP7_75t_L g3142 ( 
.A(n_2736),
.B(n_2302),
.Y(n_3142)
);

BUFx3_ASAP7_75t_L g3143 ( 
.A(n_2843),
.Y(n_3143)
);

NOR2xp33_ASAP7_75t_L g3144 ( 
.A(n_2736),
.B(n_2302),
.Y(n_3144)
);

NOR2xp33_ASAP7_75t_L g3145 ( 
.A(n_2814),
.B(n_2304),
.Y(n_3145)
);

AOI22x1_ASAP7_75t_L g3146 ( 
.A1(n_3043),
.A2(n_2163),
.B1(n_2166),
.B2(n_2264),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_L g3147 ( 
.A(n_3101),
.B(n_2534),
.Y(n_3147)
);

INVx2_ASAP7_75t_L g3148 ( 
.A(n_2738),
.Y(n_3148)
);

NOR2xp33_ASAP7_75t_SL g3149 ( 
.A(n_3045),
.B(n_1953),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_L g3150 ( 
.A(n_3101),
.B(n_2266),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_2944),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_3115),
.B(n_2266),
.Y(n_3152)
);

INVx2_ASAP7_75t_L g3153 ( 
.A(n_2739),
.Y(n_3153)
);

AND2x2_ASAP7_75t_L g3154 ( 
.A(n_2924),
.B(n_2939),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_L g3155 ( 
.A(n_3115),
.B(n_2272),
.Y(n_3155)
);

NAND2xp5_ASAP7_75t_L g3156 ( 
.A(n_2814),
.B(n_2272),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_2817),
.B(n_1930),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_L g3158 ( 
.A(n_2817),
.B(n_2168),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_3126),
.B(n_2172),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_3126),
.B(n_2172),
.Y(n_3160)
);

INVx2_ASAP7_75t_L g3161 ( 
.A(n_2749),
.Y(n_3161)
);

AOI22xp33_ASAP7_75t_L g3162 ( 
.A1(n_2791),
.A2(n_2182),
.B1(n_2384),
.B2(n_2371),
.Y(n_3162)
);

NOR2xp67_ASAP7_75t_L g3163 ( 
.A(n_2748),
.B(n_2083),
.Y(n_3163)
);

INVx2_ASAP7_75t_SL g3164 ( 
.A(n_2740),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_SL g3165 ( 
.A(n_2850),
.B(n_2304),
.Y(n_3165)
);

OAI22xp33_ASAP7_75t_L g3166 ( 
.A1(n_2775),
.A2(n_2790),
.B1(n_2792),
.B2(n_2791),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_3095),
.Y(n_3167)
);

O2A1O1Ixp5_ASAP7_75t_L g3168 ( 
.A1(n_2824),
.A2(n_2683),
.B(n_2697),
.C(n_2669),
.Y(n_3168)
);

OAI22xp5_ASAP7_75t_L g3169 ( 
.A1(n_2805),
.A2(n_2561),
.B1(n_2628),
.B2(n_2585),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_3097),
.Y(n_3170)
);

AOI22xp5_ASAP7_75t_L g3171 ( 
.A1(n_2975),
.A2(n_2099),
.B1(n_2083),
.B2(n_2305),
.Y(n_3171)
);

INVx4_ASAP7_75t_L g3172 ( 
.A(n_2748),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_SL g3173 ( 
.A(n_2891),
.B(n_2218),
.Y(n_3173)
);

NAND3xp33_ASAP7_75t_L g3174 ( 
.A(n_2805),
.B(n_2257),
.C(n_2235),
.Y(n_3174)
);

NOR2xp33_ASAP7_75t_L g3175 ( 
.A(n_2997),
.B(n_2178),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2758),
.Y(n_3176)
);

AND2x2_ASAP7_75t_L g3177 ( 
.A(n_3039),
.B(n_2178),
.Y(n_3177)
);

NOR2xp33_ASAP7_75t_L g3178 ( 
.A(n_3042),
.B(n_2180),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_3116),
.B(n_2180),
.Y(n_3179)
);

OAI221xp5_ASAP7_75t_L g3180 ( 
.A1(n_2934),
.A2(n_2044),
.B1(n_2305),
.B2(n_2270),
.C(n_2288),
.Y(n_3180)
);

INVx2_ASAP7_75t_L g3181 ( 
.A(n_2761),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_SL g3182 ( 
.A(n_2824),
.B(n_2222),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_L g3183 ( 
.A(n_2772),
.B(n_2792),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_SL g3184 ( 
.A(n_2908),
.B(n_2239),
.Y(n_3184)
);

AO22x1_ASAP7_75t_L g3185 ( 
.A1(n_2889),
.A2(n_2300),
.B1(n_1980),
.B2(n_2011),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_2775),
.B(n_2703),
.Y(n_3186)
);

BUFx3_ASAP7_75t_L g3187 ( 
.A(n_2747),
.Y(n_3187)
);

AOI22xp33_ASAP7_75t_L g3188 ( 
.A1(n_2868),
.A2(n_2393),
.B1(n_2313),
.B2(n_2452),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_2790),
.B(n_2451),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_2759),
.Y(n_3190)
);

NOR2xp33_ASAP7_75t_L g3191 ( 
.A(n_2908),
.B(n_2292),
.Y(n_3191)
);

AND2x2_ASAP7_75t_L g3192 ( 
.A(n_2776),
.B(n_1996),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_SL g3193 ( 
.A(n_3011),
.B(n_2240),
.Y(n_3193)
);

AOI22xp33_ASAP7_75t_L g3194 ( 
.A1(n_2868),
.A2(n_2456),
.B1(n_2480),
.B2(n_2466),
.Y(n_3194)
);

HB1xp67_ASAP7_75t_SL g3195 ( 
.A(n_2894),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2766),
.Y(n_3196)
);

AOI22xp5_ASAP7_75t_L g3197 ( 
.A1(n_3047),
.A2(n_3104),
.B1(n_3071),
.B2(n_2752),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_2773),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_L g3199 ( 
.A(n_2799),
.B(n_3040),
.Y(n_3199)
);

INVx2_ASAP7_75t_L g3200 ( 
.A(n_2769),
.Y(n_3200)
);

OR2x2_ASAP7_75t_L g3201 ( 
.A(n_2813),
.B(n_2310),
.Y(n_3201)
);

NAND3xp33_ASAP7_75t_L g3202 ( 
.A(n_3107),
.B(n_2964),
.C(n_2895),
.Y(n_3202)
);

CKINVDCx5p33_ASAP7_75t_R g3203 ( 
.A(n_2897),
.Y(n_3203)
);

INVxp67_ASAP7_75t_L g3204 ( 
.A(n_3007),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_SL g3205 ( 
.A(n_2827),
.B(n_2649),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_SL g3206 ( 
.A(n_2827),
.B(n_2652),
.Y(n_3206)
);

INVx2_ASAP7_75t_SL g3207 ( 
.A(n_2740),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_SL g3208 ( 
.A(n_2984),
.B(n_2652),
.Y(n_3208)
);

AOI22xp33_ASAP7_75t_L g3209 ( 
.A1(n_2964),
.A2(n_2456),
.B1(n_2480),
.B2(n_2466),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_L g3210 ( 
.A(n_2799),
.B(n_2005),
.Y(n_3210)
);

INVx3_ASAP7_75t_L g3211 ( 
.A(n_2884),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_2779),
.Y(n_3212)
);

INVxp67_ASAP7_75t_L g3213 ( 
.A(n_3007),
.Y(n_3213)
);

INVx2_ASAP7_75t_L g3214 ( 
.A(n_2771),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_SL g3215 ( 
.A(n_3011),
.B(n_2249),
.Y(n_3215)
);

BUFx3_ASAP7_75t_L g3216 ( 
.A(n_2780),
.Y(n_3216)
);

INVx2_ASAP7_75t_L g3217 ( 
.A(n_2801),
.Y(n_3217)
);

AOI22xp5_ASAP7_75t_L g3218 ( 
.A1(n_2750),
.A2(n_2294),
.B1(n_2299),
.B2(n_2176),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2782),
.Y(n_3219)
);

NOR2xp33_ASAP7_75t_L g3220 ( 
.A(n_2895),
.B(n_2295),
.Y(n_3220)
);

AND2x6_ASAP7_75t_L g3221 ( 
.A(n_3075),
.B(n_2656),
.Y(n_3221)
);

OAI22xp5_ASAP7_75t_L g3222 ( 
.A1(n_3107),
.A2(n_2597),
.B1(n_2560),
.B2(n_2261),
.Y(n_3222)
);

NOR2xp33_ASAP7_75t_L g3223 ( 
.A(n_2750),
.B(n_2256),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_2787),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_2751),
.B(n_1996),
.Y(n_3225)
);

INVx2_ASAP7_75t_L g3226 ( 
.A(n_2823),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_2751),
.B(n_2461),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_L g3228 ( 
.A(n_2767),
.B(n_2271),
.Y(n_3228)
);

AOI22xp33_ASAP7_75t_L g3229 ( 
.A1(n_2741),
.A2(n_2492),
.B1(n_2498),
.B2(n_2337),
.Y(n_3229)
);

INVx2_ASAP7_75t_L g3230 ( 
.A(n_2826),
.Y(n_3230)
);

INVx2_ASAP7_75t_SL g3231 ( 
.A(n_2744),
.Y(n_3231)
);

BUFx6f_ASAP7_75t_L g3232 ( 
.A(n_2845),
.Y(n_3232)
);

AND2x2_ASAP7_75t_L g3233 ( 
.A(n_2847),
.B(n_2017),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_SL g3234 ( 
.A(n_3059),
.B(n_2267),
.Y(n_3234)
);

AND2x2_ASAP7_75t_L g3235 ( 
.A(n_3048),
.B(n_2017),
.Y(n_3235)
);

NOR2xp33_ASAP7_75t_L g3236 ( 
.A(n_2752),
.B(n_2279),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_2795),
.Y(n_3237)
);

NOR2xp33_ASAP7_75t_L g3238 ( 
.A(n_2762),
.B(n_2175),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_L g3239 ( 
.A(n_2767),
.B(n_2039),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_L g3240 ( 
.A(n_2753),
.B(n_2039),
.Y(n_3240)
);

INVx2_ASAP7_75t_SL g3241 ( 
.A(n_2744),
.Y(n_3241)
);

NOR2xp33_ASAP7_75t_L g3242 ( 
.A(n_2762),
.B(n_2184),
.Y(n_3242)
);

O2A1O1Ixp33_ASAP7_75t_L g3243 ( 
.A1(n_2905),
.A2(n_2569),
.B(n_2104),
.C(n_2669),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_2753),
.B(n_1973),
.Y(n_3244)
);

AND2x6_ASAP7_75t_SL g3245 ( 
.A(n_2764),
.B(n_1994),
.Y(n_3245)
);

INVx2_ASAP7_75t_L g3246 ( 
.A(n_2854),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_2786),
.B(n_1973),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_SL g3248 ( 
.A(n_2984),
.B(n_2656),
.Y(n_3248)
);

BUFx3_ASAP7_75t_L g3249 ( 
.A(n_2784),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_SL g3250 ( 
.A(n_3068),
.B(n_2075),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_2786),
.B(n_1973),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_3060),
.B(n_2087),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_2905),
.B(n_2094),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_3012),
.B(n_2110),
.Y(n_3254)
);

INVx2_ASAP7_75t_L g3255 ( 
.A(n_2857),
.Y(n_3255)
);

OR2x2_ASAP7_75t_L g3256 ( 
.A(n_2965),
.B(n_2310),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_L g3257 ( 
.A(n_3012),
.B(n_2340),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_3014),
.B(n_2104),
.Y(n_3258)
);

NOR2xp33_ASAP7_75t_L g3259 ( 
.A(n_2774),
.B(n_2187),
.Y(n_3259)
);

NOR2xp33_ASAP7_75t_L g3260 ( 
.A(n_2774),
.B(n_2189),
.Y(n_3260)
);

AND2x2_ASAP7_75t_L g3261 ( 
.A(n_2871),
.B(n_2190),
.Y(n_3261)
);

AND2x6_ASAP7_75t_SL g3262 ( 
.A(n_2764),
.B(n_1994),
.Y(n_3262)
);

INVx2_ASAP7_75t_SL g3263 ( 
.A(n_2887),
.Y(n_3263)
);

NOR3xp33_ASAP7_75t_L g3264 ( 
.A(n_3055),
.B(n_2044),
.C(n_2618),
.Y(n_3264)
);

INVx2_ASAP7_75t_SL g3265 ( 
.A(n_2853),
.Y(n_3265)
);

INVx2_ASAP7_75t_SL g3266 ( 
.A(n_2853),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_3014),
.B(n_2591),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_2800),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_SL g3269 ( 
.A(n_3080),
.B(n_2134),
.Y(n_3269)
);

NAND2xp33_ASAP7_75t_SL g3270 ( 
.A(n_2831),
.B(n_1980),
.Y(n_3270)
);

NOR2xp33_ASAP7_75t_L g3271 ( 
.A(n_3017),
.B(n_2192),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_2803),
.Y(n_3272)
);

AOI22xp33_ASAP7_75t_L g3273 ( 
.A1(n_2741),
.A2(n_2492),
.B1(n_2498),
.B2(n_2310),
.Y(n_3273)
);

NOR2xp33_ASAP7_75t_SL g3274 ( 
.A(n_2912),
.B(n_2079),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_2804),
.Y(n_3275)
);

OAI22xp33_ASAP7_75t_L g3276 ( 
.A1(n_3081),
.A2(n_2668),
.B1(n_2674),
.B2(n_2666),
.Y(n_3276)
);

AOI22xp5_ASAP7_75t_L g3277 ( 
.A1(n_2783),
.A2(n_1985),
.B1(n_2028),
.B2(n_2011),
.Y(n_3277)
);

NOR2xp33_ASAP7_75t_L g3278 ( 
.A(n_2770),
.B(n_2196),
.Y(n_3278)
);

OR2x2_ASAP7_75t_L g3279 ( 
.A(n_3004),
.B(n_2144),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_L g3280 ( 
.A(n_2830),
.B(n_2837),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_2830),
.B(n_2676),
.Y(n_3281)
);

INVx2_ASAP7_75t_SL g3282 ( 
.A(n_2968),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_L g3283 ( 
.A(n_2837),
.B(n_2677),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_3090),
.B(n_2679),
.Y(n_3284)
);

NOR2xp33_ASAP7_75t_L g3285 ( 
.A(n_2770),
.B(n_2202),
.Y(n_3285)
);

NOR2xp33_ASAP7_75t_L g3286 ( 
.A(n_2898),
.B(n_2783),
.Y(n_3286)
);

INVxp67_ASAP7_75t_SL g3287 ( 
.A(n_2932),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_3090),
.B(n_1956),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_2806),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_2802),
.B(n_1956),
.Y(n_3290)
);

INVx4_ASAP7_75t_L g3291 ( 
.A(n_2755),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_L g3292 ( 
.A(n_2802),
.B(n_1956),
.Y(n_3292)
);

INVx2_ASAP7_75t_L g3293 ( 
.A(n_2862),
.Y(n_3293)
);

AOI22xp5_ASAP7_75t_L g3294 ( 
.A1(n_2835),
.A2(n_2028),
.B1(n_2038),
.B2(n_1985),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_2811),
.B(n_2508),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_2810),
.Y(n_3296)
);

INVx2_ASAP7_75t_L g3297 ( 
.A(n_2863),
.Y(n_3297)
);

NOR2xp33_ASAP7_75t_L g3298 ( 
.A(n_2898),
.B(n_2208),
.Y(n_3298)
);

AND2x6_ASAP7_75t_SL g3299 ( 
.A(n_2764),
.B(n_2032),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_SL g3300 ( 
.A(n_3062),
.B(n_2664),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_L g3301 ( 
.A(n_2811),
.B(n_2914),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_SL g3302 ( 
.A(n_2929),
.B(n_2020),
.Y(n_3302)
);

OAI22x1_ASAP7_75t_SL g3303 ( 
.A1(n_2880),
.A2(n_2139),
.B1(n_2224),
.B2(n_2100),
.Y(n_3303)
);

NAND3xp33_ASAP7_75t_L g3304 ( 
.A(n_3099),
.B(n_2065),
.C(n_2038),
.Y(n_3304)
);

INVx2_ASAP7_75t_L g3305 ( 
.A(n_2867),
.Y(n_3305)
);

NOR2xp33_ASAP7_75t_L g3306 ( 
.A(n_2995),
.B(n_2211),
.Y(n_3306)
);

NAND3xp33_ASAP7_75t_L g3307 ( 
.A(n_3099),
.B(n_2065),
.C(n_2300),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_2914),
.B(n_3034),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_2815),
.Y(n_3309)
);

INVx4_ASAP7_75t_L g3310 ( 
.A(n_2755),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_3034),
.B(n_2046),
.Y(n_3311)
);

NOR2xp33_ASAP7_75t_L g3312 ( 
.A(n_3018),
.B(n_2502),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_2818),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_2819),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_2881),
.Y(n_3315)
);

OR2x2_ASAP7_75t_L g3316 ( 
.A(n_2973),
.B(n_2829),
.Y(n_3316)
);

BUFx8_ASAP7_75t_L g3317 ( 
.A(n_2851),
.Y(n_3317)
);

OAI22xp5_ASAP7_75t_L g3318 ( 
.A1(n_2825),
.A2(n_2343),
.B1(n_2523),
.B2(n_2500),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_2902),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_L g3320 ( 
.A(n_3046),
.B(n_2616),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_3046),
.B(n_2589),
.Y(n_3321)
);

OAI22xp5_ASAP7_75t_L g3322 ( 
.A1(n_2825),
.A2(n_2343),
.B1(n_2523),
.B2(n_2500),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_SL g3323 ( 
.A(n_3062),
.B(n_2664),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_SL g3324 ( 
.A(n_2929),
.B(n_2020),
.Y(n_3324)
);

AOI21x1_ASAP7_75t_L g3325 ( 
.A1(n_2915),
.A2(n_2624),
.B(n_2623),
.Y(n_3325)
);

OAI22xp33_ASAP7_75t_L g3326 ( 
.A1(n_3109),
.A2(n_2497),
.B1(n_2525),
.B2(n_2520),
.Y(n_3326)
);

AO221x1_ASAP7_75t_L g3327 ( 
.A1(n_2974),
.A2(n_1988),
.B1(n_2472),
.B2(n_2550),
.C(n_2259),
.Y(n_3327)
);

INVx4_ASAP7_75t_L g3328 ( 
.A(n_2785),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_2821),
.Y(n_3329)
);

AND2x2_ASAP7_75t_L g3330 ( 
.A(n_3024),
.B(n_2269),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_3127),
.B(n_2589),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_3127),
.B(n_2608),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_SL g3333 ( 
.A(n_2937),
.B(n_2307),
.Y(n_3333)
);

AND2x2_ASAP7_75t_L g3334 ( 
.A(n_3024),
.B(n_2490),
.Y(n_3334)
);

NAND2xp33_ASAP7_75t_L g3335 ( 
.A(n_2951),
.B(n_2090),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_3008),
.B(n_2608),
.Y(n_3336)
);

AND2x4_ASAP7_75t_SL g3337 ( 
.A(n_2785),
.B(n_2100),
.Y(n_3337)
);

NOR2xp33_ASAP7_75t_L g3338 ( 
.A(n_3031),
.B(n_2502),
.Y(n_3338)
);

AND2x2_ASAP7_75t_L g3339 ( 
.A(n_3031),
.B(n_2307),
.Y(n_3339)
);

BUFx12f_ASAP7_75t_L g3340 ( 
.A(n_2846),
.Y(n_3340)
);

NAND2x1p5_ASAP7_75t_L g3341 ( 
.A(n_2861),
.B(n_2359),
.Y(n_3341)
);

NOR2xp33_ASAP7_75t_L g3342 ( 
.A(n_3119),
.B(n_2546),
.Y(n_3342)
);

NAND2xp33_ASAP7_75t_L g3343 ( 
.A(n_2951),
.B(n_2998),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_3008),
.B(n_2638),
.Y(n_3344)
);

NOR2xp33_ASAP7_75t_L g3345 ( 
.A(n_3130),
.B(n_2546),
.Y(n_3345)
);

INVx2_ASAP7_75t_L g3346 ( 
.A(n_2907),
.Y(n_3346)
);

INVx2_ASAP7_75t_L g3347 ( 
.A(n_2911),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_SL g3348 ( 
.A(n_2861),
.B(n_2665),
.Y(n_3348)
);

AOI22xp33_ASAP7_75t_SL g3349 ( 
.A1(n_2974),
.A2(n_2224),
.B1(n_2253),
.B2(n_2139),
.Y(n_3349)
);

INVx2_ASAP7_75t_SL g3350 ( 
.A(n_2745),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_2937),
.B(n_2638),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_2943),
.B(n_2662),
.Y(n_3352)
);

NAND3xp33_ASAP7_75t_L g3353 ( 
.A(n_3130),
.B(n_3140),
.C(n_3135),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_SL g3354 ( 
.A(n_2943),
.B(n_2618),
.Y(n_3354)
);

AND2x4_ASAP7_75t_L g3355 ( 
.A(n_2760),
.B(n_2683),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_3010),
.B(n_2662),
.Y(n_3356)
);

CKINVDCx5p33_ASAP7_75t_R g3357 ( 
.A(n_2841),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_L g3358 ( 
.A(n_3010),
.B(n_3021),
.Y(n_3358)
);

AOI21xp5_ASAP7_75t_L g3359 ( 
.A1(n_2932),
.A2(n_2625),
.B(n_2624),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_SL g3360 ( 
.A(n_3055),
.B(n_2633),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_3021),
.B(n_2667),
.Y(n_3361)
);

XNOR2xp5_ASAP7_75t_L g3362 ( 
.A(n_2778),
.B(n_1839),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_2834),
.Y(n_3363)
);

AOI22xp33_ASAP7_75t_SL g3364 ( 
.A1(n_2974),
.A2(n_2275),
.B1(n_2317),
.B2(n_2253),
.Y(n_3364)
);

AND2x2_ASAP7_75t_L g3365 ( 
.A(n_2969),
.B(n_2260),
.Y(n_3365)
);

BUFx5_ASAP7_75t_L g3366 ( 
.A(n_2788),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_L g3367 ( 
.A(n_3036),
.B(n_3050),
.Y(n_3367)
);

OAI22xp5_ASAP7_75t_L g3368 ( 
.A1(n_2832),
.A2(n_2524),
.B1(n_2531),
.B2(n_2523),
.Y(n_3368)
);

NOR2xp33_ASAP7_75t_L g3369 ( 
.A(n_3135),
.B(n_2573),
.Y(n_3369)
);

AND2x2_ASAP7_75t_L g3370 ( 
.A(n_2945),
.B(n_2114),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_2855),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_L g3372 ( 
.A(n_3036),
.B(n_2667),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_3050),
.B(n_2573),
.Y(n_3373)
);

INVx2_ASAP7_75t_SL g3374 ( 
.A(n_2809),
.Y(n_3374)
);

AND2x6_ASAP7_75t_L g3375 ( 
.A(n_3075),
.B(n_2665),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_SL g3376 ( 
.A(n_2922),
.B(n_2717),
.Y(n_3376)
);

BUFx6f_ASAP7_75t_L g3377 ( 
.A(n_2845),
.Y(n_3377)
);

AOI221xp5_ASAP7_75t_L g3378 ( 
.A1(n_3125),
.A2(n_2696),
.B1(n_2717),
.B2(n_2633),
.C(n_2308),
.Y(n_3378)
);

INVx1_ASAP7_75t_L g3379 ( 
.A(n_2856),
.Y(n_3379)
);

NOR2xp33_ASAP7_75t_L g3380 ( 
.A(n_3140),
.B(n_3001),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_2860),
.Y(n_3381)
);

INVx2_ASAP7_75t_SL g3382 ( 
.A(n_2789),
.Y(n_3382)
);

INVx2_ASAP7_75t_L g3383 ( 
.A(n_2927),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_3065),
.B(n_2697),
.Y(n_3384)
);

INVx2_ASAP7_75t_L g3385 ( 
.A(n_2933),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_SL g3386 ( 
.A(n_2832),
.B(n_2729),
.Y(n_3386)
);

AOI21xp5_ASAP7_75t_L g3387 ( 
.A1(n_2990),
.A2(n_2639),
.B(n_2625),
.Y(n_3387)
);

OAI221xp5_ASAP7_75t_L g3388 ( 
.A1(n_3125),
.A2(n_2273),
.B1(n_2167),
.B2(n_2115),
.C(n_2696),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_3065),
.B(n_3112),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_3112),
.B(n_2177),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_2972),
.B(n_2536),
.Y(n_3391)
);

AOI22xp33_ASAP7_75t_L g3392 ( 
.A1(n_2765),
.A2(n_2073),
.B1(n_2103),
.B2(n_2072),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_2865),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_2972),
.B(n_2537),
.Y(n_3394)
);

O2A1O1Ixp33_ASAP7_75t_L g3395 ( 
.A1(n_3136),
.A2(n_2081),
.B(n_2162),
.C(n_2702),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_2760),
.B(n_2544),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_2763),
.B(n_2439),
.Y(n_3397)
);

O2A1O1Ixp5_ASAP7_75t_L g3398 ( 
.A1(n_3038),
.A2(n_2296),
.B(n_2639),
.C(n_2368),
.Y(n_3398)
);

BUFx3_ASAP7_75t_L g3399 ( 
.A(n_3041),
.Y(n_3399)
);

NOR2xp33_ASAP7_75t_SL g3400 ( 
.A(n_2873),
.B(n_2079),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_2763),
.B(n_2729),
.Y(n_3401)
);

INVx2_ASAP7_75t_SL g3402 ( 
.A(n_2789),
.Y(n_3402)
);

INVx2_ASAP7_75t_L g3403 ( 
.A(n_2947),
.Y(n_3403)
);

OR2x2_ASAP7_75t_L g3404 ( 
.A(n_2820),
.B(n_2308),
.Y(n_3404)
);

INVx2_ASAP7_75t_L g3405 ( 
.A(n_2950),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_SL g3406 ( 
.A(n_2831),
.B(n_2273),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_2869),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_SL g3408 ( 
.A(n_2839),
.B(n_2027),
.Y(n_3408)
);

OAI221xp5_ASAP7_75t_L g3409 ( 
.A1(n_2765),
.A2(n_2007),
.B1(n_1005),
.B2(n_1020),
.C(n_1003),
.Y(n_3409)
);

AND2x2_ASAP7_75t_L g3410 ( 
.A(n_3033),
.B(n_1967),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_SL g3411 ( 
.A(n_2839),
.B(n_2731),
.Y(n_3411)
);

NOR2xp33_ASAP7_75t_SL g3412 ( 
.A(n_2793),
.B(n_2275),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_2777),
.B(n_2731),
.Y(n_3413)
);

AND2x2_ASAP7_75t_L g3414 ( 
.A(n_2807),
.B(n_1840),
.Y(n_3414)
);

BUFx3_ASAP7_75t_L g3415 ( 
.A(n_2959),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_SL g3416 ( 
.A(n_2840),
.B(n_2359),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_2870),
.Y(n_3417)
);

INVx2_ASAP7_75t_L g3418 ( 
.A(n_2953),
.Y(n_3418)
);

AND2x2_ASAP7_75t_L g3419 ( 
.A(n_3061),
.B(n_1846),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_2777),
.B(n_2368),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_SL g3421 ( 
.A(n_2844),
.B(n_2941),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_SL g3422 ( 
.A(n_2941),
.B(n_2368),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_L g3423 ( 
.A(n_3051),
.B(n_2429),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_3051),
.B(n_2429),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_3129),
.B(n_2429),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_2874),
.Y(n_3426)
);

INVx2_ASAP7_75t_L g3427 ( 
.A(n_2966),
.Y(n_3427)
);

OAI21xp5_ASAP7_75t_L g3428 ( 
.A1(n_2848),
.A2(n_2437),
.B(n_2428),
.Y(n_3428)
);

AOI22xp33_ASAP7_75t_L g3429 ( 
.A1(n_3005),
.A2(n_2073),
.B1(n_2103),
.B2(n_2072),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_L g3430 ( 
.A(n_3129),
.B(n_2486),
.Y(n_3430)
);

NOR2xp33_ASAP7_75t_L g3431 ( 
.A(n_3001),
.B(n_3100),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_SL g3432 ( 
.A(n_2822),
.B(n_2486),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_2948),
.B(n_2486),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_2875),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_2948),
.B(n_2659),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_2878),
.Y(n_3436)
);

AND2x2_ASAP7_75t_SL g3437 ( 
.A(n_3049),
.B(n_3005),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_SL g3438 ( 
.A(n_2798),
.B(n_2516),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_2879),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_2962),
.B(n_2660),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_2882),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_2883),
.Y(n_3442)
);

CKINVDCx5p33_ASAP7_75t_R g3443 ( 
.A(n_2742),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_2888),
.Y(n_3444)
);

CKINVDCx20_ASAP7_75t_R g3445 ( 
.A(n_2742),
.Y(n_3445)
);

NOR3xp33_ASAP7_75t_L g3446 ( 
.A(n_3136),
.B(n_2032),
.C(n_1003),
.Y(n_3446)
);

AOI22xp33_ASAP7_75t_L g3447 ( 
.A1(n_3026),
.A2(n_3132),
.B1(n_3133),
.B2(n_3121),
.Y(n_3447)
);

AOI22xp33_ASAP7_75t_L g3448 ( 
.A1(n_3026),
.A2(n_2073),
.B1(n_2103),
.B2(n_2072),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_2962),
.B(n_2661),
.Y(n_3449)
);

A2O1A1Ixp33_ASAP7_75t_L g3450 ( 
.A1(n_2798),
.A2(n_2721),
.B(n_2723),
.C(n_2720),
.Y(n_3450)
);

NAND2xp33_ASAP7_75t_SL g3451 ( 
.A(n_2816),
.B(n_2524),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_SL g3452 ( 
.A(n_2822),
.B(n_2663),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_2978),
.B(n_2986),
.Y(n_3453)
);

INVxp67_ASAP7_75t_L g3454 ( 
.A(n_2812),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_2893),
.Y(n_3455)
);

NOR2xp33_ASAP7_75t_L g3456 ( 
.A(n_3001),
.B(n_2524),
.Y(n_3456)
);

AOI22xp5_ASAP7_75t_L g3457 ( 
.A1(n_2812),
.A2(n_2317),
.B1(n_1848),
.B2(n_1872),
.Y(n_3457)
);

BUFx3_ASAP7_75t_L g3458 ( 
.A(n_2866),
.Y(n_3458)
);

NOR2xp33_ASAP7_75t_L g3459 ( 
.A(n_3100),
.B(n_2531),
.Y(n_3459)
);

AOI21xp5_ASAP7_75t_L g3460 ( 
.A1(n_2990),
.A2(n_2539),
.B(n_2531),
.Y(n_3460)
);

OAI221xp5_ASAP7_75t_L g3461 ( 
.A1(n_2940),
.A2(n_1020),
.B1(n_1023),
.B2(n_1005),
.C(n_996),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_2978),
.B(n_2704),
.Y(n_3462)
);

INVx2_ASAP7_75t_L g3463 ( 
.A(n_2977),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_L g3464 ( 
.A(n_2986),
.B(n_2705),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_2983),
.Y(n_3465)
);

INVx2_ASAP7_75t_L g3466 ( 
.A(n_2994),
.Y(n_3466)
);

NOR2xp33_ASAP7_75t_L g3467 ( 
.A(n_3100),
.B(n_2539),
.Y(n_3467)
);

INVx3_ASAP7_75t_L g3468 ( 
.A(n_2884),
.Y(n_3468)
);

OAI22xp33_ASAP7_75t_L g3469 ( 
.A1(n_2842),
.A2(n_1063),
.B1(n_1076),
.B2(n_1030),
.Y(n_3469)
);

INVxp33_ASAP7_75t_L g3470 ( 
.A(n_2985),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_SL g3471 ( 
.A(n_2836),
.B(n_2710),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_2903),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_L g3473 ( 
.A(n_2909),
.B(n_2713),
.Y(n_3473)
);

AOI22xp33_ASAP7_75t_L g3474 ( 
.A1(n_3134),
.A2(n_2103),
.B1(n_2073),
.B2(n_2424),
.Y(n_3474)
);

NOR2xp33_ASAP7_75t_L g3475 ( 
.A(n_2816),
.B(n_2539),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_2918),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_2919),
.B(n_2716),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_2926),
.B(n_2730),
.Y(n_3478)
);

OAI22x1_ASAP7_75t_R g3479 ( 
.A1(n_2896),
.A2(n_1848),
.B1(n_1872),
.B2(n_1846),
.Y(n_3479)
);

BUFx5_ASAP7_75t_L g3480 ( 
.A(n_2788),
.Y(n_3480)
);

INVxp67_ASAP7_75t_L g3481 ( 
.A(n_2896),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_2935),
.B(n_2732),
.Y(n_3482)
);

OAI22xp5_ASAP7_75t_SL g3483 ( 
.A1(n_2930),
.A2(n_1890),
.B1(n_1886),
.B2(n_887),
.Y(n_3483)
);

INVx3_ASAP7_75t_L g3484 ( 
.A(n_2904),
.Y(n_3484)
);

AOI22xp5_ASAP7_75t_L g3485 ( 
.A1(n_2930),
.A2(n_2960),
.B1(n_2971),
.B2(n_2957),
.Y(n_3485)
);

BUFx3_ASAP7_75t_L g3486 ( 
.A(n_2793),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_2942),
.B(n_2733),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_2946),
.B(n_2571),
.Y(n_3488)
);

NOR2xp33_ASAP7_75t_L g3489 ( 
.A(n_3058),
.B(n_2571),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_2963),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_2967),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_L g3492 ( 
.A(n_2970),
.B(n_2571),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_2976),
.B(n_2428),
.Y(n_3493)
);

OAI22xp5_ASAP7_75t_L g3494 ( 
.A1(n_2848),
.A2(n_2631),
.B1(n_2632),
.B2(n_2601),
.Y(n_3494)
);

INVx3_ASAP7_75t_L g3495 ( 
.A(n_2904),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_L g3496 ( 
.A(n_2979),
.B(n_2437),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_2982),
.B(n_2438),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_2988),
.Y(n_3498)
);

OAI22xp33_ASAP7_75t_L g3499 ( 
.A1(n_2842),
.A2(n_2991),
.B1(n_3009),
.B2(n_2999),
.Y(n_3499)
);

INVxp67_ASAP7_75t_SL g3500 ( 
.A(n_3120),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_SL g3501 ( 
.A(n_2845),
.B(n_2542),
.Y(n_3501)
);

A2O1A1Ixp33_ASAP7_75t_L g3502 ( 
.A1(n_2949),
.A2(n_2438),
.B(n_2441),
.C(n_2440),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_3019),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3025),
.Y(n_3504)
);

INVx2_ASAP7_75t_SL g3505 ( 
.A(n_2796),
.Y(n_3505)
);

AOI221xp5_ASAP7_75t_L g3506 ( 
.A1(n_2768),
.A2(n_1508),
.B1(n_1511),
.B2(n_1507),
.C(n_1505),
.Y(n_3506)
);

NOR2xp33_ASAP7_75t_L g3507 ( 
.A(n_3087),
.B(n_3091),
.Y(n_3507)
);

NOR3x1_ASAP7_75t_L g3508 ( 
.A(n_2916),
.B(n_1028),
.C(n_1023),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_3029),
.Y(n_3509)
);

NOR2xp33_ASAP7_75t_L g3510 ( 
.A(n_3085),
.B(n_2949),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_2836),
.B(n_2440),
.Y(n_3511)
);

INVx2_ASAP7_75t_L g3512 ( 
.A(n_3002),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_L g3513 ( 
.A(n_2849),
.B(n_2441),
.Y(n_3513)
);

OR2x2_ASAP7_75t_L g3514 ( 
.A(n_3131),
.B(n_1886),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3032),
.Y(n_3515)
);

AOI22xp33_ASAP7_75t_L g3516 ( 
.A1(n_3044),
.A2(n_2427),
.B1(n_2504),
.B2(n_2503),
.Y(n_3516)
);

INVx2_ASAP7_75t_L g3517 ( 
.A(n_3016),
.Y(n_3517)
);

INVx2_ASAP7_75t_L g3518 ( 
.A(n_3148),
.Y(n_3518)
);

BUFx3_ASAP7_75t_L g3519 ( 
.A(n_3187),
.Y(n_3519)
);

OR2x2_ASAP7_75t_L g3520 ( 
.A(n_3201),
.B(n_3131),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3142),
.B(n_2849),
.Y(n_3521)
);

OAI22xp5_ASAP7_75t_L g3522 ( 
.A1(n_3191),
.A2(n_2980),
.B1(n_2952),
.B2(n_2936),
.Y(n_3522)
);

AOI22xp33_ASAP7_75t_L g3523 ( 
.A1(n_3349),
.A2(n_3364),
.B1(n_3327),
.B2(n_3362),
.Y(n_3523)
);

NOR2xp33_ASAP7_75t_SL g3524 ( 
.A(n_3437),
.B(n_2796),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3151),
.Y(n_3525)
);

NOR2xp33_ASAP7_75t_L g3526 ( 
.A(n_3223),
.B(n_1890),
.Y(n_3526)
);

INVx1_ASAP7_75t_L g3527 ( 
.A(n_3167),
.Y(n_3527)
);

NOR2xp33_ASAP7_75t_L g3528 ( 
.A(n_3223),
.B(n_2901),
.Y(n_3528)
);

NOR2xp33_ASAP7_75t_L g3529 ( 
.A(n_3236),
.B(n_2858),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_3153),
.Y(n_3530)
);

INVx4_ASAP7_75t_L g3531 ( 
.A(n_3232),
.Y(n_3531)
);

AND3x1_ASAP7_75t_SL g3532 ( 
.A(n_3180),
.B(n_3088),
.C(n_1029),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3170),
.Y(n_3533)
);

BUFx4f_ASAP7_75t_SL g3534 ( 
.A(n_3445),
.Y(n_3534)
);

INVx3_ASAP7_75t_L g3535 ( 
.A(n_3232),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_3142),
.B(n_2858),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3176),
.Y(n_3537)
);

HB1xp67_ASAP7_75t_L g3538 ( 
.A(n_3399),
.Y(n_3538)
);

AOI22xp33_ASAP7_75t_L g3539 ( 
.A1(n_3349),
.A2(n_2885),
.B1(n_2876),
.B2(n_2794),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_3161),
.Y(n_3540)
);

HB1xp67_ASAP7_75t_L g3541 ( 
.A(n_3235),
.Y(n_3541)
);

BUFx2_ASAP7_75t_L g3542 ( 
.A(n_3317),
.Y(n_3542)
);

INVx2_ASAP7_75t_SL g3543 ( 
.A(n_3317),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_SL g3544 ( 
.A(n_3145),
.B(n_3093),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_SL g3545 ( 
.A(n_3145),
.B(n_3093),
.Y(n_3545)
);

AOI22xp5_ASAP7_75t_L g3546 ( 
.A1(n_3446),
.A2(n_3110),
.B1(n_2885),
.B2(n_2876),
.Y(n_3546)
);

NAND2x2_ASAP7_75t_L g3547 ( 
.A(n_3143),
.B(n_2980),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_L g3548 ( 
.A(n_3144),
.B(n_2797),
.Y(n_3548)
);

AND2x4_ASAP7_75t_L g3549 ( 
.A(n_3355),
.B(n_2797),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3190),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_SL g3551 ( 
.A(n_3144),
.B(n_3122),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_SL g3552 ( 
.A(n_3191),
.B(n_3156),
.Y(n_3552)
);

NAND2xp33_ASAP7_75t_L g3553 ( 
.A(n_3264),
.B(n_2998),
.Y(n_3553)
);

AOI22xp33_ASAP7_75t_SL g3554 ( 
.A1(n_3483),
.A2(n_2794),
.B1(n_2876),
.B2(n_3003),
.Y(n_3554)
);

NAND3xp33_ASAP7_75t_SL g3555 ( 
.A(n_3446),
.B(n_890),
.C(n_886),
.Y(n_3555)
);

NOR2xp33_ASAP7_75t_L g3556 ( 
.A(n_3236),
.B(n_2992),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3196),
.Y(n_3557)
);

AND2x2_ASAP7_75t_L g3558 ( 
.A(n_3154),
.B(n_3003),
.Y(n_3558)
);

OR2x6_ASAP7_75t_L g3559 ( 
.A(n_3355),
.B(n_3131),
.Y(n_3559)
);

AOI22xp33_ASAP7_75t_L g3560 ( 
.A1(n_3364),
.A2(n_2876),
.B1(n_2794),
.B2(n_2892),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3198),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_3233),
.B(n_2743),
.Y(n_3562)
);

INVx2_ASAP7_75t_L g3563 ( 
.A(n_3181),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_3240),
.B(n_2754),
.Y(n_3564)
);

AND2x4_ASAP7_75t_L g3565 ( 
.A(n_3172),
.B(n_3075),
.Y(n_3565)
);

INVx2_ASAP7_75t_L g3566 ( 
.A(n_3200),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3212),
.Y(n_3567)
);

INVx2_ASAP7_75t_L g3568 ( 
.A(n_3214),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_SL g3569 ( 
.A(n_3158),
.B(n_3122),
.Y(n_3569)
);

AND2x6_ASAP7_75t_SL g3570 ( 
.A(n_3271),
.B(n_3410),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3238),
.B(n_2757),
.Y(n_3571)
);

BUFx3_ASAP7_75t_L g3572 ( 
.A(n_3216),
.Y(n_3572)
);

INVx2_ASAP7_75t_SL g3573 ( 
.A(n_3337),
.Y(n_3573)
);

OAI21xp5_ASAP7_75t_L g3574 ( 
.A1(n_3202),
.A2(n_3120),
.B(n_3006),
.Y(n_3574)
);

INVx1_ASAP7_75t_SL g3575 ( 
.A(n_3443),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_3217),
.Y(n_3576)
);

BUFx6f_ASAP7_75t_L g3577 ( 
.A(n_3232),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3219),
.Y(n_3578)
);

OAI22xp5_ASAP7_75t_L g3579 ( 
.A1(n_3287),
.A2(n_3006),
.B1(n_2921),
.B2(n_2928),
.Y(n_3579)
);

INVx5_ASAP7_75t_L g3580 ( 
.A(n_3221),
.Y(n_3580)
);

HB1xp67_ASAP7_75t_L g3581 ( 
.A(n_3370),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_SL g3582 ( 
.A(n_3157),
.B(n_3271),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3224),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3237),
.Y(n_3584)
);

AOI22xp33_ASAP7_75t_L g3585 ( 
.A1(n_3279),
.A2(n_2794),
.B1(n_2892),
.B2(n_3052),
.Y(n_3585)
);

NOR2xp33_ASAP7_75t_L g3586 ( 
.A(n_3149),
.B(n_3128),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3268),
.Y(n_3587)
);

INVx2_ASAP7_75t_L g3588 ( 
.A(n_3226),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_SL g3589 ( 
.A(n_3358),
.B(n_2737),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3238),
.B(n_3020),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_3230),
.Y(n_3591)
);

A2O1A1Ixp33_ASAP7_75t_L g3592 ( 
.A1(n_3243),
.A2(n_2921),
.B(n_2928),
.C(n_2852),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_3242),
.B(n_3020),
.Y(n_3593)
);

INVx2_ASAP7_75t_L g3594 ( 
.A(n_3246),
.Y(n_3594)
);

NAND2x1p5_ASAP7_75t_L g3595 ( 
.A(n_3249),
.B(n_2737),
.Y(n_3595)
);

OAI21xp33_ASAP7_75t_L g3596 ( 
.A1(n_3220),
.A2(n_898),
.B(n_894),
.Y(n_3596)
);

NOR3xp33_ASAP7_75t_SL g3597 ( 
.A(n_3307),
.B(n_900),
.C(n_899),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3272),
.Y(n_3598)
);

INVx2_ASAP7_75t_L g3599 ( 
.A(n_3255),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_3275),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3289),
.Y(n_3601)
);

INVxp67_ASAP7_75t_L g3602 ( 
.A(n_3306),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_3242),
.B(n_3037),
.Y(n_3603)
);

INVx2_ASAP7_75t_SL g3604 ( 
.A(n_3415),
.Y(n_3604)
);

INVx2_ASAP7_75t_L g3605 ( 
.A(n_3293),
.Y(n_3605)
);

AND2x4_ASAP7_75t_SL g3606 ( 
.A(n_3172),
.B(n_3037),
.Y(n_3606)
);

INVx4_ASAP7_75t_L g3607 ( 
.A(n_3232),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3259),
.B(n_2737),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_SL g3609 ( 
.A(n_3367),
.B(n_2746),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3296),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_L g3611 ( 
.A(n_3259),
.B(n_2746),
.Y(n_3611)
);

INVx2_ASAP7_75t_SL g3612 ( 
.A(n_3486),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3309),
.Y(n_3613)
);

AND2x4_ASAP7_75t_L g3614 ( 
.A(n_3291),
.B(n_2746),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3313),
.Y(n_3615)
);

NOR2xp33_ASAP7_75t_L g3616 ( 
.A(n_3260),
.B(n_2952),
.Y(n_3616)
);

NOR2xp33_ASAP7_75t_L g3617 ( 
.A(n_3260),
.B(n_2210),
.Y(n_3617)
);

BUFx6f_ASAP7_75t_L g3618 ( 
.A(n_3377),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_L g3619 ( 
.A(n_3225),
.B(n_2998),
.Y(n_3619)
);

NAND2x1p5_ASAP7_75t_L g3620 ( 
.A(n_3282),
.B(n_2845),
.Y(n_3620)
);

INVx5_ASAP7_75t_L g3621 ( 
.A(n_3221),
.Y(n_3621)
);

AOI22xp5_ASAP7_75t_L g3622 ( 
.A1(n_3175),
.A2(n_2917),
.B1(n_2892),
.B2(n_2998),
.Y(n_3622)
);

AND2x4_ASAP7_75t_L g3623 ( 
.A(n_3291),
.B(n_3092),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_SL g3624 ( 
.A(n_3389),
.B(n_2996),
.Y(n_3624)
);

AOI22xp5_ASAP7_75t_L g3625 ( 
.A1(n_3175),
.A2(n_2892),
.B1(n_3084),
.B2(n_3023),
.Y(n_3625)
);

AOI22xp5_ASAP7_75t_L g3626 ( 
.A1(n_3178),
.A2(n_3023),
.B1(n_3084),
.B2(n_2951),
.Y(n_3626)
);

BUFx8_ASAP7_75t_SL g3627 ( 
.A(n_3357),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3210),
.B(n_3023),
.Y(n_3628)
);

INVx2_ASAP7_75t_L g3629 ( 
.A(n_3297),
.Y(n_3629)
);

AND2x2_ASAP7_75t_L g3630 ( 
.A(n_3141),
.B(n_1512),
.Y(n_3630)
);

AOI22xp5_ASAP7_75t_L g3631 ( 
.A1(n_3178),
.A2(n_3023),
.B1(n_3084),
.B2(n_2951),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_3177),
.B(n_3084),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3192),
.B(n_3057),
.Y(n_3633)
);

INVx3_ASAP7_75t_L g3634 ( 
.A(n_3377),
.Y(n_3634)
);

INVx2_ASAP7_75t_L g3635 ( 
.A(n_3305),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_3227),
.B(n_3063),
.Y(n_3636)
);

INVx5_ASAP7_75t_L g3637 ( 
.A(n_3221),
.Y(n_3637)
);

INVx2_ASAP7_75t_SL g3638 ( 
.A(n_3340),
.Y(n_3638)
);

HB1xp67_ASAP7_75t_L g3639 ( 
.A(n_3204),
.Y(n_3639)
);

INVx2_ASAP7_75t_SL g3640 ( 
.A(n_3203),
.Y(n_3640)
);

AOI22xp5_ASAP7_75t_L g3641 ( 
.A1(n_3264),
.A2(n_2958),
.B1(n_3053),
.B2(n_2920),
.Y(n_3641)
);

AOI22xp5_ASAP7_75t_L g3642 ( 
.A1(n_3360),
.A2(n_3369),
.B1(n_3345),
.B2(n_3166),
.Y(n_3642)
);

BUFx6f_ASAP7_75t_L g3643 ( 
.A(n_3377),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_3147),
.B(n_3066),
.Y(n_3644)
);

INVxp67_ASAP7_75t_L g3645 ( 
.A(n_3306),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_L g3646 ( 
.A(n_3286),
.B(n_3067),
.Y(n_3646)
);

BUFx2_ASAP7_75t_L g3647 ( 
.A(n_3204),
.Y(n_3647)
);

A2O1A1Ixp33_ASAP7_75t_L g3648 ( 
.A1(n_3220),
.A2(n_2913),
.B(n_3098),
.C(n_3079),
.Y(n_3648)
);

NOR2x2_ASAP7_75t_L g3649 ( 
.A(n_3303),
.B(n_2671),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3314),
.Y(n_3650)
);

INVx2_ASAP7_75t_SL g3651 ( 
.A(n_3458),
.Y(n_3651)
);

INVx2_ASAP7_75t_SL g3652 ( 
.A(n_3263),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_SL g3653 ( 
.A(n_3499),
.B(n_3286),
.Y(n_3653)
);

BUFx12f_ASAP7_75t_L g3654 ( 
.A(n_3245),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3329),
.Y(n_3655)
);

AND2x2_ASAP7_75t_L g3656 ( 
.A(n_3334),
.B(n_1513),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3363),
.Y(n_3657)
);

INVx2_ASAP7_75t_L g3658 ( 
.A(n_3315),
.Y(n_3658)
);

INVx2_ASAP7_75t_L g3659 ( 
.A(n_3319),
.Y(n_3659)
);

CKINVDCx5p33_ASAP7_75t_R g3660 ( 
.A(n_3195),
.Y(n_3660)
);

NOR2xp33_ASAP7_75t_L g3661 ( 
.A(n_3171),
.B(n_3103),
.Y(n_3661)
);

A2O1A1Ixp33_ASAP7_75t_L g3662 ( 
.A1(n_3345),
.A2(n_3070),
.B(n_3078),
.C(n_3074),
.Y(n_3662)
);

NOR3xp33_ASAP7_75t_SL g3663 ( 
.A(n_3304),
.B(n_905),
.C(n_903),
.Y(n_3663)
);

HB1xp67_ASAP7_75t_L g3664 ( 
.A(n_3213),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_SL g3665 ( 
.A(n_3499),
.B(n_2996),
.Y(n_3665)
);

INVx5_ASAP7_75t_L g3666 ( 
.A(n_3221),
.Y(n_3666)
);

OAI22xp5_ASAP7_75t_L g3667 ( 
.A1(n_3287),
.A2(n_2910),
.B1(n_2859),
.B2(n_3022),
.Y(n_3667)
);

CKINVDCx5p33_ASAP7_75t_R g3668 ( 
.A(n_3185),
.Y(n_3668)
);

AO22x1_ASAP7_75t_L g3669 ( 
.A1(n_3470),
.A2(n_2925),
.B1(n_2920),
.B2(n_2958),
.Y(n_3669)
);

AND2x4_ASAP7_75t_L g3670 ( 
.A(n_3310),
.B(n_3092),
.Y(n_3670)
);

INVx2_ASAP7_75t_L g3671 ( 
.A(n_3346),
.Y(n_3671)
);

AOI22xp33_ASAP7_75t_SL g3672 ( 
.A1(n_3437),
.A2(n_2925),
.B1(n_2920),
.B2(n_2958),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3371),
.Y(n_3673)
);

NOR2xp33_ASAP7_75t_L g3674 ( 
.A(n_3294),
.B(n_3082),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3379),
.Y(n_3675)
);

NOR2xp33_ASAP7_75t_L g3676 ( 
.A(n_3277),
.B(n_3083),
.Y(n_3676)
);

BUFx4f_ASAP7_75t_L g3677 ( 
.A(n_3377),
.Y(n_3677)
);

INVx2_ASAP7_75t_SL g3678 ( 
.A(n_3339),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_L g3679 ( 
.A(n_3239),
.B(n_3086),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3381),
.Y(n_3680)
);

AOI22xp33_ASAP7_75t_L g3681 ( 
.A1(n_3162),
.A2(n_3108),
.B1(n_3089),
.B2(n_2788),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_3393),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3407),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_SL g3684 ( 
.A(n_3453),
.B(n_2996),
.Y(n_3684)
);

INVx3_ASAP7_75t_L g3685 ( 
.A(n_3221),
.Y(n_3685)
);

INVx2_ASAP7_75t_L g3686 ( 
.A(n_3347),
.Y(n_3686)
);

HB1xp67_ASAP7_75t_L g3687 ( 
.A(n_3213),
.Y(n_3687)
);

BUFx12f_ASAP7_75t_L g3688 ( 
.A(n_3262),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_SL g3689 ( 
.A(n_3308),
.B(n_2996),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_L g3690 ( 
.A(n_3183),
.B(n_2958),
.Y(n_3690)
);

OR2x6_ASAP7_75t_L g3691 ( 
.A(n_3454),
.B(n_2859),
.Y(n_3691)
);

AOI22xp33_ASAP7_75t_L g3692 ( 
.A1(n_3162),
.A2(n_2788),
.B1(n_3073),
.B2(n_3028),
.Y(n_3692)
);

NOR3xp33_ASAP7_75t_SL g3693 ( 
.A(n_3270),
.B(n_907),
.C(n_906),
.Y(n_3693)
);

BUFx6f_ASAP7_75t_L g3694 ( 
.A(n_3310),
.Y(n_3694)
);

BUFx6f_ASAP7_75t_L g3695 ( 
.A(n_3328),
.Y(n_3695)
);

INVx2_ASAP7_75t_L g3696 ( 
.A(n_3383),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3417),
.Y(n_3697)
);

NOR2xp33_ASAP7_75t_L g3698 ( 
.A(n_3218),
.B(n_2910),
.Y(n_3698)
);

INVx2_ASAP7_75t_SL g3699 ( 
.A(n_3479),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_SL g3700 ( 
.A(n_3353),
.B(n_3069),
.Y(n_3700)
);

AND2x2_ASAP7_75t_L g3701 ( 
.A(n_3261),
.B(n_3365),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_L g3702 ( 
.A(n_3278),
.B(n_2925),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_3278),
.B(n_2925),
.Y(n_3703)
);

NAND2xp5_ASAP7_75t_L g3704 ( 
.A(n_3285),
.B(n_2925),
.Y(n_3704)
);

INVx2_ASAP7_75t_L g3705 ( 
.A(n_3385),
.Y(n_3705)
);

OAI22xp5_ASAP7_75t_L g3706 ( 
.A1(n_3500),
.A2(n_3072),
.B1(n_3105),
.B2(n_3022),
.Y(n_3706)
);

AND2x2_ASAP7_75t_L g3707 ( 
.A(n_3330),
.B(n_1514),
.Y(n_3707)
);

BUFx4f_ASAP7_75t_L g3708 ( 
.A(n_3350),
.Y(n_3708)
);

AOI22xp5_ASAP7_75t_L g3709 ( 
.A1(n_3369),
.A2(n_2920),
.B1(n_930),
.B2(n_946),
.Y(n_3709)
);

INVx2_ASAP7_75t_SL g3710 ( 
.A(n_3514),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_3285),
.B(n_2920),
.Y(n_3711)
);

INVx4_ASAP7_75t_L g3712 ( 
.A(n_3328),
.Y(n_3712)
);

HB1xp67_ASAP7_75t_L g3713 ( 
.A(n_3454),
.Y(n_3713)
);

NAND2xp5_ASAP7_75t_L g3714 ( 
.A(n_3298),
.B(n_3137),
.Y(n_3714)
);

NAND2x1p5_ASAP7_75t_L g3715 ( 
.A(n_3163),
.B(n_3069),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3426),
.Y(n_3716)
);

INVx3_ASAP7_75t_L g3717 ( 
.A(n_3375),
.Y(n_3717)
);

BUFx6f_ASAP7_75t_L g3718 ( 
.A(n_3375),
.Y(n_3718)
);

AOI22xp33_ASAP7_75t_SL g3719 ( 
.A1(n_3169),
.A2(n_1029),
.B1(n_1030),
.B2(n_1028),
.Y(n_3719)
);

HB1xp67_ASAP7_75t_L g3720 ( 
.A(n_3481),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_3434),
.Y(n_3721)
);

INVx1_ASAP7_75t_SL g3722 ( 
.A(n_3256),
.Y(n_3722)
);

OAI22xp5_ASAP7_75t_L g3723 ( 
.A1(n_3500),
.A2(n_3072),
.B1(n_3105),
.B2(n_2900),
.Y(n_3723)
);

AND2x4_ASAP7_75t_L g3724 ( 
.A(n_3431),
.B(n_3092),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_SL g3725 ( 
.A(n_3197),
.B(n_3069),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3436),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_3439),
.Y(n_3727)
);

AOI22xp5_ASAP7_75t_L g3728 ( 
.A1(n_3166),
.A2(n_935),
.B1(n_952),
.B2(n_917),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_3298),
.B(n_3199),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_3441),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_SL g3731 ( 
.A(n_3378),
.B(n_3069),
.Y(n_3731)
);

AOI22xp5_ASAP7_75t_L g3732 ( 
.A1(n_3222),
.A2(n_937),
.B1(n_957),
.B2(n_919),
.Y(n_3732)
);

AOI22xp5_ASAP7_75t_L g3733 ( 
.A1(n_3253),
.A2(n_941),
.B1(n_964),
.B2(n_921),
.Y(n_3733)
);

AOI22xp5_ASAP7_75t_SL g3734 ( 
.A1(n_3288),
.A2(n_1039),
.B1(n_1040),
.B2(n_1038),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_L g3735 ( 
.A(n_3179),
.B(n_3077),
.Y(n_3735)
);

AOI22xp33_ASAP7_75t_L g3736 ( 
.A1(n_3419),
.A2(n_2788),
.B1(n_3118),
.B2(n_3102),
.Y(n_3736)
);

INVx5_ASAP7_75t_L g3737 ( 
.A(n_3375),
.Y(n_3737)
);

INVx2_ASAP7_75t_SL g3738 ( 
.A(n_3374),
.Y(n_3738)
);

AOI22xp5_ASAP7_75t_L g3739 ( 
.A1(n_3380),
.A2(n_945),
.B1(n_970),
.B2(n_924),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3442),
.Y(n_3740)
);

BUFx2_ASAP7_75t_L g3741 ( 
.A(n_3404),
.Y(n_3741)
);

INVx2_ASAP7_75t_L g3742 ( 
.A(n_3403),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3444),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3455),
.Y(n_3744)
);

BUFx3_ASAP7_75t_L g3745 ( 
.A(n_3265),
.Y(n_3745)
);

INVx4_ASAP7_75t_L g3746 ( 
.A(n_3375),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_L g3747 ( 
.A(n_3257),
.B(n_3123),
.Y(n_3747)
);

NAND2xp5_ASAP7_75t_SL g3748 ( 
.A(n_3380),
.B(n_3076),
.Y(n_3748)
);

AO22x1_ASAP7_75t_L g3749 ( 
.A1(n_3508),
.A2(n_955),
.B1(n_976),
.B2(n_925),
.Y(n_3749)
);

OAI21xp33_ASAP7_75t_L g3750 ( 
.A1(n_3174),
.A2(n_910),
.B(n_909),
.Y(n_3750)
);

NAND2xp33_ASAP7_75t_L g3751 ( 
.A(n_3301),
.B(n_3076),
.Y(n_3751)
);

BUFx8_ASAP7_75t_L g3752 ( 
.A(n_3414),
.Y(n_3752)
);

NAND2xp5_ASAP7_75t_L g3753 ( 
.A(n_3311),
.B(n_3139),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_SL g3754 ( 
.A(n_3247),
.B(n_3076),
.Y(n_3754)
);

NOR2x1_ASAP7_75t_L g3755 ( 
.A(n_3406),
.B(n_2756),
.Y(n_3755)
);

NAND2xp5_ASAP7_75t_L g3756 ( 
.A(n_3159),
.B(n_2900),
.Y(n_3756)
);

NOR2xp33_ASAP7_75t_L g3757 ( 
.A(n_3316),
.B(n_2890),
.Y(n_3757)
);

NOR2x1p5_ASAP7_75t_L g3758 ( 
.A(n_3351),
.B(n_2890),
.Y(n_3758)
);

INVx2_ASAP7_75t_L g3759 ( 
.A(n_3405),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_3472),
.Y(n_3760)
);

BUFx2_ASAP7_75t_L g3761 ( 
.A(n_3481),
.Y(n_3761)
);

NAND3xp33_ASAP7_75t_SL g3762 ( 
.A(n_3209),
.B(n_914),
.C(n_911),
.Y(n_3762)
);

AOI21xp5_ASAP7_75t_L g3763 ( 
.A1(n_3359),
.A2(n_2961),
.B(n_3076),
.Y(n_3763)
);

HB1xp67_ASAP7_75t_L g3764 ( 
.A(n_3160),
.Y(n_3764)
);

INVx2_ASAP7_75t_L g3765 ( 
.A(n_3418),
.Y(n_3765)
);

INVx2_ASAP7_75t_L g3766 ( 
.A(n_3427),
.Y(n_3766)
);

INVx2_ASAP7_75t_L g3767 ( 
.A(n_3463),
.Y(n_3767)
);

BUFx5_ASAP7_75t_L g3768 ( 
.A(n_3375),
.Y(n_3768)
);

INVx2_ASAP7_75t_L g3769 ( 
.A(n_3465),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_3254),
.B(n_2931),
.Y(n_3770)
);

INVx2_ASAP7_75t_L g3771 ( 
.A(n_3466),
.Y(n_3771)
);

INVx8_ASAP7_75t_L g3772 ( 
.A(n_3299),
.Y(n_3772)
);

OR2x6_ASAP7_75t_L g3773 ( 
.A(n_3397),
.B(n_2923),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_3228),
.B(n_2931),
.Y(n_3774)
);

AOI22xp33_ASAP7_75t_L g3775 ( 
.A1(n_3457),
.A2(n_2427),
.B1(n_2504),
.B2(n_2503),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3476),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3490),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_3189),
.B(n_2938),
.Y(n_3778)
);

HB1xp67_ASAP7_75t_L g3779 ( 
.A(n_3267),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_3150),
.B(n_2938),
.Y(n_3780)
);

AOI22xp33_ASAP7_75t_L g3781 ( 
.A1(n_3229),
.A2(n_2509),
.B1(n_2526),
.B2(n_2507),
.Y(n_3781)
);

NAND2xp5_ASAP7_75t_L g3782 ( 
.A(n_3152),
.B(n_2954),
.Y(n_3782)
);

NAND2xp5_ASAP7_75t_L g3783 ( 
.A(n_3155),
.B(n_2954),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_SL g3784 ( 
.A(n_3251),
.B(n_2756),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_SL g3785 ( 
.A(n_3276),
.B(n_2808),
.Y(n_3785)
);

INVx2_ASAP7_75t_SL g3786 ( 
.A(n_3164),
.Y(n_3786)
);

OAI21xp33_ASAP7_75t_L g3787 ( 
.A1(n_3280),
.A2(n_927),
.B(n_926),
.Y(n_3787)
);

OAI22x1_ASAP7_75t_R g3788 ( 
.A1(n_3400),
.A2(n_936),
.B1(n_939),
.B2(n_929),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_L g3789 ( 
.A(n_3186),
.B(n_2981),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_L g3790 ( 
.A(n_3729),
.B(n_3582),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_SL g3791 ( 
.A(n_3642),
.B(n_3732),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_SL g3792 ( 
.A(n_3642),
.B(n_3326),
.Y(n_3792)
);

NAND2xp33_ASAP7_75t_SL g3793 ( 
.A(n_3668),
.B(n_3266),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_SL g3794 ( 
.A(n_3732),
.B(n_3326),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_SL g3795 ( 
.A(n_3653),
.B(n_3276),
.Y(n_3795)
);

NAND2xp33_ASAP7_75t_SL g3796 ( 
.A(n_3571),
.B(n_3408),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_SL g3797 ( 
.A(n_3706),
.B(n_3356),
.Y(n_3797)
);

NAND2xp33_ASAP7_75t_SL g3798 ( 
.A(n_3693),
.B(n_3173),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_SL g3799 ( 
.A(n_3579),
.B(n_3361),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_SL g3800 ( 
.A(n_3579),
.B(n_3372),
.Y(n_3800)
);

NAND2xp5_ASAP7_75t_SL g3801 ( 
.A(n_3552),
.B(n_3384),
.Y(n_3801)
);

NAND2xp5_ASAP7_75t_SL g3802 ( 
.A(n_3723),
.B(n_3451),
.Y(n_3802)
);

NAND2xp5_ASAP7_75t_SL g3803 ( 
.A(n_3616),
.B(n_3373),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_SL g3804 ( 
.A(n_3702),
.B(n_3433),
.Y(n_3804)
);

AND2x2_ASAP7_75t_L g3805 ( 
.A(n_3701),
.B(n_3412),
.Y(n_3805)
);

NAND2xp5_ASAP7_75t_SL g3806 ( 
.A(n_3548),
.B(n_3447),
.Y(n_3806)
);

NAND2xp5_ASAP7_75t_L g3807 ( 
.A(n_3602),
.B(n_3491),
.Y(n_3807)
);

NAND2xp33_ASAP7_75t_SL g3808 ( 
.A(n_3712),
.B(n_3182),
.Y(n_3808)
);

NAND2xp5_ASAP7_75t_SL g3809 ( 
.A(n_3529),
.B(n_3528),
.Y(n_3809)
);

AND2x2_ASAP7_75t_L g3810 ( 
.A(n_3541),
.B(n_3312),
.Y(n_3810)
);

NAND2xp33_ASAP7_75t_SL g3811 ( 
.A(n_3712),
.B(n_3184),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_SL g3812 ( 
.A(n_3590),
.B(n_3447),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_L g3813 ( 
.A(n_3645),
.B(n_3526),
.Y(n_3813)
);

AND2x2_ASAP7_75t_L g3814 ( 
.A(n_3656),
.B(n_3312),
.Y(n_3814)
);

NAND2xp33_ASAP7_75t_SL g3815 ( 
.A(n_3597),
.B(n_3165),
.Y(n_3815)
);

NAND2xp33_ASAP7_75t_SL g3816 ( 
.A(n_3663),
.B(n_3258),
.Y(n_3816)
);

NAND2xp33_ASAP7_75t_SL g3817 ( 
.A(n_3660),
.B(n_3244),
.Y(n_3817)
);

NAND2xp5_ASAP7_75t_SL g3818 ( 
.A(n_3593),
.B(n_3209),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_SL g3819 ( 
.A(n_3603),
.B(n_3510),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3646),
.B(n_3498),
.Y(n_3820)
);

AND2x4_ASAP7_75t_L g3821 ( 
.A(n_3559),
.B(n_3438),
.Y(n_3821)
);

NAND2xp5_ASAP7_75t_SL g3822 ( 
.A(n_3556),
.B(n_3622),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_SL g3823 ( 
.A(n_3622),
.B(n_3608),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_SL g3824 ( 
.A(n_3611),
.B(n_3510),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_L g3825 ( 
.A(n_3779),
.B(n_3503),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_SL g3826 ( 
.A(n_3661),
.B(n_3194),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_SL g3827 ( 
.A(n_3626),
.B(n_3631),
.Y(n_3827)
);

NAND2xp5_ASAP7_75t_L g3828 ( 
.A(n_3581),
.B(n_3390),
.Y(n_3828)
);

AND2x2_ASAP7_75t_L g3829 ( 
.A(n_3707),
.B(n_3193),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_SL g3830 ( 
.A(n_3626),
.B(n_3194),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_L g3831 ( 
.A(n_3562),
.B(n_3504),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_SL g3832 ( 
.A(n_3631),
.B(n_3284),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_SL g3833 ( 
.A(n_3625),
.B(n_3188),
.Y(n_3833)
);

NAND2xp5_ASAP7_75t_SL g3834 ( 
.A(n_3625),
.B(n_3188),
.Y(n_3834)
);

NAND2xp5_ASAP7_75t_L g3835 ( 
.A(n_3722),
.B(n_3509),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_SL g3836 ( 
.A(n_3676),
.B(n_3283),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_SL g3837 ( 
.A(n_3703),
.B(n_3273),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_SL g3838 ( 
.A(n_3704),
.B(n_3273),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_L g3839 ( 
.A(n_3722),
.B(n_3630),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_SL g3840 ( 
.A(n_3711),
.B(n_3709),
.Y(n_3840)
);

NAND2xp33_ASAP7_75t_SL g3841 ( 
.A(n_3640),
.B(n_3234),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_SL g3842 ( 
.A(n_3709),
.B(n_3168),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_SL g3843 ( 
.A(n_3674),
.B(n_3435),
.Y(n_3843)
);

NAND2xp5_ASAP7_75t_SL g3844 ( 
.A(n_3544),
.B(n_3440),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_SL g3845 ( 
.A(n_3545),
.B(n_3449),
.Y(n_3845)
);

NAND2xp5_ASAP7_75t_SL g3846 ( 
.A(n_3521),
.B(n_3462),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_SL g3847 ( 
.A(n_3536),
.B(n_3464),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_SL g3848 ( 
.A(n_3546),
.B(n_3229),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_SL g3849 ( 
.A(n_3546),
.B(n_3146),
.Y(n_3849)
);

NAND2xp33_ASAP7_75t_SL g3850 ( 
.A(n_3694),
.B(n_3391),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_SL g3851 ( 
.A(n_3698),
.B(n_3524),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_SL g3852 ( 
.A(n_3524),
.B(n_3338),
.Y(n_3852)
);

NAND2xp5_ASAP7_75t_SL g3853 ( 
.A(n_3714),
.B(n_3338),
.Y(n_3853)
);

NAND2xp33_ASAP7_75t_SL g3854 ( 
.A(n_3694),
.B(n_3394),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_SL g3855 ( 
.A(n_3619),
.B(n_3507),
.Y(n_3855)
);

NAND2xp5_ASAP7_75t_L g3856 ( 
.A(n_3633),
.B(n_3515),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_SL g3857 ( 
.A(n_3554),
.B(n_3507),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_SL g3858 ( 
.A(n_3551),
.B(n_3475),
.Y(n_3858)
);

NAND2xp5_ASAP7_75t_SL g3859 ( 
.A(n_3522),
.B(n_3475),
.Y(n_3859)
);

AND2x2_ASAP7_75t_L g3860 ( 
.A(n_3558),
.B(n_3215),
.Y(n_3860)
);

NAND2xp33_ASAP7_75t_SL g3861 ( 
.A(n_3694),
.B(n_3250),
.Y(n_3861)
);

AND2x2_ASAP7_75t_L g3862 ( 
.A(n_3647),
.B(n_3342),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_SL g3863 ( 
.A(n_3580),
.B(n_3342),
.Y(n_3863)
);

NAND2xp33_ASAP7_75t_SL g3864 ( 
.A(n_3695),
.B(n_3411),
.Y(n_3864)
);

AND2x2_ASAP7_75t_L g3865 ( 
.A(n_3761),
.B(n_3431),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_SL g3866 ( 
.A(n_3580),
.B(n_3448),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_SL g3867 ( 
.A(n_3580),
.B(n_3448),
.Y(n_3867)
);

AND2x2_ASAP7_75t_SL g3868 ( 
.A(n_3553),
.B(n_3343),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_SL g3869 ( 
.A(n_3621),
.B(n_3290),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_SL g3870 ( 
.A(n_3621),
.B(n_3292),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_SL g3871 ( 
.A(n_3621),
.B(n_3489),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_SL g3872 ( 
.A(n_3637),
.B(n_3489),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_3764),
.B(n_3469),
.Y(n_3873)
);

NAND2xp33_ASAP7_75t_SL g3874 ( 
.A(n_3695),
.B(n_3488),
.Y(n_3874)
);

NAND2xp5_ASAP7_75t_SL g3875 ( 
.A(n_3637),
.B(n_3274),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_L g3876 ( 
.A(n_3678),
.B(n_3469),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_SL g3877 ( 
.A(n_3637),
.B(n_3321),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_L g3878 ( 
.A(n_3636),
.B(n_3639),
.Y(n_3878)
);

AND2x4_ASAP7_75t_L g3879 ( 
.A(n_3559),
.B(n_3438),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_SL g3880 ( 
.A(n_3666),
.B(n_3331),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_L g3881 ( 
.A(n_3664),
.B(n_3320),
.Y(n_3881)
);

NAND2xp33_ASAP7_75t_SL g3882 ( 
.A(n_3695),
.B(n_3492),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_SL g3883 ( 
.A(n_3666),
.B(n_3332),
.Y(n_3883)
);

NAND2xp33_ASAP7_75t_SL g3884 ( 
.A(n_3687),
.B(n_3423),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_L g3885 ( 
.A(n_3713),
.B(n_3252),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_SL g3886 ( 
.A(n_3666),
.B(n_3366),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_SL g3887 ( 
.A(n_3737),
.B(n_3366),
.Y(n_3887)
);

NAND2xp33_ASAP7_75t_SL g3888 ( 
.A(n_3746),
.B(n_3424),
.Y(n_3888)
);

NAND2xp5_ASAP7_75t_SL g3889 ( 
.A(n_3737),
.B(n_3366),
.Y(n_3889)
);

NAND2xp5_ASAP7_75t_SL g3890 ( 
.A(n_3737),
.B(n_3366),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_SL g3891 ( 
.A(n_3560),
.B(n_3366),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_SL g3892 ( 
.A(n_3628),
.B(n_3366),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_L g3893 ( 
.A(n_3720),
.B(n_3281),
.Y(n_3893)
);

NAND2xp33_ASAP7_75t_SL g3894 ( 
.A(n_3746),
.B(n_3425),
.Y(n_3894)
);

NAND2xp5_ASAP7_75t_SL g3895 ( 
.A(n_3585),
.B(n_3480),
.Y(n_3895)
);

NAND2xp33_ASAP7_75t_SL g3896 ( 
.A(n_3741),
.B(n_3430),
.Y(n_3896)
);

NAND2xp5_ASAP7_75t_SL g3897 ( 
.A(n_3719),
.B(n_3480),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_SL g3898 ( 
.A(n_3677),
.B(n_3480),
.Y(n_3898)
);

NAND2xp33_ASAP7_75t_SL g3899 ( 
.A(n_3718),
.B(n_3538),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_SL g3900 ( 
.A(n_3677),
.B(n_3480),
.Y(n_3900)
);

NAND2xp5_ASAP7_75t_SL g3901 ( 
.A(n_3728),
.B(n_3480),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_SL g3902 ( 
.A(n_3728),
.B(n_3480),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_SL g3903 ( 
.A(n_3641),
.B(n_3395),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_SL g3904 ( 
.A(n_3641),
.B(n_3352),
.Y(n_3904)
);

NAND2xp33_ASAP7_75t_SL g3905 ( 
.A(n_3718),
.B(n_3207),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_SL g3906 ( 
.A(n_3718),
.B(n_3336),
.Y(n_3906)
);

NAND2xp33_ASAP7_75t_SL g3907 ( 
.A(n_3604),
.B(n_3231),
.Y(n_3907)
);

AND2x4_ASAP7_75t_L g3908 ( 
.A(n_3559),
.B(n_3205),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_SL g3909 ( 
.A(n_3586),
.B(n_3344),
.Y(n_3909)
);

NAND2xp5_ASAP7_75t_SL g3910 ( 
.A(n_3574),
.B(n_3456),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_L g3911 ( 
.A(n_3644),
.B(n_3456),
.Y(n_3911)
);

NAND2xp33_ASAP7_75t_SL g3912 ( 
.A(n_3542),
.B(n_3241),
.Y(n_3912)
);

NAND2xp5_ASAP7_75t_SL g3913 ( 
.A(n_3574),
.B(n_3459),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_SL g3914 ( 
.A(n_3665),
.B(n_3672),
.Y(n_3914)
);

NAND2xp33_ASAP7_75t_SL g3915 ( 
.A(n_3543),
.B(n_3396),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_SL g3916 ( 
.A(n_3617),
.B(n_3459),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_SL g3917 ( 
.A(n_3734),
.B(n_3467),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_SL g3918 ( 
.A(n_3734),
.B(n_3467),
.Y(n_3918)
);

NAND2xp5_ASAP7_75t_SL g3919 ( 
.A(n_3569),
.B(n_3318),
.Y(n_3919)
);

NAND2xp5_ASAP7_75t_SL g3920 ( 
.A(n_3757),
.B(n_3322),
.Y(n_3920)
);

NAND2xp33_ASAP7_75t_SL g3921 ( 
.A(n_3786),
.B(n_3382),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_L g3922 ( 
.A(n_3564),
.B(n_3485),
.Y(n_3922)
);

NAND2xp33_ASAP7_75t_SL g3923 ( 
.A(n_3651),
.B(n_3402),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_SL g3924 ( 
.A(n_3679),
.B(n_3269),
.Y(n_3924)
);

NAND2xp5_ASAP7_75t_SL g3925 ( 
.A(n_3539),
.B(n_3474),
.Y(n_3925)
);

NAND2xp33_ASAP7_75t_SL g3926 ( 
.A(n_3623),
.B(n_3670),
.Y(n_3926)
);

NAND2xp5_ASAP7_75t_SL g3927 ( 
.A(n_3577),
.B(n_3474),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_SL g3928 ( 
.A(n_3577),
.B(n_3368),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_SL g3929 ( 
.A(n_3577),
.B(n_2781),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_SL g3930 ( 
.A(n_3618),
.B(n_2781),
.Y(n_3930)
);

NAND2xp5_ASAP7_75t_SL g3931 ( 
.A(n_3618),
.B(n_2781),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_L g3932 ( 
.A(n_3747),
.B(n_3473),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_SL g3933 ( 
.A(n_3618),
.B(n_2828),
.Y(n_3933)
);

AND2x2_ASAP7_75t_SL g3934 ( 
.A(n_3523),
.B(n_3392),
.Y(n_3934)
);

NAND2xp33_ASAP7_75t_SL g3935 ( 
.A(n_3623),
.B(n_3505),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_L g3936 ( 
.A(n_3770),
.B(n_3477),
.Y(n_3936)
);

NAND2xp5_ASAP7_75t_SL g3937 ( 
.A(n_3643),
.B(n_3690),
.Y(n_3937)
);

NAND2xp5_ASAP7_75t_SL g3938 ( 
.A(n_3643),
.B(n_2828),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_SL g3939 ( 
.A(n_3643),
.B(n_3648),
.Y(n_3939)
);

NAND2xp5_ASAP7_75t_SL g3940 ( 
.A(n_3632),
.B(n_2828),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_SL g3941 ( 
.A(n_3755),
.B(n_2838),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_SL g3942 ( 
.A(n_3575),
.B(n_2838),
.Y(n_3942)
);

AND2x2_ASAP7_75t_L g3943 ( 
.A(n_3575),
.B(n_3333),
.Y(n_3943)
);

NAND2xp5_ASAP7_75t_SL g3944 ( 
.A(n_3774),
.B(n_2838),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_SL g3945 ( 
.A(n_3785),
.B(n_2864),
.Y(n_3945)
);

NAND2xp33_ASAP7_75t_SL g3946 ( 
.A(n_3670),
.B(n_3211),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_SL g3947 ( 
.A(n_3662),
.B(n_2864),
.Y(n_3947)
);

AND3x1_ASAP7_75t_L g3948 ( 
.A(n_3638),
.B(n_1039),
.C(n_1038),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_SL g3949 ( 
.A(n_3778),
.B(n_2864),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_L g3950 ( 
.A(n_3753),
.B(n_3478),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_SL g3951 ( 
.A(n_3750),
.B(n_2877),
.Y(n_3951)
);

AND2x2_ASAP7_75t_L g3952 ( 
.A(n_3710),
.B(n_1040),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3525),
.B(n_3482),
.Y(n_3953)
);

AND2x2_ASAP7_75t_L g3954 ( 
.A(n_3699),
.B(n_1043),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_L g3955 ( 
.A(n_3527),
.B(n_3487),
.Y(n_3955)
);

NAND2xp33_ASAP7_75t_SL g3956 ( 
.A(n_3573),
.B(n_3565),
.Y(n_3956)
);

NAND2xp5_ASAP7_75t_L g3957 ( 
.A(n_3533),
.B(n_3376),
.Y(n_3957)
);

NAND2xp33_ASAP7_75t_SL g3958 ( 
.A(n_3565),
.B(n_3211),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_SL g3959 ( 
.A(n_3750),
.B(n_3549),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_SL g3960 ( 
.A(n_3549),
.B(n_2877),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_SL g3961 ( 
.A(n_3535),
.B(n_2877),
.Y(n_3961)
);

NAND2xp33_ASAP7_75t_SL g3962 ( 
.A(n_3738),
.B(n_3468),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_SL g3963 ( 
.A(n_3535),
.B(n_2886),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_L g3964 ( 
.A(n_3537),
.B(n_3550),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_SL g3965 ( 
.A(n_3634),
.B(n_2886),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_L g3966 ( 
.A(n_3557),
.B(n_3295),
.Y(n_3966)
);

NAND2xp5_ASAP7_75t_L g3967 ( 
.A(n_3561),
.B(n_3421),
.Y(n_3967)
);

NAND2xp5_ASAP7_75t_SL g3968 ( 
.A(n_3634),
.B(n_2886),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_SL g3969 ( 
.A(n_3754),
.B(n_2899),
.Y(n_3969)
);

NAND2xp5_ASAP7_75t_SL g3970 ( 
.A(n_3725),
.B(n_2899),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_SL g3971 ( 
.A(n_3789),
.B(n_2899),
.Y(n_3971)
);

NAND2xp5_ASAP7_75t_SL g3972 ( 
.A(n_3787),
.B(n_3531),
.Y(n_3972)
);

NAND2xp33_ASAP7_75t_SL g3973 ( 
.A(n_3612),
.B(n_3468),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_SL g3974 ( 
.A(n_3787),
.B(n_2955),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_SL g3975 ( 
.A(n_3531),
.B(n_2955),
.Y(n_3975)
);

NAND2xp5_ASAP7_75t_SL g3976 ( 
.A(n_3607),
.B(n_2955),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_SL g3977 ( 
.A(n_3607),
.B(n_3685),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_L g3978 ( 
.A(n_3567),
.B(n_3493),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_SL g3979 ( 
.A(n_3685),
.B(n_2956),
.Y(n_3979)
);

NAND2xp33_ASAP7_75t_SL g3980 ( 
.A(n_3758),
.B(n_3484),
.Y(n_3980)
);

NAND2xp5_ASAP7_75t_SL g3981 ( 
.A(n_3717),
.B(n_2956),
.Y(n_3981)
);

NAND2xp33_ASAP7_75t_SL g3982 ( 
.A(n_3717),
.B(n_3484),
.Y(n_3982)
);

NAND2xp33_ASAP7_75t_SL g3983 ( 
.A(n_3652),
.B(n_3495),
.Y(n_3983)
);

NAND2xp33_ASAP7_75t_SL g3984 ( 
.A(n_3614),
.B(n_3495),
.Y(n_3984)
);

NAND2xp5_ASAP7_75t_L g3985 ( 
.A(n_3578),
.B(n_3496),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_3583),
.B(n_3497),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_SL g3987 ( 
.A(n_3684),
.B(n_3700),
.Y(n_3987)
);

NAND2xp5_ASAP7_75t_SL g3988 ( 
.A(n_3596),
.B(n_3667),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_SL g3989 ( 
.A(n_3596),
.B(n_2956),
.Y(n_3989)
);

NAND2xp5_ASAP7_75t_SL g3990 ( 
.A(n_3748),
.B(n_2987),
.Y(n_3990)
);

NAND2xp33_ASAP7_75t_SL g3991 ( 
.A(n_3614),
.B(n_3354),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_SL g3992 ( 
.A(n_3745),
.B(n_2987),
.Y(n_3992)
);

AND2x4_ASAP7_75t_L g3993 ( 
.A(n_3724),
.B(n_3205),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_SL g3994 ( 
.A(n_3624),
.B(n_2987),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_SL g3995 ( 
.A(n_3731),
.B(n_3013),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_SL g3996 ( 
.A(n_3534),
.B(n_3013),
.Y(n_3996)
);

NAND2xp5_ASAP7_75t_SL g3997 ( 
.A(n_3724),
.B(n_3013),
.Y(n_3997)
);

NAND2xp5_ASAP7_75t_SL g3998 ( 
.A(n_3689),
.B(n_3015),
.Y(n_3998)
);

NAND2xp5_ASAP7_75t_SL g3999 ( 
.A(n_3780),
.B(n_3015),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_SL g4000 ( 
.A(n_3782),
.B(n_3015),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_SL g4001 ( 
.A(n_3783),
.B(n_3768),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_SL g4002 ( 
.A(n_3768),
.B(n_3035),
.Y(n_4002)
);

AND2x4_ASAP7_75t_L g4003 ( 
.A(n_3691),
.B(n_3206),
.Y(n_4003)
);

NAND2xp5_ASAP7_75t_SL g4004 ( 
.A(n_3768),
.B(n_3035),
.Y(n_4004)
);

NAND2xp33_ASAP7_75t_SL g4005 ( 
.A(n_3784),
.B(n_2923),
.Y(n_4005)
);

NAND2xp5_ASAP7_75t_SL g4006 ( 
.A(n_3768),
.B(n_3756),
.Y(n_4006)
);

NAND2xp5_ASAP7_75t_SL g4007 ( 
.A(n_3768),
.B(n_3035),
.Y(n_4007)
);

NAND2xp5_ASAP7_75t_SL g4008 ( 
.A(n_3739),
.B(n_3054),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_SL g4009 ( 
.A(n_3739),
.B(n_3054),
.Y(n_4009)
);

NAND2xp5_ASAP7_75t_SL g4010 ( 
.A(n_3736),
.B(n_3054),
.Y(n_4010)
);

NAND2xp5_ASAP7_75t_L g4011 ( 
.A(n_3584),
.B(n_3587),
.Y(n_4011)
);

NAND2xp5_ASAP7_75t_L g4012 ( 
.A(n_3598),
.B(n_3401),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_SL g4013 ( 
.A(n_3733),
.B(n_3056),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_SL g4014 ( 
.A(n_3733),
.B(n_3056),
.Y(n_4014)
);

NAND2xp33_ASAP7_75t_SL g4015 ( 
.A(n_3589),
.B(n_3056),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_SL g4016 ( 
.A(n_3681),
.B(n_3609),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_SL g4017 ( 
.A(n_3620),
.B(n_3094),
.Y(n_4017)
);

NAND2xp5_ASAP7_75t_SL g4018 ( 
.A(n_3592),
.B(n_3094),
.Y(n_4018)
);

AND2x2_ASAP7_75t_L g4019 ( 
.A(n_3595),
.B(n_1043),
.Y(n_4019)
);

NAND2xp33_ASAP7_75t_SL g4020 ( 
.A(n_3520),
.B(n_3094),
.Y(n_4020)
);

NAND2xp5_ASAP7_75t_SL g4021 ( 
.A(n_3735),
.B(n_3106),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_SL g4022 ( 
.A(n_3715),
.B(n_3106),
.Y(n_4022)
);

NAND2xp5_ASAP7_75t_L g4023 ( 
.A(n_3600),
.B(n_3413),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_SL g4024 ( 
.A(n_3519),
.B(n_3106),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_SL g4025 ( 
.A(n_3572),
.B(n_3114),
.Y(n_4025)
);

AND2x2_ASAP7_75t_L g4026 ( 
.A(n_3601),
.B(n_1046),
.Y(n_4026)
);

NAND2xp5_ASAP7_75t_SL g4027 ( 
.A(n_3610),
.B(n_3114),
.Y(n_4027)
);

NAND2xp5_ASAP7_75t_L g4028 ( 
.A(n_3613),
.B(n_3420),
.Y(n_4028)
);

NAND2xp5_ASAP7_75t_SL g4029 ( 
.A(n_3692),
.B(n_3450),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_SL g4030 ( 
.A(n_3763),
.B(n_3429),
.Y(n_4030)
);

AND2x4_ASAP7_75t_L g4031 ( 
.A(n_3691),
.B(n_3206),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_SL g4032 ( 
.A(n_3615),
.B(n_3429),
.Y(n_4032)
);

NAND2xp5_ASAP7_75t_SL g4033 ( 
.A(n_3650),
.B(n_3494),
.Y(n_4033)
);

AND2x2_ASAP7_75t_L g4034 ( 
.A(n_3655),
.B(n_3657),
.Y(n_4034)
);

AND2x2_ASAP7_75t_L g4035 ( 
.A(n_3673),
.B(n_3675),
.Y(n_4035)
);

AND2x2_ASAP7_75t_L g4036 ( 
.A(n_3680),
.B(n_1046),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_SL g4037 ( 
.A(n_3682),
.B(n_3114),
.Y(n_4037)
);

INVx3_ASAP7_75t_L g4038 ( 
.A(n_3865),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_L g4039 ( 
.A(n_3878),
.B(n_3683),
.Y(n_4039)
);

BUFx6f_ASAP7_75t_L g4040 ( 
.A(n_3875),
.Y(n_4040)
);

INVx2_ASAP7_75t_L g4041 ( 
.A(n_4034),
.Y(n_4041)
);

AND2x4_ASAP7_75t_L g4042 ( 
.A(n_3821),
.B(n_3691),
.Y(n_4042)
);

CKINVDCx5p33_ASAP7_75t_R g4043 ( 
.A(n_3841),
.Y(n_4043)
);

AND2x4_ASAP7_75t_L g4044 ( 
.A(n_3821),
.B(n_3697),
.Y(n_4044)
);

INVx1_ASAP7_75t_L g4045 ( 
.A(n_3964),
.Y(n_4045)
);

NAND2xp5_ASAP7_75t_L g4046 ( 
.A(n_3836),
.B(n_3716),
.Y(n_4046)
);

NAND2x1_ASAP7_75t_L g4047 ( 
.A(n_4003),
.B(n_4031),
.Y(n_4047)
);

AND2x2_ASAP7_75t_L g4048 ( 
.A(n_3810),
.B(n_3721),
.Y(n_4048)
);

BUFx6f_ASAP7_75t_L g4049 ( 
.A(n_3997),
.Y(n_4049)
);

BUFx4f_ASAP7_75t_L g4050 ( 
.A(n_3814),
.Y(n_4050)
);

OAI22xp5_ASAP7_75t_L g4051 ( 
.A1(n_3791),
.A2(n_3794),
.B1(n_3792),
.B2(n_3826),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_4011),
.Y(n_4052)
);

AND2x2_ASAP7_75t_L g4053 ( 
.A(n_3862),
.B(n_3805),
.Y(n_4053)
);

INVx3_ASAP7_75t_L g4054 ( 
.A(n_3993),
.Y(n_4054)
);

AND2x2_ASAP7_75t_L g4055 ( 
.A(n_4035),
.B(n_3726),
.Y(n_4055)
);

OAI21xp5_ASAP7_75t_L g4056 ( 
.A1(n_3794),
.A2(n_3762),
.B(n_3555),
.Y(n_4056)
);

BUFx6f_ASAP7_75t_L g4057 ( 
.A(n_3839),
.Y(n_4057)
);

BUFx3_ASAP7_75t_L g4058 ( 
.A(n_3943),
.Y(n_4058)
);

BUFx6f_ASAP7_75t_L g4059 ( 
.A(n_3996),
.Y(n_4059)
);

INVxp67_ASAP7_75t_L g4060 ( 
.A(n_3807),
.Y(n_4060)
);

OAI22xp5_ASAP7_75t_L g4061 ( 
.A1(n_3791),
.A2(n_3547),
.B1(n_3388),
.B2(n_3392),
.Y(n_4061)
);

AOI22xp5_ASAP7_75t_L g4062 ( 
.A1(n_3934),
.A2(n_3532),
.B1(n_3749),
.B2(n_3688),
.Y(n_4062)
);

AO32x1_ASAP7_75t_L g4063 ( 
.A1(n_4026),
.A2(n_3727),
.A3(n_3743),
.B1(n_3740),
.B2(n_3730),
.Y(n_4063)
);

BUFx8_ASAP7_75t_SL g4064 ( 
.A(n_3813),
.Y(n_4064)
);

INVxp67_ASAP7_75t_L g4065 ( 
.A(n_3885),
.Y(n_4065)
);

AND2x4_ASAP7_75t_L g4066 ( 
.A(n_3821),
.B(n_3744),
.Y(n_4066)
);

A2O1A1Ixp33_ASAP7_75t_L g4067 ( 
.A1(n_3792),
.A2(n_3409),
.B(n_3461),
.C(n_3335),
.Y(n_4067)
);

NAND2xp5_ASAP7_75t_L g4068 ( 
.A(n_3893),
.B(n_3760),
.Y(n_4068)
);

OAI22xp33_ASAP7_75t_L g4069 ( 
.A1(n_3848),
.A2(n_3795),
.B1(n_3822),
.B2(n_3833),
.Y(n_4069)
);

NOR2xp33_ASAP7_75t_L g4070 ( 
.A(n_3790),
.B(n_3627),
.Y(n_4070)
);

A2O1A1Ixp33_ASAP7_75t_SL g4071 ( 
.A1(n_3957),
.A2(n_1049),
.B(n_1054),
.C(n_1047),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_L g4072 ( 
.A(n_3828),
.B(n_3776),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_L g4073 ( 
.A(n_3843),
.B(n_3777),
.Y(n_4073)
);

HB1xp67_ASAP7_75t_L g4074 ( 
.A(n_3881),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_L g4075 ( 
.A(n_3820),
.B(n_3570),
.Y(n_4075)
);

NAND2xp5_ASAP7_75t_L g4076 ( 
.A(n_3911),
.B(n_3825),
.Y(n_4076)
);

BUFx6f_ASAP7_75t_L g4077 ( 
.A(n_3960),
.Y(n_4077)
);

AOI22xp33_ASAP7_75t_L g4078 ( 
.A1(n_3934),
.A2(n_3795),
.B1(n_3834),
.B2(n_3925),
.Y(n_4078)
);

AOI22xp33_ASAP7_75t_L g4079 ( 
.A1(n_3830),
.A2(n_3812),
.B1(n_3849),
.B2(n_3806),
.Y(n_4079)
);

INVx2_ASAP7_75t_L g4080 ( 
.A(n_4028),
.Y(n_4080)
);

BUFx8_ASAP7_75t_L g4081 ( 
.A(n_3954),
.Y(n_4081)
);

INVx1_ASAP7_75t_L g4082 ( 
.A(n_3835),
.Y(n_4082)
);

AOI21xp5_ASAP7_75t_L g4083 ( 
.A1(n_3802),
.A2(n_3751),
.B(n_3387),
.Y(n_4083)
);

A2O1A1Ixp33_ASAP7_75t_L g4084 ( 
.A1(n_3798),
.A2(n_3570),
.B(n_3788),
.C(n_3772),
.Y(n_4084)
);

NAND2x2_ASAP7_75t_L g4085 ( 
.A(n_3796),
.B(n_3772),
.Y(n_4085)
);

AND2x2_ASAP7_75t_L g4086 ( 
.A(n_3860),
.B(n_3773),
.Y(n_4086)
);

CKINVDCx5p33_ASAP7_75t_R g4087 ( 
.A(n_3793),
.Y(n_4087)
);

BUFx6f_ASAP7_75t_L g4088 ( 
.A(n_3868),
.Y(n_4088)
);

INVx3_ASAP7_75t_L g4089 ( 
.A(n_3993),
.Y(n_4089)
);

OAI22xp33_ASAP7_75t_L g4090 ( 
.A1(n_3857),
.A2(n_3772),
.B1(n_3654),
.B2(n_3773),
.Y(n_4090)
);

HB1xp67_ASAP7_75t_L g4091 ( 
.A(n_3804),
.Y(n_4091)
);

HB1xp67_ASAP7_75t_L g4092 ( 
.A(n_3804),
.Y(n_4092)
);

INVx2_ASAP7_75t_L g4093 ( 
.A(n_4012),
.Y(n_4093)
);

AND2x4_ASAP7_75t_L g4094 ( 
.A(n_3879),
.B(n_3773),
.Y(n_4094)
);

AOI221xp5_ASAP7_75t_L g4095 ( 
.A1(n_3948),
.A2(n_1054),
.B1(n_1058),
.B2(n_1049),
.C(n_1047),
.Y(n_4095)
);

OAI22xp5_ASAP7_75t_L g4096 ( 
.A1(n_3903),
.A2(n_3708),
.B1(n_3416),
.B2(n_3324),
.Y(n_4096)
);

INVx4_ASAP7_75t_L g4097 ( 
.A(n_3868),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_SL g4098 ( 
.A(n_3817),
.B(n_3708),
.Y(n_4098)
);

CKINVDCx5p33_ASAP7_75t_R g4099 ( 
.A(n_3912),
.Y(n_4099)
);

A2O1A1Ixp33_ASAP7_75t_L g4100 ( 
.A1(n_3988),
.A2(n_3302),
.B(n_3606),
.C(n_1063),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3966),
.Y(n_4101)
);

BUFx8_ASAP7_75t_SL g4102 ( 
.A(n_3829),
.Y(n_4102)
);

INVx2_ASAP7_75t_L g4103 ( 
.A(n_4023),
.Y(n_4103)
);

NAND2xp5_ASAP7_75t_L g4104 ( 
.A(n_3831),
.B(n_3518),
.Y(n_4104)
);

NAND2xp5_ASAP7_75t_SL g4105 ( 
.A(n_3896),
.B(n_3752),
.Y(n_4105)
);

AND2x2_ASAP7_75t_L g4106 ( 
.A(n_3809),
.B(n_1058),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_L g4107 ( 
.A(n_3856),
.B(n_3530),
.Y(n_4107)
);

NAND2xp5_ASAP7_75t_SL g4108 ( 
.A(n_3915),
.B(n_3752),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_L g4109 ( 
.A(n_3936),
.B(n_3540),
.Y(n_4109)
);

BUFx2_ASAP7_75t_L g4110 ( 
.A(n_3907),
.Y(n_4110)
);

HB1xp67_ASAP7_75t_L g4111 ( 
.A(n_3967),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_3803),
.B(n_3563),
.Y(n_4112)
);

NAND2xp5_ASAP7_75t_L g4113 ( 
.A(n_3803),
.B(n_3566),
.Y(n_4113)
);

CKINVDCx20_ASAP7_75t_R g4114 ( 
.A(n_3923),
.Y(n_4114)
);

BUFx2_ASAP7_75t_L g4115 ( 
.A(n_3921),
.Y(n_4115)
);

INVx4_ASAP7_75t_L g4116 ( 
.A(n_4019),
.Y(n_4116)
);

BUFx2_ASAP7_75t_L g4117 ( 
.A(n_3973),
.Y(n_4117)
);

BUFx6f_ASAP7_75t_L g4118 ( 
.A(n_4003),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_3978),
.Y(n_4119)
);

INVx2_ASAP7_75t_L g4120 ( 
.A(n_3985),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_L g4121 ( 
.A(n_3922),
.B(n_3568),
.Y(n_4121)
);

OAI22xp5_ASAP7_75t_L g4122 ( 
.A1(n_3797),
.A2(n_3775),
.B1(n_2833),
.B2(n_2808),
.Y(n_4122)
);

O2A1O1Ixp33_ASAP7_75t_L g4123 ( 
.A1(n_3842),
.A2(n_1070),
.B(n_1076),
.C(n_1073),
.Y(n_4123)
);

A2O1A1Ixp33_ASAP7_75t_L g4124 ( 
.A1(n_3815),
.A2(n_1070),
.B(n_1073),
.C(n_1069),
.Y(n_4124)
);

INVx5_ASAP7_75t_L g4125 ( 
.A(n_4003),
.Y(n_4125)
);

AOI22xp33_ASAP7_75t_L g4126 ( 
.A1(n_3818),
.A2(n_3512),
.B1(n_3517),
.B2(n_3576),
.Y(n_4126)
);

OAI21xp5_ASAP7_75t_L g4127 ( 
.A1(n_3797),
.A2(n_3386),
.B(n_3398),
.Y(n_4127)
);

NAND2x1p5_ASAP7_75t_L g4128 ( 
.A(n_4024),
.B(n_3111),
.Y(n_4128)
);

AOI22x1_ASAP7_75t_L g4129 ( 
.A1(n_3808),
.A2(n_947),
.B1(n_956),
.B2(n_944),
.Y(n_4129)
);

INVx4_ASAP7_75t_L g4130 ( 
.A(n_3993),
.Y(n_4130)
);

BUFx3_ASAP7_75t_L g4131 ( 
.A(n_3952),
.Y(n_4131)
);

NAND2xp5_ASAP7_75t_L g4132 ( 
.A(n_3853),
.B(n_3588),
.Y(n_4132)
);

BUFx2_ASAP7_75t_L g4133 ( 
.A(n_3983),
.Y(n_4133)
);

INVx4_ASAP7_75t_L g4134 ( 
.A(n_4036),
.Y(n_4134)
);

INVx5_ASAP7_75t_L g4135 ( 
.A(n_4031),
.Y(n_4135)
);

INVxp67_ASAP7_75t_SL g4136 ( 
.A(n_3799),
.Y(n_4136)
);

INVx3_ASAP7_75t_L g4137 ( 
.A(n_4031),
.Y(n_4137)
);

BUFx2_ASAP7_75t_L g4138 ( 
.A(n_3962),
.Y(n_4138)
);

BUFx2_ASAP7_75t_L g4139 ( 
.A(n_3884),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_L g4140 ( 
.A(n_3953),
.B(n_3591),
.Y(n_4140)
);

BUFx8_ASAP7_75t_L g4141 ( 
.A(n_3879),
.Y(n_4141)
);

INVx3_ASAP7_75t_L g4142 ( 
.A(n_3908),
.Y(n_4142)
);

AOI21xp5_ASAP7_75t_L g4143 ( 
.A1(n_3802),
.A2(n_3669),
.B(n_3460),
.Y(n_4143)
);

AND2x4_ASAP7_75t_L g4144 ( 
.A(n_3879),
.B(n_3501),
.Y(n_4144)
);

BUFx2_ASAP7_75t_L g4145 ( 
.A(n_3956),
.Y(n_4145)
);

AOI21xp5_ASAP7_75t_L g4146 ( 
.A1(n_3799),
.A2(n_3501),
.B(n_3386),
.Y(n_4146)
);

AOI22xp33_ASAP7_75t_SL g4147 ( 
.A1(n_3873),
.A2(n_3876),
.B1(n_3908),
.B2(n_3950),
.Y(n_4147)
);

AOI21x1_ASAP7_75t_L g4148 ( 
.A1(n_4018),
.A2(n_3325),
.B(n_1221),
.Y(n_4148)
);

INVx4_ASAP7_75t_L g4149 ( 
.A(n_3908),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_3986),
.Y(n_4150)
);

BUFx3_ASAP7_75t_L g4151 ( 
.A(n_3955),
.Y(n_4151)
);

NOR2xp33_ASAP7_75t_L g4152 ( 
.A(n_3819),
.B(n_958),
.Y(n_4152)
);

A2O1A1Ixp33_ASAP7_75t_L g4153 ( 
.A1(n_3816),
.A2(n_1080),
.B(n_1082),
.C(n_1069),
.Y(n_4153)
);

O2A1O1Ixp33_ASAP7_75t_SL g4154 ( 
.A1(n_3858),
.A2(n_1082),
.B(n_1086),
.C(n_1080),
.Y(n_4154)
);

AOI21xp5_ASAP7_75t_L g4155 ( 
.A1(n_3800),
.A2(n_3859),
.B(n_3888),
.Y(n_4155)
);

AOI21xp5_ASAP7_75t_L g4156 ( 
.A1(n_3800),
.A2(n_3894),
.B(n_3982),
.Y(n_4156)
);

INVx4_ASAP7_75t_L g4157 ( 
.A(n_3861),
.Y(n_4157)
);

INVx1_ASAP7_75t_SL g4158 ( 
.A(n_3899),
.Y(n_4158)
);

INVx4_ASAP7_75t_L g4159 ( 
.A(n_3811),
.Y(n_4159)
);

AND2x4_ASAP7_75t_L g4160 ( 
.A(n_3851),
.B(n_3594),
.Y(n_4160)
);

AOI21xp5_ASAP7_75t_L g4161 ( 
.A1(n_3874),
.A2(n_3248),
.B(n_3208),
.Y(n_4161)
);

INVx2_ASAP7_75t_L g4162 ( 
.A(n_4027),
.Y(n_4162)
);

AOI22xp5_ASAP7_75t_L g4163 ( 
.A1(n_3917),
.A2(n_3452),
.B1(n_3471),
.B2(n_3432),
.Y(n_4163)
);

INVx5_ASAP7_75t_L g4164 ( 
.A(n_3905),
.Y(n_4164)
);

BUFx6f_ASAP7_75t_L g4165 ( 
.A(n_3863),
.Y(n_4165)
);

AOI22xp33_ASAP7_75t_L g4166 ( 
.A1(n_3914),
.A2(n_3599),
.B1(n_3629),
.B2(n_3605),
.Y(n_4166)
);

CKINVDCx6p67_ASAP7_75t_R g4167 ( 
.A(n_3916),
.Y(n_4167)
);

OR2x6_ASAP7_75t_L g4168 ( 
.A(n_3959),
.B(n_3348),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_4032),
.Y(n_4169)
);

INVx3_ASAP7_75t_L g4170 ( 
.A(n_3932),
.Y(n_4170)
);

NAND2xp5_ASAP7_75t_L g4171 ( 
.A(n_3846),
.B(n_3635),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_SL g4172 ( 
.A(n_3980),
.B(n_3124),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_4032),
.Y(n_4173)
);

NOR2xp33_ASAP7_75t_L g4174 ( 
.A(n_3942),
.B(n_963),
.Y(n_4174)
);

NOR2xp33_ASAP7_75t_L g4175 ( 
.A(n_3824),
.B(n_965),
.Y(n_4175)
);

BUFx6f_ASAP7_75t_L g4176 ( 
.A(n_3939),
.Y(n_4176)
);

INVx2_ASAP7_75t_L g4177 ( 
.A(n_4037),
.Y(n_4177)
);

BUFx2_ASAP7_75t_L g4178 ( 
.A(n_3926),
.Y(n_4178)
);

AOI22xp5_ASAP7_75t_L g4179 ( 
.A1(n_3918),
.A2(n_3422),
.B1(n_3506),
.B2(n_3348),
.Y(n_4179)
);

OAI22xp5_ASAP7_75t_L g4180 ( 
.A1(n_3920),
.A2(n_2833),
.B1(n_3341),
.B2(n_3781),
.Y(n_4180)
);

OR2x2_ASAP7_75t_SL g4181 ( 
.A(n_3935),
.B(n_3649),
.Y(n_4181)
);

INVx2_ASAP7_75t_L g4182 ( 
.A(n_4021),
.Y(n_4182)
);

INVx2_ASAP7_75t_L g4183 ( 
.A(n_3937),
.Y(n_4183)
);

OR2x2_ASAP7_75t_L g4184 ( 
.A(n_3823),
.B(n_3658),
.Y(n_4184)
);

AOI21xp5_ASAP7_75t_L g4185 ( 
.A1(n_3882),
.A2(n_3248),
.B(n_3208),
.Y(n_4185)
);

AOI22xp33_ASAP7_75t_L g4186 ( 
.A1(n_3914),
.A2(n_3659),
.B1(n_3686),
.B2(n_3671),
.Y(n_4186)
);

BUFx6f_ASAP7_75t_L g4187 ( 
.A(n_4025),
.Y(n_4187)
);

OR2x2_ASAP7_75t_L g4188 ( 
.A(n_3909),
.B(n_3827),
.Y(n_4188)
);

BUFx6f_ASAP7_75t_L g4189 ( 
.A(n_3929),
.Y(n_4189)
);

NOR2xp33_ASAP7_75t_L g4190 ( 
.A(n_3801),
.B(n_969),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_4033),
.Y(n_4191)
);

OR2x6_ASAP7_75t_L g4192 ( 
.A(n_3866),
.B(n_3341),
.Y(n_4192)
);

BUFx6f_ASAP7_75t_L g4193 ( 
.A(n_3930),
.Y(n_4193)
);

OAI22xp5_ASAP7_75t_L g4194 ( 
.A1(n_3840),
.A2(n_1089),
.B1(n_1093),
.B2(n_1086),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_L g4195 ( 
.A(n_3847),
.B(n_3696),
.Y(n_4195)
);

AND2x2_ASAP7_75t_L g4196 ( 
.A(n_3904),
.B(n_1089),
.Y(n_4196)
);

OAI22xp5_ASAP7_75t_SL g4197 ( 
.A1(n_3946),
.A2(n_1096),
.B1(n_1100),
.B2(n_1093),
.Y(n_4197)
);

AO22x1_ASAP7_75t_L g4198 ( 
.A1(n_4020),
.A2(n_3742),
.B1(n_3759),
.B2(n_3705),
.Y(n_4198)
);

AOI21xp5_ASAP7_75t_L g4199 ( 
.A1(n_3832),
.A2(n_3323),
.B(n_3300),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_4033),
.Y(n_4200)
);

OAI22xp5_ASAP7_75t_L g4201 ( 
.A1(n_3919),
.A2(n_1100),
.B1(n_1104),
.B2(n_1096),
.Y(n_4201)
);

AOI21xp5_ASAP7_75t_L g4202 ( 
.A1(n_4030),
.A2(n_3958),
.B(n_3947),
.Y(n_4202)
);

INVx2_ASAP7_75t_SL g4203 ( 
.A(n_3992),
.Y(n_4203)
);

AOI21xp33_ASAP7_75t_L g4204 ( 
.A1(n_3974),
.A2(n_3096),
.B(n_3511),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_3801),
.Y(n_4205)
);

OAI22xp5_ASAP7_75t_L g4206 ( 
.A1(n_3910),
.A2(n_1105),
.B1(n_1107),
.B2(n_1104),
.Y(n_4206)
);

AOI22xp5_ASAP7_75t_L g4207 ( 
.A1(n_3852),
.A2(n_3323),
.B1(n_3300),
.B2(n_974),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_3855),
.B(n_3765),
.Y(n_4208)
);

AND2x2_ASAP7_75t_L g4209 ( 
.A(n_4013),
.B(n_1105),
.Y(n_4209)
);

INVx2_ASAP7_75t_L g4210 ( 
.A(n_3906),
.Y(n_4210)
);

NAND2xp5_ASAP7_75t_L g4211 ( 
.A(n_3924),
.B(n_3844),
.Y(n_4211)
);

AOI21xp5_ASAP7_75t_L g4212 ( 
.A1(n_4030),
.A2(n_3096),
.B(n_3428),
.Y(n_4212)
);

O2A1O1Ixp33_ASAP7_75t_L g4213 ( 
.A1(n_3845),
.A2(n_1124),
.B(n_1127),
.C(n_1107),
.Y(n_4213)
);

OAI22xp5_ASAP7_75t_L g4214 ( 
.A1(n_3913),
.A2(n_1124),
.B1(n_1127),
.B2(n_1122),
.Y(n_4214)
);

CKINVDCx5p33_ASAP7_75t_R g4215 ( 
.A(n_3850),
.Y(n_4215)
);

CKINVDCx5p33_ASAP7_75t_R g4216 ( 
.A(n_3854),
.Y(n_4216)
);

BUFx3_ASAP7_75t_L g4217 ( 
.A(n_3991),
.Y(n_4217)
);

INVx2_ASAP7_75t_L g4218 ( 
.A(n_3999),
.Y(n_4218)
);

NAND2xp5_ASAP7_75t_SL g4219 ( 
.A(n_3984),
.B(n_3124),
.Y(n_4219)
);

INVx1_ASAP7_75t_SL g4220 ( 
.A(n_3864),
.Y(n_4220)
);

AOI222xp33_ASAP7_75t_L g4221 ( 
.A1(n_4029),
.A2(n_1132),
.B1(n_1128),
.B2(n_1129),
.C1(n_1122),
.C2(n_980),
.Y(n_4221)
);

NOR2xp33_ASAP7_75t_L g4222 ( 
.A(n_3972),
.B(n_972),
.Y(n_4222)
);

INVx2_ASAP7_75t_L g4223 ( 
.A(n_4000),
.Y(n_4223)
);

O2A1O1Ixp33_ASAP7_75t_L g4224 ( 
.A1(n_3951),
.A2(n_1132),
.B(n_1128),
.C(n_1129),
.Y(n_4224)
);

INVx6_ASAP7_75t_L g4225 ( 
.A(n_3977),
.Y(n_4225)
);

AOI21xp5_ASAP7_75t_L g4226 ( 
.A1(n_4029),
.A2(n_3502),
.B(n_3138),
.Y(n_4226)
);

INVx4_ASAP7_75t_L g4227 ( 
.A(n_4015),
.Y(n_4227)
);

O2A1O1Ixp33_ASAP7_75t_L g4228 ( 
.A1(n_4014),
.A2(n_1516),
.B(n_1519),
.C(n_1515),
.Y(n_4228)
);

AO32x2_ASAP7_75t_L g4229 ( 
.A1(n_3837),
.A2(n_3111),
.A3(n_3767),
.B1(n_3769),
.B2(n_3766),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_4006),
.Y(n_4230)
);

INVx2_ASAP7_75t_L g4231 ( 
.A(n_3940),
.Y(n_4231)
);

OR2x2_ASAP7_75t_L g4232 ( 
.A(n_3838),
.B(n_3771),
.Y(n_4232)
);

BUFx3_ASAP7_75t_L g4233 ( 
.A(n_3931),
.Y(n_4233)
);

BUFx6f_ASAP7_75t_SL g4234 ( 
.A(n_4008),
.Y(n_4234)
);

INVx2_ASAP7_75t_L g4235 ( 
.A(n_3949),
.Y(n_4235)
);

NOR2xp33_ASAP7_75t_L g4236 ( 
.A(n_3987),
.B(n_978),
.Y(n_4236)
);

O2A1O1Ixp33_ASAP7_75t_SL g4237 ( 
.A1(n_3928),
.A2(n_1530),
.B(n_1531),
.C(n_1521),
.Y(n_4237)
);

AO32x2_ASAP7_75t_L g4238 ( 
.A1(n_4001),
.A2(n_1225),
.A3(n_1227),
.B1(n_1226),
.B2(n_1215),
.Y(n_4238)
);

INVx2_ASAP7_75t_SL g4239 ( 
.A(n_3933),
.Y(n_4239)
);

OAI22xp5_ASAP7_75t_L g4240 ( 
.A1(n_3901),
.A2(n_3513),
.B1(n_2989),
.B2(n_2993),
.Y(n_4240)
);

HB1xp67_ASAP7_75t_L g4241 ( 
.A(n_3945),
.Y(n_4241)
);

AOI21xp5_ASAP7_75t_L g4242 ( 
.A1(n_3867),
.A2(n_3138),
.B(n_3124),
.Y(n_4242)
);

INVx2_ASAP7_75t_L g4243 ( 
.A(n_3971),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_L g4244 ( 
.A(n_4009),
.B(n_4016),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_3944),
.Y(n_4245)
);

O2A1O1Ixp33_ASAP7_75t_L g4246 ( 
.A1(n_3989),
.A2(n_1542),
.B(n_1543),
.C(n_1537),
.Y(n_4246)
);

AOI21xp5_ASAP7_75t_L g4247 ( 
.A1(n_3869),
.A2(n_3138),
.B(n_2989),
.Y(n_4247)
);

NOR2xp33_ASAP7_75t_R g4248 ( 
.A(n_4005),
.B(n_2981),
.Y(n_4248)
);

INVx4_ASAP7_75t_L g4249 ( 
.A(n_3975),
.Y(n_4249)
);

AND2x4_ASAP7_75t_L g4250 ( 
.A(n_3871),
.B(n_3113),
.Y(n_4250)
);

AOI21xp5_ASAP7_75t_L g4251 ( 
.A1(n_3870),
.A2(n_3000),
.B(n_2993),
.Y(n_4251)
);

BUFx12f_ASAP7_75t_L g4252 ( 
.A(n_3938),
.Y(n_4252)
);

A2O1A1Ixp33_ASAP7_75t_SL g4253 ( 
.A1(n_3994),
.A2(n_1228),
.B(n_1230),
.C(n_1229),
.Y(n_4253)
);

AOI21x1_ASAP7_75t_L g4254 ( 
.A1(n_3927),
.A2(n_3969),
.B(n_3872),
.Y(n_4254)
);

OAI22xp5_ASAP7_75t_SL g4255 ( 
.A1(n_3902),
.A2(n_1009),
.B1(n_1041),
.B2(n_995),
.Y(n_4255)
);

AND2x2_ASAP7_75t_L g4256 ( 
.A(n_3990),
.B(n_1232),
.Y(n_4256)
);

HB1xp67_ASAP7_75t_L g4257 ( 
.A(n_3892),
.Y(n_4257)
);

OAI22xp5_ASAP7_75t_L g4258 ( 
.A1(n_3897),
.A2(n_3027),
.B1(n_3030),
.B2(n_3000),
.Y(n_4258)
);

AND2x4_ASAP7_75t_L g4259 ( 
.A(n_3970),
.B(n_3027),
.Y(n_4259)
);

BUFx8_ASAP7_75t_L g4260 ( 
.A(n_3976),
.Y(n_4260)
);

BUFx8_ASAP7_75t_SL g4261 ( 
.A(n_3961),
.Y(n_4261)
);

BUFx12f_ASAP7_75t_L g4262 ( 
.A(n_4017),
.Y(n_4262)
);

AOI21xp5_ASAP7_75t_L g4263 ( 
.A1(n_3886),
.A2(n_3064),
.B(n_3030),
.Y(n_4263)
);

BUFx3_ASAP7_75t_L g4264 ( 
.A(n_3963),
.Y(n_4264)
);

BUFx12f_ASAP7_75t_L g4265 ( 
.A(n_4022),
.Y(n_4265)
);

AOI21xp5_ASAP7_75t_L g4266 ( 
.A1(n_3887),
.A2(n_3113),
.B(n_3064),
.Y(n_4266)
);

BUFx12f_ASAP7_75t_L g4267 ( 
.A(n_3965),
.Y(n_4267)
);

OR2x6_ASAP7_75t_L g4268 ( 
.A(n_3877),
.B(n_3117),
.Y(n_4268)
);

INVx2_ASAP7_75t_L g4269 ( 
.A(n_3998),
.Y(n_4269)
);

AOI22xp33_ASAP7_75t_L g4270 ( 
.A1(n_4010),
.A2(n_3516),
.B1(n_2509),
.B2(n_2526),
.Y(n_4270)
);

INVx2_ASAP7_75t_L g4271 ( 
.A(n_3880),
.Y(n_4271)
);

BUFx6f_ASAP7_75t_L g4272 ( 
.A(n_3968),
.Y(n_4272)
);

NOR2xp33_ASAP7_75t_SL g4273 ( 
.A(n_3883),
.B(n_3117),
.Y(n_4273)
);

BUFx10_ASAP7_75t_L g4274 ( 
.A(n_3941),
.Y(n_4274)
);

INVx2_ASAP7_75t_L g4275 ( 
.A(n_3995),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_4002),
.Y(n_4276)
);

INVx2_ASAP7_75t_L g4277 ( 
.A(n_3895),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_L g4278 ( 
.A(n_4060),
.B(n_4076),
.Y(n_4278)
);

OAI21x1_ASAP7_75t_L g4279 ( 
.A1(n_4083),
.A2(n_4148),
.B(n_4212),
.Y(n_4279)
);

NAND2xp5_ASAP7_75t_L g4280 ( 
.A(n_4065),
.B(n_1234),
.Y(n_4280)
);

BUFx2_ASAP7_75t_SL g4281 ( 
.A(n_4114),
.Y(n_4281)
);

NAND2xp5_ASAP7_75t_SL g4282 ( 
.A(n_4159),
.B(n_3898),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_4205),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_4091),
.Y(n_4284)
);

O2A1O1Ixp33_ASAP7_75t_L g4285 ( 
.A1(n_4056),
.A2(n_1235),
.B(n_1238),
.C(n_1236),
.Y(n_4285)
);

BUFx2_ASAP7_75t_L g4286 ( 
.A(n_4110),
.Y(n_4286)
);

OAI21x1_ASAP7_75t_L g4287 ( 
.A1(n_4155),
.A2(n_3890),
.B(n_3889),
.Y(n_4287)
);

INVx1_ASAP7_75t_L g4288 ( 
.A(n_4092),
.Y(n_4288)
);

NAND2xp5_ASAP7_75t_L g4289 ( 
.A(n_4170),
.B(n_1242),
.Y(n_4289)
);

NAND2xp5_ASAP7_75t_L g4290 ( 
.A(n_4111),
.B(n_1243),
.Y(n_4290)
);

AOI221x1_ASAP7_75t_L g4291 ( 
.A1(n_4051),
.A2(n_1251),
.B1(n_1264),
.B2(n_1261),
.C(n_1259),
.Y(n_4291)
);

AOI21xp5_ASAP7_75t_L g4292 ( 
.A1(n_4156),
.A2(n_4007),
.B(n_4004),
.Y(n_4292)
);

INVx2_ASAP7_75t_L g4293 ( 
.A(n_4057),
.Y(n_4293)
);

AO31x2_ASAP7_75t_L g4294 ( 
.A1(n_4169),
.A2(n_1265),
.A3(n_1273),
.B(n_1272),
.Y(n_4294)
);

A2O1A1Ixp33_ASAP7_75t_L g4295 ( 
.A1(n_4084),
.A2(n_3891),
.B(n_1276),
.C(n_1277),
.Y(n_4295)
);

AOI21xp5_ASAP7_75t_L g4296 ( 
.A1(n_4069),
.A2(n_3900),
.B(n_3979),
.Y(n_4296)
);

NOR2xp33_ASAP7_75t_L g4297 ( 
.A(n_4064),
.B(n_3),
.Y(n_4297)
);

BUFx10_ASAP7_75t_L g4298 ( 
.A(n_4070),
.Y(n_4298)
);

OAI21xp5_ASAP7_75t_L g4299 ( 
.A1(n_4079),
.A2(n_3981),
.B(n_1280),
.Y(n_4299)
);

OAI21x1_ASAP7_75t_L g4300 ( 
.A1(n_4143),
.A2(n_3516),
.B(n_2714),
.Y(n_4300)
);

OAI21x1_ASAP7_75t_L g4301 ( 
.A1(n_4127),
.A2(n_2714),
.B(n_1281),
.Y(n_4301)
);

AND2x4_ASAP7_75t_L g4302 ( 
.A(n_4125),
.B(n_1274),
.Y(n_4302)
);

NOR2xp33_ASAP7_75t_L g4303 ( 
.A(n_4043),
.B(n_4),
.Y(n_4303)
);

NOR2xp33_ASAP7_75t_L g4304 ( 
.A(n_4102),
.B(n_6),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_4041),
.Y(n_4305)
);

NOR2xp67_ASAP7_75t_L g4306 ( 
.A(n_4164),
.B(n_1284),
.Y(n_4306)
);

INVx1_ASAP7_75t_L g4307 ( 
.A(n_4045),
.Y(n_4307)
);

INVx2_ASAP7_75t_L g4308 ( 
.A(n_4057),
.Y(n_4308)
);

OAI21xp5_ASAP7_75t_L g4309 ( 
.A1(n_4061),
.A2(n_1288),
.B(n_1286),
.Y(n_4309)
);

OAI21xp33_ASAP7_75t_L g4310 ( 
.A1(n_4136),
.A2(n_1031),
.B(n_1002),
.Y(n_4310)
);

CKINVDCx11_ASAP7_75t_R g4311 ( 
.A(n_4057),
.Y(n_4311)
);

NOR2xp67_ASAP7_75t_SL g4312 ( 
.A(n_4164),
.B(n_1289),
.Y(n_4312)
);

NOR2xp67_ASAP7_75t_L g4313 ( 
.A(n_4164),
.B(n_1290),
.Y(n_4313)
);

BUFx4f_ASAP7_75t_L g4314 ( 
.A(n_4167),
.Y(n_4314)
);

OAI21xp5_ASAP7_75t_L g4315 ( 
.A1(n_4124),
.A2(n_1293),
.B(n_1292),
.Y(n_4315)
);

BUFx10_ASAP7_75t_L g4316 ( 
.A(n_4099),
.Y(n_4316)
);

INVxp67_ASAP7_75t_SL g4317 ( 
.A(n_4139),
.Y(n_4317)
);

OAI22xp33_ASAP7_75t_L g4318 ( 
.A1(n_4062),
.A2(n_987),
.B1(n_990),
.B2(n_979),
.Y(n_4318)
);

NOR2xp33_ASAP7_75t_L g4319 ( 
.A(n_4087),
.B(n_9),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_4052),
.Y(n_4320)
);

O2A1O1Ixp5_ASAP7_75t_SL g4321 ( 
.A1(n_4105),
.A2(n_4191),
.B(n_4200),
.C(n_4173),
.Y(n_4321)
);

AOI21xp5_ASAP7_75t_L g4322 ( 
.A1(n_4172),
.A2(n_4202),
.B(n_4145),
.Y(n_4322)
);

AOI21xp5_ASAP7_75t_L g4323 ( 
.A1(n_4219),
.A2(n_2554),
.B(n_2542),
.Y(n_4323)
);

O2A1O1Ixp33_ASAP7_75t_L g4324 ( 
.A1(n_4153),
.A2(n_1295),
.B(n_1301),
.C(n_1294),
.Y(n_4324)
);

NOR2xp67_ASAP7_75t_L g4325 ( 
.A(n_4159),
.B(n_1305),
.Y(n_4325)
);

OAI22xp33_ASAP7_75t_L g4326 ( 
.A1(n_4134),
.A2(n_997),
.B1(n_999),
.B2(n_994),
.Y(n_4326)
);

AOI21xp5_ASAP7_75t_L g4327 ( 
.A1(n_4117),
.A2(n_2554),
.B(n_2542),
.Y(n_4327)
);

A2O1A1Ixp33_ASAP7_75t_L g4328 ( 
.A1(n_4078),
.A2(n_1307),
.B(n_1006),
.C(n_1007),
.Y(n_4328)
);

NAND2xp33_ASAP7_75t_L g4329 ( 
.A(n_4088),
.B(n_1001),
.Y(n_4329)
);

AOI21xp5_ASAP7_75t_L g4330 ( 
.A1(n_4237),
.A2(n_2554),
.B(n_2542),
.Y(n_4330)
);

AO31x2_ASAP7_75t_L g4331 ( 
.A1(n_4277),
.A2(n_1266),
.A3(n_1267),
.B(n_1224),
.Y(n_4331)
);

CKINVDCx16_ASAP7_75t_R g4332 ( 
.A(n_4131),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_4074),
.Y(n_4333)
);

BUFx6f_ASAP7_75t_L g4334 ( 
.A(n_4059),
.Y(n_4334)
);

CKINVDCx5p33_ASAP7_75t_R g4335 ( 
.A(n_4081),
.Y(n_4335)
);

OAI21x1_ASAP7_75t_L g4336 ( 
.A1(n_4226),
.A2(n_2714),
.B(n_2482),
.Y(n_4336)
);

O2A1O1Ixp33_ASAP7_75t_L g4337 ( 
.A1(n_4201),
.A2(n_1267),
.B(n_1285),
.C(n_1266),
.Y(n_4337)
);

OAI21x1_ASAP7_75t_L g4338 ( 
.A1(n_4254),
.A2(n_2631),
.B(n_2601),
.Y(n_4338)
);

OAI21xp5_ASAP7_75t_L g4339 ( 
.A1(n_4152),
.A2(n_1010),
.B(n_1008),
.Y(n_4339)
);

AOI21xp5_ASAP7_75t_L g4340 ( 
.A1(n_4133),
.A2(n_2556),
.B(n_2554),
.Y(n_4340)
);

AOI21xp5_ASAP7_75t_L g4341 ( 
.A1(n_4138),
.A2(n_2567),
.B(n_2556),
.Y(n_4341)
);

NOR2xp33_ASAP7_75t_L g4342 ( 
.A(n_4038),
.B(n_9),
.Y(n_4342)
);

AOI21x1_ASAP7_75t_L g4343 ( 
.A1(n_4108),
.A2(n_1303),
.B(n_1285),
.Y(n_4343)
);

OAI21xp5_ASAP7_75t_L g4344 ( 
.A1(n_4067),
.A2(n_1016),
.B(n_1015),
.Y(n_4344)
);

AO21x2_ASAP7_75t_L g4345 ( 
.A1(n_4204),
.A2(n_1321),
.B(n_1303),
.Y(n_4345)
);

INVx3_ASAP7_75t_L g4346 ( 
.A(n_4134),
.Y(n_4346)
);

AO31x2_ASAP7_75t_L g4347 ( 
.A1(n_4075),
.A2(n_1350),
.A3(n_1355),
.B(n_1321),
.Y(n_4347)
);

AO31x2_ASAP7_75t_L g4348 ( 
.A1(n_4244),
.A2(n_1355),
.A3(n_1385),
.B(n_1350),
.Y(n_4348)
);

OAI21x1_ASAP7_75t_L g4349 ( 
.A1(n_4146),
.A2(n_2631),
.B(n_2601),
.Y(n_4349)
);

A2O1A1Ixp33_ASAP7_75t_L g4350 ( 
.A1(n_4190),
.A2(n_1034),
.B(n_1042),
.C(n_1035),
.Y(n_4350)
);

AOI21xp5_ASAP7_75t_L g4351 ( 
.A1(n_4217),
.A2(n_2567),
.B(n_2556),
.Y(n_4351)
);

AOI21xp5_ASAP7_75t_L g4352 ( 
.A1(n_4227),
.A2(n_2567),
.B(n_2556),
.Y(n_4352)
);

AOI221x1_ASAP7_75t_L g4353 ( 
.A1(n_4222),
.A2(n_1409),
.B1(n_1432),
.B2(n_1402),
.C(n_1385),
.Y(n_4353)
);

AO31x2_ASAP7_75t_L g4354 ( 
.A1(n_4182),
.A2(n_1409),
.A3(n_1432),
.B(n_1402),
.Y(n_4354)
);

OAI21xp5_ASAP7_75t_L g4355 ( 
.A1(n_4175),
.A2(n_1048),
.B(n_1024),
.Y(n_4355)
);

NOR2xp33_ASAP7_75t_L g4356 ( 
.A(n_4050),
.B(n_10),
.Y(n_4356)
);

AO31x2_ASAP7_75t_L g4357 ( 
.A1(n_4258),
.A2(n_1434),
.A3(n_1436),
.B(n_1433),
.Y(n_4357)
);

NAND2xp33_ASAP7_75t_SL g4358 ( 
.A(n_4115),
.B(n_1050),
.Y(n_4358)
);

AOI22xp5_ASAP7_75t_L g4359 ( 
.A1(n_4221),
.A2(n_1052),
.B1(n_1055),
.B2(n_1051),
.Y(n_4359)
);

CKINVDCx11_ASAP7_75t_R g4360 ( 
.A(n_4085),
.Y(n_4360)
);

AND2x4_ASAP7_75t_L g4361 ( 
.A(n_4125),
.B(n_1433),
.Y(n_4361)
);

CKINVDCx5p33_ASAP7_75t_R g4362 ( 
.A(n_4081),
.Y(n_4362)
);

O2A1O1Ixp33_ASAP7_75t_SL g4363 ( 
.A1(n_4098),
.A2(n_12),
.B(n_10),
.C(n_11),
.Y(n_4363)
);

AO31x2_ASAP7_75t_L g4364 ( 
.A1(n_4275),
.A2(n_1436),
.A3(n_1448),
.B(n_1434),
.Y(n_4364)
);

AOI21xp5_ASAP7_75t_L g4365 ( 
.A1(n_4227),
.A2(n_2572),
.B(n_2567),
.Y(n_4365)
);

AOI21xp5_ASAP7_75t_L g4366 ( 
.A1(n_4178),
.A2(n_2578),
.B(n_2572),
.Y(n_4366)
);

AO31x2_ASAP7_75t_L g4367 ( 
.A1(n_4218),
.A2(n_1466),
.A3(n_1478),
.B(n_1448),
.Y(n_4367)
);

NOR2x1_ASAP7_75t_R g4368 ( 
.A(n_4116),
.B(n_1061),
.Y(n_4368)
);

O2A1O1Ixp33_ASAP7_75t_L g4369 ( 
.A1(n_4194),
.A2(n_1478),
.B(n_1479),
.C(n_1466),
.Y(n_4369)
);

BUFx6f_ASAP7_75t_L g4370 ( 
.A(n_4059),
.Y(n_4370)
);

O2A1O1Ixp5_ASAP7_75t_L g4371 ( 
.A1(n_4157),
.A2(n_1510),
.B(n_1525),
.C(n_1479),
.Y(n_4371)
);

INVx4_ASAP7_75t_L g4372 ( 
.A(n_4059),
.Y(n_4372)
);

A2O1A1Ixp33_ASAP7_75t_L g4373 ( 
.A1(n_4123),
.A2(n_1057),
.B(n_1059),
.C(n_1056),
.Y(n_4373)
);

BUFx2_ASAP7_75t_SL g4374 ( 
.A(n_4157),
.Y(n_4374)
);

AOI221x1_ASAP7_75t_L g4375 ( 
.A1(n_4211),
.A2(n_1510),
.B1(n_1552),
.B2(n_1525),
.C(n_1490),
.Y(n_4375)
);

NAND2xp5_ASAP7_75t_L g4376 ( 
.A(n_4151),
.B(n_13),
.Y(n_4376)
);

AO21x2_ASAP7_75t_L g4377 ( 
.A1(n_4112),
.A2(n_2528),
.B(n_2507),
.Y(n_4377)
);

AO31x2_ASAP7_75t_L g4378 ( 
.A1(n_4223),
.A2(n_2543),
.A3(n_2549),
.B(n_2528),
.Y(n_4378)
);

NOR2xp33_ASAP7_75t_L g4379 ( 
.A(n_4261),
.B(n_4225),
.Y(n_4379)
);

NAND2xp5_ASAP7_75t_L g4380 ( 
.A(n_4055),
.B(n_13),
.Y(n_4380)
);

A2O1A1Ixp33_ASAP7_75t_L g4381 ( 
.A1(n_4236),
.A2(n_4196),
.B(n_4174),
.C(n_4224),
.Y(n_4381)
);

NAND2xp5_ASAP7_75t_SL g4382 ( 
.A(n_4215),
.B(n_4216),
.Y(n_4382)
);

BUFx3_ASAP7_75t_L g4383 ( 
.A(n_4058),
.Y(n_4383)
);

BUFx12f_ASAP7_75t_L g4384 ( 
.A(n_4181),
.Y(n_4384)
);

AOI21xp5_ASAP7_75t_L g4385 ( 
.A1(n_4199),
.A2(n_2578),
.B(n_2572),
.Y(n_4385)
);

AND2x2_ASAP7_75t_L g4386 ( 
.A(n_4053),
.B(n_14),
.Y(n_4386)
);

A2O1A1Ixp33_ASAP7_75t_L g4387 ( 
.A1(n_4095),
.A2(n_1068),
.B(n_1071),
.C(n_1064),
.Y(n_4387)
);

NOR2x1_ASAP7_75t_R g4388 ( 
.A(n_4116),
.B(n_1087),
.Y(n_4388)
);

A2O1A1Ixp33_ASAP7_75t_L g4389 ( 
.A1(n_4106),
.A2(n_1077),
.B(n_1081),
.C(n_1072),
.Y(n_4389)
);

OAI21x1_ASAP7_75t_L g4390 ( 
.A1(n_4161),
.A2(n_2641),
.B(n_2632),
.Y(n_4390)
);

O2A1O1Ixp33_ASAP7_75t_SL g4391 ( 
.A1(n_4090),
.A2(n_16),
.B(n_14),
.C(n_15),
.Y(n_4391)
);

OAI21x1_ASAP7_75t_L g4392 ( 
.A1(n_4185),
.A2(n_2641),
.B(n_2632),
.Y(n_4392)
);

NAND2x1_ASAP7_75t_L g4393 ( 
.A(n_4097),
.B(n_4088),
.Y(n_4393)
);

BUFx6f_ASAP7_75t_L g4394 ( 
.A(n_4187),
.Y(n_4394)
);

NOR2xp33_ASAP7_75t_L g4395 ( 
.A(n_4225),
.B(n_15),
.Y(n_4395)
);

NAND2xp5_ASAP7_75t_L g4396 ( 
.A(n_4048),
.B(n_16),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4082),
.Y(n_4397)
);

BUFx10_ASAP7_75t_L g4398 ( 
.A(n_4189),
.Y(n_4398)
);

INVx5_ASAP7_75t_L g4399 ( 
.A(n_4088),
.Y(n_4399)
);

AOI21x1_ASAP7_75t_L g4400 ( 
.A1(n_4209),
.A2(n_2549),
.B(n_2543),
.Y(n_4400)
);

O2A1O1Ixp33_ASAP7_75t_L g4401 ( 
.A1(n_4206),
.A2(n_2448),
.B(n_2450),
.C(n_2442),
.Y(n_4401)
);

OAI22xp5_ASAP7_75t_L g4402 ( 
.A1(n_4097),
.A2(n_1088),
.B1(n_1090),
.B2(n_1083),
.Y(n_4402)
);

OA21x2_ASAP7_75t_L g4403 ( 
.A1(n_4230),
.A2(n_1094),
.B(n_1091),
.Y(n_4403)
);

AO31x2_ASAP7_75t_L g4404 ( 
.A1(n_4235),
.A2(n_2563),
.A3(n_2579),
.B(n_2555),
.Y(n_4404)
);

NAND2xp5_ASAP7_75t_L g4405 ( 
.A(n_4101),
.B(n_18),
.Y(n_4405)
);

INVxp67_ASAP7_75t_L g4406 ( 
.A(n_4039),
.Y(n_4406)
);

A2O1A1Ixp33_ASAP7_75t_L g4407 ( 
.A1(n_4100),
.A2(n_1097),
.B(n_1098),
.C(n_1095),
.Y(n_4407)
);

AOI21xp5_ASAP7_75t_L g4408 ( 
.A1(n_4122),
.A2(n_2578),
.B(n_2572),
.Y(n_4408)
);

OAI22xp5_ASAP7_75t_L g4409 ( 
.A1(n_4197),
.A2(n_1103),
.B1(n_1111),
.B2(n_1099),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4120),
.Y(n_4410)
);

AOI21xp5_ASAP7_75t_L g4411 ( 
.A1(n_4198),
.A2(n_2582),
.B(n_2578),
.Y(n_4411)
);

O2A1O1Ixp33_ASAP7_75t_L g4412 ( 
.A1(n_4214),
.A2(n_4154),
.B(n_4071),
.C(n_4213),
.Y(n_4412)
);

OAI21x1_ASAP7_75t_L g4413 ( 
.A1(n_4240),
.A2(n_4242),
.B(n_4180),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_4080),
.Y(n_4414)
);

BUFx3_ASAP7_75t_L g4415 ( 
.A(n_4260),
.Y(n_4415)
);

AO31x2_ASAP7_75t_L g4416 ( 
.A1(n_4243),
.A2(n_2563),
.A3(n_2579),
.B(n_2555),
.Y(n_4416)
);

AOI21xp5_ASAP7_75t_SL g4417 ( 
.A1(n_4234),
.A2(n_1113),
.B(n_1112),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_4046),
.Y(n_4418)
);

AOI21xp5_ASAP7_75t_L g4419 ( 
.A1(n_4158),
.A2(n_4273),
.B(n_4220),
.Y(n_4419)
);

AOI21xp5_ASAP7_75t_L g4420 ( 
.A1(n_4096),
.A2(n_2595),
.B(n_2582),
.Y(n_4420)
);

OAI21x1_ASAP7_75t_L g4421 ( 
.A1(n_4113),
.A2(n_2690),
.B(n_2641),
.Y(n_4421)
);

CKINVDCx20_ASAP7_75t_R g4422 ( 
.A(n_4260),
.Y(n_4422)
);

AO31x2_ASAP7_75t_L g4423 ( 
.A1(n_4210),
.A2(n_2588),
.A3(n_2448),
.B(n_2450),
.Y(n_4423)
);

OAI22xp5_ASAP7_75t_L g4424 ( 
.A1(n_4188),
.A2(n_4179),
.B1(n_4129),
.B2(n_4255),
.Y(n_4424)
);

INVx3_ASAP7_75t_L g4425 ( 
.A(n_4233),
.Y(n_4425)
);

INVx3_ASAP7_75t_SL g4426 ( 
.A(n_4187),
.Y(n_4426)
);

INVx2_ASAP7_75t_L g4427 ( 
.A(n_4183),
.Y(n_4427)
);

OAI22xp5_ASAP7_75t_L g4428 ( 
.A1(n_4147),
.A2(n_1116),
.B1(n_1117),
.B2(n_1114),
.Y(n_4428)
);

OAI21xp5_ASAP7_75t_L g4429 ( 
.A1(n_4228),
.A2(n_1121),
.B(n_1119),
.Y(n_4429)
);

AO31x2_ASAP7_75t_L g4430 ( 
.A1(n_4271),
.A2(n_2588),
.A3(n_2458),
.B(n_2464),
.Y(n_4430)
);

O2A1O1Ixp33_ASAP7_75t_SL g4431 ( 
.A1(n_4073),
.A2(n_22),
.B(n_18),
.C(n_20),
.Y(n_4431)
);

OA21x2_ASAP7_75t_L g4432 ( 
.A1(n_4276),
.A2(n_1126),
.B(n_1125),
.Y(n_4432)
);

OAI21x1_ASAP7_75t_L g4433 ( 
.A1(n_4247),
.A2(n_2700),
.B(n_2690),
.Y(n_4433)
);

OAI21x1_ASAP7_75t_L g4434 ( 
.A1(n_4263),
.A2(n_2700),
.B(n_2690),
.Y(n_4434)
);

AO21x1_ASAP7_75t_L g4435 ( 
.A1(n_4072),
.A2(n_20),
.B(n_22),
.Y(n_4435)
);

NAND2xp5_ASAP7_75t_L g4436 ( 
.A(n_4119),
.B(n_23),
.Y(n_4436)
);

INVx4_ASAP7_75t_L g4437 ( 
.A(n_4265),
.Y(n_4437)
);

AO31x2_ASAP7_75t_L g4438 ( 
.A1(n_4162),
.A2(n_2458),
.A3(n_2464),
.B(n_2442),
.Y(n_4438)
);

OAI21x1_ASAP7_75t_L g4439 ( 
.A1(n_4266),
.A2(n_2706),
.B(n_2700),
.Y(n_4439)
);

OAI21xp5_ASAP7_75t_L g4440 ( 
.A1(n_4241),
.A2(n_1133),
.B(n_1130),
.Y(n_4440)
);

AOI21xp5_ASAP7_75t_L g4441 ( 
.A1(n_4063),
.A2(n_2595),
.B(n_2582),
.Y(n_4441)
);

INVx2_ASAP7_75t_L g4442 ( 
.A(n_4093),
.Y(n_4442)
);

INVx2_ASAP7_75t_SL g4443 ( 
.A(n_4274),
.Y(n_4443)
);

OA21x2_ASAP7_75t_L g4444 ( 
.A1(n_4245),
.A2(n_4208),
.B(n_4121),
.Y(n_4444)
);

AND2x2_ASAP7_75t_L g4445 ( 
.A(n_4086),
.B(n_4130),
.Y(n_4445)
);

OAI21xp5_ASAP7_75t_L g4446 ( 
.A1(n_4246),
.A2(n_1135),
.B(n_1134),
.Y(n_4446)
);

INVx1_ASAP7_75t_L g4447 ( 
.A(n_4068),
.Y(n_4447)
);

OAI22xp5_ASAP7_75t_L g4448 ( 
.A1(n_4207),
.A2(n_2474),
.B1(n_2479),
.B2(n_2469),
.Y(n_4448)
);

INVx1_ASAP7_75t_L g4449 ( 
.A(n_4150),
.Y(n_4449)
);

INVx1_ASAP7_75t_L g4450 ( 
.A(n_4103),
.Y(n_4450)
);

AND2x4_ASAP7_75t_L g4451 ( 
.A(n_4125),
.B(n_1484),
.Y(n_4451)
);

NOR2x1_ASAP7_75t_L g4452 ( 
.A(n_4249),
.B(n_2706),
.Y(n_4452)
);

INVx1_ASAP7_75t_L g4453 ( 
.A(n_4104),
.Y(n_4453)
);

BUFx3_ASAP7_75t_L g4454 ( 
.A(n_4141),
.Y(n_4454)
);

INVx1_ASAP7_75t_SL g4455 ( 
.A(n_4264),
.Y(n_4455)
);

AOI22xp33_ASAP7_75t_L g4456 ( 
.A1(n_4160),
.A2(n_2474),
.B1(n_2479),
.B2(n_2469),
.Y(n_4456)
);

A2O1A1Ixp33_ASAP7_75t_L g4457 ( 
.A1(n_4176),
.A2(n_4163),
.B(n_4047),
.C(n_4160),
.Y(n_4457)
);

AOI211x1_ASAP7_75t_L g4458 ( 
.A1(n_4132),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_4458)
);

NOR2xp33_ASAP7_75t_L g4459 ( 
.A(n_4262),
.B(n_26),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_4107),
.Y(n_4460)
);

BUFx6f_ASAP7_75t_L g4461 ( 
.A(n_4187),
.Y(n_4461)
);

AOI21xp5_ASAP7_75t_L g4462 ( 
.A1(n_4063),
.A2(n_2595),
.B(n_2582),
.Y(n_4462)
);

INVx2_ASAP7_75t_L g4463 ( 
.A(n_4044),
.Y(n_4463)
);

AO31x2_ASAP7_75t_L g4464 ( 
.A1(n_4177),
.A2(n_2485),
.A3(n_2488),
.B(n_2483),
.Y(n_4464)
);

NAND2xp5_ASAP7_75t_SL g4465 ( 
.A(n_4176),
.B(n_2595),
.Y(n_4465)
);

AO31x2_ASAP7_75t_L g4466 ( 
.A1(n_4231),
.A2(n_2485),
.A3(n_2488),
.B(n_2483),
.Y(n_4466)
);

BUFx3_ASAP7_75t_L g4467 ( 
.A(n_4141),
.Y(n_4467)
);

INVx2_ASAP7_75t_L g4468 ( 
.A(n_4044),
.Y(n_4468)
);

O2A1O1Ixp33_ASAP7_75t_SL g4469 ( 
.A1(n_4203),
.A2(n_30),
.B(n_27),
.C(n_29),
.Y(n_4469)
);

INVx1_ASAP7_75t_L g4470 ( 
.A(n_4232),
.Y(n_4470)
);

INVx1_ASAP7_75t_L g4471 ( 
.A(n_4140),
.Y(n_4471)
);

AOI221xp5_ASAP7_75t_SL g4472 ( 
.A1(n_4176),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.C(n_32),
.Y(n_4472)
);

OAI21x1_ASAP7_75t_L g4473 ( 
.A1(n_4269),
.A2(n_2706),
.B(n_2501),
.Y(n_4473)
);

A2O1A1Ixp33_ASAP7_75t_L g4474 ( 
.A1(n_4047),
.A2(n_2501),
.B(n_2684),
.C(n_2671),
.Y(n_4474)
);

NAND2xp5_ASAP7_75t_L g4475 ( 
.A(n_4109),
.B(n_31),
.Y(n_4475)
);

CKINVDCx20_ASAP7_75t_R g4476 ( 
.A(n_4130),
.Y(n_4476)
);

OAI21xp5_ASAP7_75t_SL g4477 ( 
.A1(n_4094),
.A2(n_32),
.B(n_33),
.Y(n_4477)
);

INVx1_ASAP7_75t_SL g4478 ( 
.A(n_4248),
.Y(n_4478)
);

INVx5_ASAP7_75t_L g4479 ( 
.A(n_4252),
.Y(n_4479)
);

AOI21xp5_ASAP7_75t_L g4480 ( 
.A1(n_4251),
.A2(n_2648),
.B(n_2621),
.Y(n_4480)
);

AOI221x1_ASAP7_75t_L g4481 ( 
.A1(n_4171),
.A2(n_1540),
.B1(n_1490),
.B2(n_1304),
.C(n_1344),
.Y(n_4481)
);

NAND2xp5_ASAP7_75t_L g4482 ( 
.A(n_4066),
.B(n_34),
.Y(n_4482)
);

OAI21x1_ASAP7_75t_L g4483 ( 
.A1(n_4195),
.A2(n_2688),
.B(n_2684),
.Y(n_4483)
);

AO32x2_ASAP7_75t_L g4484 ( 
.A1(n_4149),
.A2(n_37),
.A3(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_4484)
);

AO31x2_ASAP7_75t_L g4485 ( 
.A1(n_4149),
.A2(n_2699),
.A3(n_2709),
.B(n_2688),
.Y(n_4485)
);

OA21x2_ASAP7_75t_L g4486 ( 
.A1(n_4166),
.A2(n_2709),
.B(n_2699),
.Y(n_4486)
);

OAI21x1_ASAP7_75t_L g4487 ( 
.A1(n_4128),
.A2(n_2712),
.B(n_2711),
.Y(n_4487)
);

OAI21x1_ASAP7_75t_L g4488 ( 
.A1(n_4270),
.A2(n_2712),
.B(n_2711),
.Y(n_4488)
);

AOI21xp5_ASAP7_75t_L g4489 ( 
.A1(n_4257),
.A2(n_2648),
.B(n_2621),
.Y(n_4489)
);

INVx1_ASAP7_75t_L g4490 ( 
.A(n_4184),
.Y(n_4490)
);

INVx1_ASAP7_75t_SL g4491 ( 
.A(n_4066),
.Y(n_4491)
);

OA21x2_ASAP7_75t_L g4492 ( 
.A1(n_4186),
.A2(n_4144),
.B(n_4126),
.Y(n_4492)
);

AOI21xp5_ASAP7_75t_L g4493 ( 
.A1(n_4168),
.A2(n_2648),
.B(n_2621),
.Y(n_4493)
);

AOI21xp5_ASAP7_75t_L g4494 ( 
.A1(n_4168),
.A2(n_2648),
.B(n_2621),
.Y(n_4494)
);

NAND2xp5_ASAP7_75t_L g4495 ( 
.A(n_4165),
.B(n_4054),
.Y(n_4495)
);

OAI21x1_ASAP7_75t_L g4496 ( 
.A1(n_4256),
.A2(n_4137),
.B(n_4142),
.Y(n_4496)
);

INVx1_ASAP7_75t_L g4497 ( 
.A(n_4229),
.Y(n_4497)
);

NAND3xp33_ASAP7_75t_L g4498 ( 
.A(n_4249),
.B(n_1540),
.C(n_1490),
.Y(n_4498)
);

O2A1O1Ixp33_ASAP7_75t_SL g4499 ( 
.A1(n_4239),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_4499)
);

NAND2xp5_ASAP7_75t_L g4500 ( 
.A(n_4165),
.B(n_38),
.Y(n_4500)
);

NAND2xp5_ASAP7_75t_L g4501 ( 
.A(n_4165),
.B(n_4089),
.Y(n_4501)
);

OAI21xp5_ASAP7_75t_L g4502 ( 
.A1(n_4259),
.A2(n_2715),
.B(n_39),
.Y(n_4502)
);

AND2x2_ASAP7_75t_L g4503 ( 
.A(n_4118),
.B(n_41),
.Y(n_4503)
);

AOI21xp5_ASAP7_75t_L g4504 ( 
.A1(n_4253),
.A2(n_2708),
.B(n_2673),
.Y(n_4504)
);

AOI21xp5_ASAP7_75t_L g4505 ( 
.A1(n_4268),
.A2(n_2708),
.B(n_2673),
.Y(n_4505)
);

INVx1_ASAP7_75t_SL g4506 ( 
.A(n_4267),
.Y(n_4506)
);

AOI31xp67_ASAP7_75t_L g4507 ( 
.A1(n_4250),
.A2(n_2715),
.A3(n_1540),
.B(n_1490),
.Y(n_4507)
);

NAND2xp5_ASAP7_75t_L g4508 ( 
.A(n_4144),
.B(n_4077),
.Y(n_4508)
);

NAND2xp5_ASAP7_75t_L g4509 ( 
.A(n_4077),
.B(n_41),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_4229),
.Y(n_4510)
);

AOI21xp5_ASAP7_75t_L g4511 ( 
.A1(n_4268),
.A2(n_2708),
.B(n_2673),
.Y(n_4511)
);

NAND2xp5_ASAP7_75t_L g4512 ( 
.A(n_4077),
.B(n_42),
.Y(n_4512)
);

AOI21xp5_ASAP7_75t_L g4513 ( 
.A1(n_4192),
.A2(n_2708),
.B(n_2673),
.Y(n_4513)
);

NOR2x1_ASAP7_75t_R g4514 ( 
.A(n_4135),
.B(n_1490),
.Y(n_4514)
);

A2O1A1Ixp33_ASAP7_75t_L g4515 ( 
.A1(n_4094),
.A2(n_1540),
.B(n_46),
.C(n_42),
.Y(n_4515)
);

AOI21x1_ASAP7_75t_SL g4516 ( 
.A1(n_4259),
.A2(n_45),
.B(n_48),
.Y(n_4516)
);

AO31x2_ASAP7_75t_L g4517 ( 
.A1(n_4229),
.A2(n_1540),
.A3(n_50),
.B(n_45),
.Y(n_4517)
);

INVx2_ASAP7_75t_L g4518 ( 
.A(n_4427),
.Y(n_4518)
);

INVx1_ASAP7_75t_L g4519 ( 
.A(n_4283),
.Y(n_4519)
);

AO31x2_ASAP7_75t_L g4520 ( 
.A1(n_4497),
.A2(n_4238),
.A3(n_4135),
.B(n_4040),
.Y(n_4520)
);

OAI21x1_ASAP7_75t_L g4521 ( 
.A1(n_4321),
.A2(n_4238),
.B(n_4274),
.Y(n_4521)
);

OAI21x1_ASAP7_75t_L g4522 ( 
.A1(n_4327),
.A2(n_4238),
.B(n_4040),
.Y(n_4522)
);

OAI21xp5_ASAP7_75t_L g4523 ( 
.A1(n_4381),
.A2(n_4250),
.B(n_4192),
.Y(n_4523)
);

OR2x2_ASAP7_75t_L g4524 ( 
.A(n_4284),
.B(n_4118),
.Y(n_4524)
);

AOI21xp33_ASAP7_75t_L g4525 ( 
.A1(n_4403),
.A2(n_4040),
.B(n_4049),
.Y(n_4525)
);

CKINVDCx20_ASAP7_75t_R g4526 ( 
.A(n_4422),
.Y(n_4526)
);

OAI21x1_ASAP7_75t_L g4527 ( 
.A1(n_4340),
.A2(n_4135),
.B(n_4189),
.Y(n_4527)
);

INVx4_ASAP7_75t_L g4528 ( 
.A(n_4479),
.Y(n_4528)
);

AND2x2_ASAP7_75t_L g4529 ( 
.A(n_4286),
.B(n_4118),
.Y(n_4529)
);

OAI21x1_ASAP7_75t_L g4530 ( 
.A1(n_4341),
.A2(n_4193),
.B(n_4189),
.Y(n_4530)
);

NAND2x1p5_ASAP7_75t_L g4531 ( 
.A(n_4454),
.B(n_4193),
.Y(n_4531)
);

INVx1_ASAP7_75t_L g4532 ( 
.A(n_4418),
.Y(n_4532)
);

INVx5_ASAP7_75t_L g4533 ( 
.A(n_4451),
.Y(n_4533)
);

OA21x2_ASAP7_75t_L g4534 ( 
.A1(n_4510),
.A2(n_4042),
.B(n_4193),
.Y(n_4534)
);

INVx2_ASAP7_75t_SL g4535 ( 
.A(n_4383),
.Y(n_4535)
);

OAI21xp5_ASAP7_75t_L g4536 ( 
.A1(n_4477),
.A2(n_4424),
.B(n_4472),
.Y(n_4536)
);

NAND2xp5_ASAP7_75t_L g4537 ( 
.A(n_4288),
.B(n_4272),
.Y(n_4537)
);

OAI21x1_ASAP7_75t_SL g4538 ( 
.A1(n_4322),
.A2(n_49),
.B(n_50),
.Y(n_4538)
);

AND2x4_ASAP7_75t_L g4539 ( 
.A(n_4317),
.B(n_4042),
.Y(n_4539)
);

INVx2_ASAP7_75t_L g4540 ( 
.A(n_4444),
.Y(n_4540)
);

BUFx10_ASAP7_75t_L g4541 ( 
.A(n_4335),
.Y(n_4541)
);

CKINVDCx5p33_ASAP7_75t_R g4542 ( 
.A(n_4362),
.Y(n_4542)
);

AOI22xp33_ASAP7_75t_L g4543 ( 
.A1(n_4492),
.A2(n_4049),
.B1(n_4272),
.B2(n_1258),
.Y(n_4543)
);

NAND2xp5_ASAP7_75t_L g4544 ( 
.A(n_4278),
.B(n_4272),
.Y(n_4544)
);

AOI22x1_ASAP7_75t_L g4545 ( 
.A1(n_4374),
.A2(n_4049),
.B1(n_54),
.B2(n_51),
.Y(n_4545)
);

AND2x4_ASAP7_75t_L g4546 ( 
.A(n_4445),
.B(n_51),
.Y(n_4546)
);

INVx2_ASAP7_75t_L g4547 ( 
.A(n_4444),
.Y(n_4547)
);

NAND2xp5_ASAP7_75t_L g4548 ( 
.A(n_4406),
.B(n_52),
.Y(n_4548)
);

INVxp33_ASAP7_75t_L g4549 ( 
.A(n_4368),
.Y(n_4549)
);

OA21x2_ASAP7_75t_L g4550 ( 
.A1(n_4457),
.A2(n_52),
.B(n_54),
.Y(n_4550)
);

CKINVDCx5p33_ASAP7_75t_R g4551 ( 
.A(n_4281),
.Y(n_4551)
);

OA21x2_ASAP7_75t_L g4552 ( 
.A1(n_4496),
.A2(n_55),
.B(n_56),
.Y(n_4552)
);

BUFx2_ASAP7_75t_L g4553 ( 
.A(n_4476),
.Y(n_4553)
);

AOI21xp5_ASAP7_75t_L g4554 ( 
.A1(n_4420),
.A2(n_1991),
.B(n_1984),
.Y(n_4554)
);

OAI222xp33_ASAP7_75t_L g4555 ( 
.A1(n_4470),
.A2(n_4332),
.B1(n_4414),
.B2(n_4450),
.C1(n_4410),
.C2(n_4490),
.Y(n_4555)
);

OAI21x1_ASAP7_75t_L g4556 ( 
.A1(n_4489),
.A2(n_58),
.B(n_59),
.Y(n_4556)
);

AND2x4_ASAP7_75t_L g4557 ( 
.A(n_4463),
.B(n_58),
.Y(n_4557)
);

OAI21x1_ASAP7_75t_L g4558 ( 
.A1(n_4366),
.A2(n_59),
.B(n_60),
.Y(n_4558)
);

NAND2xp5_ASAP7_75t_L g4559 ( 
.A(n_4333),
.B(n_60),
.Y(n_4559)
);

INVx1_ASAP7_75t_L g4560 ( 
.A(n_4397),
.Y(n_4560)
);

OA21x2_ASAP7_75t_L g4561 ( 
.A1(n_4279),
.A2(n_61),
.B(n_62),
.Y(n_4561)
);

OAI21x1_ASAP7_75t_L g4562 ( 
.A1(n_4413),
.A2(n_62),
.B(n_63),
.Y(n_4562)
);

INVx1_ASAP7_75t_SL g4563 ( 
.A(n_4455),
.Y(n_4563)
);

AOI21xp5_ASAP7_75t_L g4564 ( 
.A1(n_4282),
.A2(n_1991),
.B(n_1984),
.Y(n_4564)
);

INVx2_ASAP7_75t_SL g4565 ( 
.A(n_4467),
.Y(n_4565)
);

INVx2_ASAP7_75t_L g4566 ( 
.A(n_4442),
.Y(n_4566)
);

OAI21x1_ASAP7_75t_L g4567 ( 
.A1(n_4385),
.A2(n_63),
.B(n_64),
.Y(n_4567)
);

NAND2xp5_ASAP7_75t_L g4568 ( 
.A(n_4447),
.B(n_66),
.Y(n_4568)
);

NAND2xp5_ASAP7_75t_L g4569 ( 
.A(n_4449),
.B(n_67),
.Y(n_4569)
);

OAI22xp33_ASAP7_75t_L g4570 ( 
.A1(n_4384),
.A2(n_1258),
.B1(n_1304),
.B2(n_1149),
.Y(n_4570)
);

O2A1O1Ixp33_ASAP7_75t_L g4571 ( 
.A1(n_4350),
.A2(n_72),
.B(n_68),
.C(n_69),
.Y(n_4571)
);

INVx2_ASAP7_75t_L g4572 ( 
.A(n_4293),
.Y(n_4572)
);

INVx2_ASAP7_75t_L g4573 ( 
.A(n_4308),
.Y(n_4573)
);

OR2x6_ASAP7_75t_SL g4574 ( 
.A(n_4376),
.B(n_68),
.Y(n_4574)
);

OAI22xp33_ASAP7_75t_L g4575 ( 
.A1(n_4502),
.A2(n_1258),
.B1(n_1304),
.B2(n_1149),
.Y(n_4575)
);

INVx2_ASAP7_75t_SL g4576 ( 
.A(n_4316),
.Y(n_4576)
);

OR2x2_ASAP7_75t_L g4577 ( 
.A(n_4307),
.B(n_69),
.Y(n_4577)
);

OAI21x1_ASAP7_75t_L g4578 ( 
.A1(n_4421),
.A2(n_74),
.B(n_76),
.Y(n_4578)
);

OR2x2_ASAP7_75t_L g4579 ( 
.A(n_4320),
.B(n_77),
.Y(n_4579)
);

OA21x2_ASAP7_75t_L g4580 ( 
.A1(n_4419),
.A2(n_78),
.B(n_80),
.Y(n_4580)
);

OA21x2_ASAP7_75t_L g4581 ( 
.A1(n_4287),
.A2(n_81),
.B(n_82),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_4305),
.Y(n_4582)
);

NAND2xp5_ASAP7_75t_L g4583 ( 
.A(n_4471),
.B(n_82),
.Y(n_4583)
);

INVx2_ASAP7_75t_L g4584 ( 
.A(n_4453),
.Y(n_4584)
);

OAI21x1_ASAP7_75t_L g4585 ( 
.A1(n_4351),
.A2(n_84),
.B(n_86),
.Y(n_4585)
);

BUFx12f_ASAP7_75t_L g4586 ( 
.A(n_4298),
.Y(n_4586)
);

OA21x2_ASAP7_75t_L g4587 ( 
.A1(n_4292),
.A2(n_84),
.B(n_88),
.Y(n_4587)
);

A2O1A1Ixp33_ASAP7_75t_L g4588 ( 
.A1(n_4358),
.A2(n_90),
.B(n_88),
.C(n_89),
.Y(n_4588)
);

OA21x2_ASAP7_75t_L g4589 ( 
.A1(n_4290),
.A2(n_89),
.B(n_91),
.Y(n_4589)
);

OAI21xp33_ASAP7_75t_L g4590 ( 
.A1(n_4344),
.A2(n_91),
.B(n_92),
.Y(n_4590)
);

BUFx2_ASAP7_75t_L g4591 ( 
.A(n_4425),
.Y(n_4591)
);

NAND2xp5_ASAP7_75t_L g4592 ( 
.A(n_4460),
.B(n_93),
.Y(n_4592)
);

INVx6_ASAP7_75t_L g4593 ( 
.A(n_4479),
.Y(n_4593)
);

OAI21x1_ASAP7_75t_L g4594 ( 
.A1(n_4352),
.A2(n_94),
.B(n_95),
.Y(n_4594)
);

AO21x2_ASAP7_75t_L g4595 ( 
.A1(n_4377),
.A2(n_94),
.B(n_95),
.Y(n_4595)
);

OAI21x1_ASAP7_75t_L g4596 ( 
.A1(n_4365),
.A2(n_96),
.B(n_97),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_4517),
.Y(n_4597)
);

BUFx6f_ASAP7_75t_L g4598 ( 
.A(n_4302),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_4517),
.Y(n_4599)
);

AO31x2_ASAP7_75t_L g4600 ( 
.A1(n_4435),
.A2(n_100),
.A3(n_97),
.B(n_98),
.Y(n_4600)
);

OAI22xp33_ASAP7_75t_L g4601 ( 
.A1(n_4478),
.A2(n_1258),
.B1(n_1304),
.B2(n_1149),
.Y(n_4601)
);

OA21x2_ASAP7_75t_L g4602 ( 
.A1(n_4495),
.A2(n_100),
.B(n_103),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_4517),
.Y(n_4603)
);

OA21x2_ASAP7_75t_L g4604 ( 
.A1(n_4501),
.A2(n_103),
.B(n_104),
.Y(n_4604)
);

AND2x2_ASAP7_75t_L g4605 ( 
.A(n_4346),
.B(n_105),
.Y(n_4605)
);

AO32x2_ASAP7_75t_L g4606 ( 
.A1(n_4443),
.A2(n_108),
.A3(n_106),
.B1(n_107),
.B2(n_110),
.Y(n_4606)
);

NAND2xp5_ASAP7_75t_L g4607 ( 
.A(n_4475),
.B(n_106),
.Y(n_4607)
);

CKINVDCx20_ASAP7_75t_R g4608 ( 
.A(n_4311),
.Y(n_4608)
);

NAND2x1p5_ASAP7_75t_L g4609 ( 
.A(n_4312),
.B(n_1149),
.Y(n_4609)
);

INVx6_ASAP7_75t_L g4610 ( 
.A(n_4479),
.Y(n_4610)
);

AO21x2_ASAP7_75t_L g4611 ( 
.A1(n_4411),
.A2(n_108),
.B(n_110),
.Y(n_4611)
);

O2A1O1Ixp33_ASAP7_75t_L g4612 ( 
.A1(n_4391),
.A2(n_115),
.B(n_111),
.C(n_112),
.Y(n_4612)
);

AOI22xp33_ASAP7_75t_L g4613 ( 
.A1(n_4492),
.A2(n_1258),
.B1(n_1304),
.B2(n_1149),
.Y(n_4613)
);

O2A1O1Ixp33_ASAP7_75t_SL g4614 ( 
.A1(n_4382),
.A2(n_118),
.B(n_115),
.C(n_116),
.Y(n_4614)
);

AO21x2_ASAP7_75t_L g4615 ( 
.A1(n_4345),
.A2(n_118),
.B(n_120),
.Y(n_4615)
);

INVx1_ASAP7_75t_L g4616 ( 
.A(n_4294),
.Y(n_4616)
);

OA21x2_ASAP7_75t_L g4617 ( 
.A1(n_4481),
.A2(n_120),
.B(n_121),
.Y(n_4617)
);

AO21x2_ASAP7_75t_L g4618 ( 
.A1(n_4441),
.A2(n_4462),
.B(n_4280),
.Y(n_4618)
);

INVx1_ASAP7_75t_SL g4619 ( 
.A(n_4506),
.Y(n_4619)
);

NAND2xp5_ASAP7_75t_L g4620 ( 
.A(n_4405),
.B(n_122),
.Y(n_4620)
);

AOI22xp33_ASAP7_75t_L g4621 ( 
.A1(n_4432),
.A2(n_1393),
.B1(n_1469),
.B2(n_1344),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4294),
.Y(n_4622)
);

NOR2xp33_ASAP7_75t_L g4623 ( 
.A(n_4379),
.B(n_123),
.Y(n_4623)
);

OAI21xp5_ASAP7_75t_L g4624 ( 
.A1(n_4440),
.A2(n_123),
.B(n_124),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_4294),
.Y(n_4625)
);

CKINVDCx5p33_ASAP7_75t_R g4626 ( 
.A(n_4415),
.Y(n_4626)
);

AOI221xp5_ASAP7_75t_L g4627 ( 
.A1(n_4458),
.A2(n_1469),
.B1(n_1393),
.B2(n_1344),
.C(n_128),
.Y(n_4627)
);

INVx1_ASAP7_75t_L g4628 ( 
.A(n_4508),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4430),
.Y(n_4629)
);

OA21x2_ASAP7_75t_L g4630 ( 
.A1(n_4338),
.A2(n_4494),
.B(n_4493),
.Y(n_4630)
);

OAI21xp5_ASAP7_75t_L g4631 ( 
.A1(n_4339),
.A2(n_126),
.B(n_127),
.Y(n_4631)
);

A2O1A1Ixp33_ASAP7_75t_L g4632 ( 
.A1(n_4310),
.A2(n_129),
.B(n_127),
.C(n_128),
.Y(n_4632)
);

NAND2xp5_ASAP7_75t_L g4633 ( 
.A(n_4436),
.B(n_4380),
.Y(n_4633)
);

HB1xp67_ASAP7_75t_L g4634 ( 
.A(n_4485),
.Y(n_4634)
);

AOI221xp5_ASAP7_75t_L g4635 ( 
.A1(n_4428),
.A2(n_1469),
.B1(n_1393),
.B2(n_1344),
.C(n_133),
.Y(n_4635)
);

INVx2_ASAP7_75t_L g4636 ( 
.A(n_4468),
.Y(n_4636)
);

OR2x6_ASAP7_75t_L g4637 ( 
.A(n_4393),
.B(n_4306),
.Y(n_4637)
);

OAI21x1_ASAP7_75t_L g4638 ( 
.A1(n_4408),
.A2(n_131),
.B(n_132),
.Y(n_4638)
);

OA21x2_ASAP7_75t_L g4639 ( 
.A1(n_4482),
.A2(n_4500),
.B(n_4483),
.Y(n_4639)
);

INVx2_ASAP7_75t_L g4640 ( 
.A(n_4491),
.Y(n_4640)
);

AND2x2_ASAP7_75t_L g4641 ( 
.A(n_4426),
.B(n_4386),
.Y(n_4641)
);

AO21x2_ASAP7_75t_L g4642 ( 
.A1(n_4309),
.A2(n_132),
.B(n_133),
.Y(n_4642)
);

INVx1_ASAP7_75t_SL g4643 ( 
.A(n_4396),
.Y(n_4643)
);

OR2x2_ASAP7_75t_L g4644 ( 
.A(n_4289),
.B(n_134),
.Y(n_4644)
);

OAI21x1_ASAP7_75t_L g4645 ( 
.A1(n_4513),
.A2(n_4343),
.B(n_4400),
.Y(n_4645)
);

AOI222xp33_ASAP7_75t_L g4646 ( 
.A1(n_4328),
.A2(n_4355),
.B1(n_4318),
.B2(n_4329),
.C1(n_4429),
.C2(n_4389),
.Y(n_4646)
);

INVx1_ASAP7_75t_L g4647 ( 
.A(n_4430),
.Y(n_4647)
);

OA21x2_ASAP7_75t_L g4648 ( 
.A1(n_4509),
.A2(n_134),
.B(n_135),
.Y(n_4648)
);

OR2x6_ASAP7_75t_L g4649 ( 
.A(n_4313),
.B(n_1344),
.Y(n_4649)
);

OAI21x1_ASAP7_75t_L g4650 ( 
.A1(n_4480),
.A2(n_135),
.B(n_136),
.Y(n_4650)
);

NAND2xp5_ASAP7_75t_L g4651 ( 
.A(n_4342),
.B(n_137),
.Y(n_4651)
);

OAI22xp5_ASAP7_75t_L g4652 ( 
.A1(n_4515),
.A2(n_140),
.B1(n_137),
.B2(n_139),
.Y(n_4652)
);

INVx2_ASAP7_75t_L g4653 ( 
.A(n_4485),
.Y(n_4653)
);

OAI21x1_ASAP7_75t_L g4654 ( 
.A1(n_4349),
.A2(n_139),
.B(n_141),
.Y(n_4654)
);

OR2x2_ASAP7_75t_L g4655 ( 
.A(n_4372),
.B(n_142),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_4430),
.Y(n_4656)
);

OAI21xp5_ASAP7_75t_L g4657 ( 
.A1(n_4432),
.A2(n_142),
.B(n_143),
.Y(n_4657)
);

INVx2_ASAP7_75t_L g4658 ( 
.A(n_4485),
.Y(n_4658)
);

OAI21x1_ASAP7_75t_SL g4659 ( 
.A1(n_4437),
.A2(n_4512),
.B(n_4296),
.Y(n_4659)
);

NAND2x1p5_ASAP7_75t_L g4660 ( 
.A(n_4314),
.B(n_1393),
.Y(n_4660)
);

INVx2_ASAP7_75t_L g4661 ( 
.A(n_4347),
.Y(n_4661)
);

INVx2_ASAP7_75t_L g4662 ( 
.A(n_4347),
.Y(n_4662)
);

AOI221xp5_ASAP7_75t_L g4663 ( 
.A1(n_4431),
.A2(n_1469),
.B1(n_1393),
.B2(n_146),
.C(n_144),
.Y(n_4663)
);

OA21x2_ASAP7_75t_L g4664 ( 
.A1(n_4498),
.A2(n_145),
.B(n_150),
.Y(n_4664)
);

OAI21x1_ASAP7_75t_L g4665 ( 
.A1(n_4473),
.A2(n_150),
.B(n_151),
.Y(n_4665)
);

INVx2_ASAP7_75t_L g4666 ( 
.A(n_4394),
.Y(n_4666)
);

OAI21x1_ASAP7_75t_L g4667 ( 
.A1(n_4390),
.A2(n_151),
.B(n_152),
.Y(n_4667)
);

INVx1_ASAP7_75t_L g4668 ( 
.A(n_4423),
.Y(n_4668)
);

OAI21x1_ASAP7_75t_L g4669 ( 
.A1(n_4392),
.A2(n_152),
.B(n_153),
.Y(n_4669)
);

OAI21x1_ASAP7_75t_L g4670 ( 
.A1(n_4516),
.A2(n_154),
.B(n_156),
.Y(n_4670)
);

INVx1_ASAP7_75t_L g4671 ( 
.A(n_4423),
.Y(n_4671)
);

AND2x6_ASAP7_75t_L g4672 ( 
.A(n_4302),
.B(n_1469),
.Y(n_4672)
);

BUFx3_ASAP7_75t_L g4673 ( 
.A(n_4334),
.Y(n_4673)
);

AND2x4_ASAP7_75t_L g4674 ( 
.A(n_4399),
.B(n_157),
.Y(n_4674)
);

OAI21x1_ASAP7_75t_L g4675 ( 
.A1(n_4452),
.A2(n_157),
.B(n_158),
.Y(n_4675)
);

OR2x2_ASAP7_75t_L g4676 ( 
.A(n_4394),
.B(n_158),
.Y(n_4676)
);

OAI21x1_ASAP7_75t_L g4677 ( 
.A1(n_4505),
.A2(n_160),
.B(n_161),
.Y(n_4677)
);

NAND3xp33_ASAP7_75t_L g4678 ( 
.A(n_4403),
.B(n_4395),
.C(n_4499),
.Y(n_4678)
);

INVx3_ASAP7_75t_L g4679 ( 
.A(n_4398),
.Y(n_4679)
);

OAI21x1_ASAP7_75t_L g4680 ( 
.A1(n_4511),
.A2(n_160),
.B(n_162),
.Y(n_4680)
);

BUFx10_ASAP7_75t_L g4681 ( 
.A(n_4356),
.Y(n_4681)
);

BUFx6f_ASAP7_75t_L g4682 ( 
.A(n_4360),
.Y(n_4682)
);

AND2x4_ASAP7_75t_L g4683 ( 
.A(n_4399),
.B(n_162),
.Y(n_4683)
);

OAI21x1_ASAP7_75t_L g4684 ( 
.A1(n_4301),
.A2(n_164),
.B(n_165),
.Y(n_4684)
);

OAI21x1_ASAP7_75t_L g4685 ( 
.A1(n_4300),
.A2(n_164),
.B(n_165),
.Y(n_4685)
);

AND2x4_ASAP7_75t_L g4686 ( 
.A(n_4399),
.B(n_4461),
.Y(n_4686)
);

INVx2_ASAP7_75t_L g4687 ( 
.A(n_4461),
.Y(n_4687)
);

OAI21xp5_ASAP7_75t_L g4688 ( 
.A1(n_4303),
.A2(n_166),
.B(n_167),
.Y(n_4688)
);

OR2x2_ASAP7_75t_L g4689 ( 
.A(n_4334),
.B(n_166),
.Y(n_4689)
);

INVx1_ASAP7_75t_L g4690 ( 
.A(n_4423),
.Y(n_4690)
);

BUFx6f_ASAP7_75t_L g4691 ( 
.A(n_4370),
.Y(n_4691)
);

AOI22xp5_ASAP7_75t_L g4692 ( 
.A1(n_4469),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.Y(n_4692)
);

BUFx6f_ASAP7_75t_L g4693 ( 
.A(n_4370),
.Y(n_4693)
);

INVx2_ASAP7_75t_L g4694 ( 
.A(n_4466),
.Y(n_4694)
);

OA21x2_ASAP7_75t_L g4695 ( 
.A1(n_4375),
.A2(n_168),
.B(n_169),
.Y(n_4695)
);

CKINVDCx20_ASAP7_75t_R g4696 ( 
.A(n_4297),
.Y(n_4696)
);

AND2x4_ASAP7_75t_L g4697 ( 
.A(n_4503),
.B(n_172),
.Y(n_4697)
);

OAI21x1_ASAP7_75t_L g4698 ( 
.A1(n_4323),
.A2(n_172),
.B(n_173),
.Y(n_4698)
);

OAI22xp5_ASAP7_75t_L g4699 ( 
.A1(n_4325),
.A2(n_4459),
.B1(n_4319),
.B2(n_4407),
.Y(n_4699)
);

HB1xp67_ASAP7_75t_L g4700 ( 
.A(n_4438),
.Y(n_4700)
);

NAND2xp5_ASAP7_75t_L g4701 ( 
.A(n_4304),
.B(n_175),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4348),
.Y(n_4702)
);

OAI21x1_ASAP7_75t_L g4703 ( 
.A1(n_4465),
.A2(n_175),
.B(n_176),
.Y(n_4703)
);

OAI21x1_ASAP7_75t_L g4704 ( 
.A1(n_4371),
.A2(n_180),
.B(n_181),
.Y(n_4704)
);

INVx2_ASAP7_75t_L g4705 ( 
.A(n_4466),
.Y(n_4705)
);

OAI221xp5_ASAP7_75t_L g4706 ( 
.A1(n_4359),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.C(n_183),
.Y(n_4706)
);

AND2x2_ASAP7_75t_L g4707 ( 
.A(n_4529),
.B(n_4484),
.Y(n_4707)
);

A2O1A1Ixp33_ASAP7_75t_L g4708 ( 
.A1(n_4536),
.A2(n_4678),
.B(n_4590),
.C(n_4657),
.Y(n_4708)
);

AO31x2_ASAP7_75t_L g4709 ( 
.A1(n_4540),
.A2(n_4353),
.A3(n_4291),
.B(n_4402),
.Y(n_4709)
);

CKINVDCx5p33_ASAP7_75t_R g4710 ( 
.A(n_4526),
.Y(n_4710)
);

NAND2xp5_ASAP7_75t_L g4711 ( 
.A(n_4532),
.B(n_4438),
.Y(n_4711)
);

OAI22xp5_ASAP7_75t_L g4712 ( 
.A1(n_4692),
.A2(n_4326),
.B1(n_4484),
.B2(n_4417),
.Y(n_4712)
);

CKINVDCx6p67_ASAP7_75t_R g4713 ( 
.A(n_4682),
.Y(n_4713)
);

AOI22xp33_ASAP7_75t_L g4714 ( 
.A1(n_4678),
.A2(n_4590),
.B1(n_4580),
.B2(n_4550),
.Y(n_4714)
);

AOI21xp33_ASAP7_75t_L g4715 ( 
.A1(n_4580),
.A2(n_4388),
.B(n_4285),
.Y(n_4715)
);

INVx3_ASAP7_75t_L g4716 ( 
.A(n_4539),
.Y(n_4716)
);

INVx2_ASAP7_75t_L g4717 ( 
.A(n_4547),
.Y(n_4717)
);

BUFx2_ASAP7_75t_L g4718 ( 
.A(n_4608),
.Y(n_4718)
);

OAI22xp33_ASAP7_75t_L g4719 ( 
.A1(n_4692),
.A2(n_4484),
.B1(n_4299),
.B2(n_4486),
.Y(n_4719)
);

OAI211xp5_ASAP7_75t_SL g4720 ( 
.A1(n_4688),
.A2(n_4373),
.B(n_4387),
.C(n_4363),
.Y(n_4720)
);

INVx4_ASAP7_75t_L g4721 ( 
.A(n_4682),
.Y(n_4721)
);

OAI22xp5_ASAP7_75t_L g4722 ( 
.A1(n_4574),
.A2(n_4412),
.B1(n_4456),
.B2(n_4295),
.Y(n_4722)
);

CKINVDCx11_ASAP7_75t_R g4723 ( 
.A(n_4541),
.Y(n_4723)
);

AOI21xp33_ASAP7_75t_L g4724 ( 
.A1(n_4550),
.A2(n_4361),
.B(n_4451),
.Y(n_4724)
);

INVx4_ASAP7_75t_L g4725 ( 
.A(n_4682),
.Y(n_4725)
);

OR2x6_ASAP7_75t_L g4726 ( 
.A(n_4637),
.B(n_4361),
.Y(n_4726)
);

AOI22xp5_ASAP7_75t_L g4727 ( 
.A1(n_4652),
.A2(n_4409),
.B1(n_4448),
.B2(n_4315),
.Y(n_4727)
);

INVx1_ASAP7_75t_L g4728 ( 
.A(n_4519),
.Y(n_4728)
);

INVx1_ASAP7_75t_L g4729 ( 
.A(n_4519),
.Y(n_4729)
);

INVx3_ASAP7_75t_L g4730 ( 
.A(n_4539),
.Y(n_4730)
);

AOI21xp5_ASAP7_75t_L g4731 ( 
.A1(n_4564),
.A2(n_4514),
.B(n_4330),
.Y(n_4731)
);

INVx2_ASAP7_75t_L g4732 ( 
.A(n_4532),
.Y(n_4732)
);

NAND2x1p5_ASAP7_75t_L g4733 ( 
.A(n_4674),
.B(n_4486),
.Y(n_4733)
);

CKINVDCx20_ASAP7_75t_R g4734 ( 
.A(n_4696),
.Y(n_4734)
);

INVx3_ASAP7_75t_L g4735 ( 
.A(n_4528),
.Y(n_4735)
);

AND2x2_ASAP7_75t_L g4736 ( 
.A(n_4591),
.B(n_4348),
.Y(n_4736)
);

AND2x2_ASAP7_75t_L g4737 ( 
.A(n_4641),
.B(n_4438),
.Y(n_4737)
);

O2A1O1Ixp33_ASAP7_75t_SL g4738 ( 
.A1(n_4701),
.A2(n_4446),
.B(n_4474),
.C(n_184),
.Y(n_4738)
);

AOI22xp33_ASAP7_75t_L g4739 ( 
.A1(n_4663),
.A2(n_4488),
.B1(n_4336),
.B2(n_4433),
.Y(n_4739)
);

OR2x2_ASAP7_75t_L g4740 ( 
.A(n_4524),
.B(n_4464),
.Y(n_4740)
);

NAND2xp5_ASAP7_75t_L g4741 ( 
.A(n_4560),
.B(n_4464),
.Y(n_4741)
);

OAI22xp5_ASAP7_75t_L g4742 ( 
.A1(n_4706),
.A2(n_4504),
.B1(n_4401),
.B2(n_4324),
.Y(n_4742)
);

INVx1_ASAP7_75t_L g4743 ( 
.A(n_4560),
.Y(n_4743)
);

AND2x2_ASAP7_75t_L g4744 ( 
.A(n_4553),
.B(n_4464),
.Y(n_4744)
);

INVx2_ASAP7_75t_L g4745 ( 
.A(n_4584),
.Y(n_4745)
);

INVx1_ASAP7_75t_L g4746 ( 
.A(n_4582),
.Y(n_4746)
);

INVx1_ASAP7_75t_L g4747 ( 
.A(n_4582),
.Y(n_4747)
);

NAND2xp33_ASAP7_75t_L g4748 ( 
.A(n_4626),
.B(n_4434),
.Y(n_4748)
);

BUFx2_ASAP7_75t_L g4749 ( 
.A(n_4528),
.Y(n_4749)
);

NAND2xp5_ASAP7_75t_L g4750 ( 
.A(n_4643),
.B(n_4544),
.Y(n_4750)
);

AND2x2_ASAP7_75t_L g4751 ( 
.A(n_4535),
.B(n_4357),
.Y(n_4751)
);

AOI22xp5_ASAP7_75t_L g4752 ( 
.A1(n_4631),
.A2(n_4624),
.B1(n_4627),
.B2(n_4699),
.Y(n_4752)
);

AOI22xp5_ASAP7_75t_L g4753 ( 
.A1(n_4642),
.A2(n_4487),
.B1(n_4439),
.B2(n_4337),
.Y(n_4753)
);

NOR3xp33_ASAP7_75t_SL g4754 ( 
.A(n_4542),
.B(n_4369),
.C(n_182),
.Y(n_4754)
);

AND2x4_ASAP7_75t_L g4755 ( 
.A(n_4533),
.B(n_4666),
.Y(n_4755)
);

NAND2xp33_ASAP7_75t_SL g4756 ( 
.A(n_4551),
.B(n_183),
.Y(n_4756)
);

AND2x2_ASAP7_75t_L g4757 ( 
.A(n_4563),
.B(n_4357),
.Y(n_4757)
);

NAND2xp5_ASAP7_75t_L g4758 ( 
.A(n_4639),
.B(n_4466),
.Y(n_4758)
);

OAI22xp5_ASAP7_75t_L g4759 ( 
.A1(n_4545),
.A2(n_4507),
.B1(n_186),
.B2(n_184),
.Y(n_4759)
);

NAND2xp5_ASAP7_75t_L g4760 ( 
.A(n_4639),
.B(n_4357),
.Y(n_4760)
);

AND2x4_ASAP7_75t_L g4761 ( 
.A(n_4533),
.B(n_4331),
.Y(n_4761)
);

OAI21x1_ASAP7_75t_L g4762 ( 
.A1(n_4527),
.A2(n_4331),
.B(n_4354),
.Y(n_4762)
);

INVx2_ASAP7_75t_L g4763 ( 
.A(n_4518),
.Y(n_4763)
);

INVx2_ASAP7_75t_L g4764 ( 
.A(n_4572),
.Y(n_4764)
);

CKINVDCx5p33_ASAP7_75t_R g4765 ( 
.A(n_4586),
.Y(n_4765)
);

CKINVDCx5p33_ASAP7_75t_R g4766 ( 
.A(n_4541),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_4628),
.Y(n_4767)
);

AOI21xp5_ASAP7_75t_L g4768 ( 
.A1(n_4612),
.A2(n_4575),
.B(n_4587),
.Y(n_4768)
);

NOR2xp33_ASAP7_75t_L g4769 ( 
.A(n_4576),
.B(n_185),
.Y(n_4769)
);

OAI22xp33_ASAP7_75t_L g4770 ( 
.A1(n_4523),
.A2(n_4367),
.B1(n_4354),
.B2(n_4364),
.Y(n_4770)
);

INVx6_ASAP7_75t_L g4771 ( 
.A(n_4593),
.Y(n_4771)
);

OR2x2_ASAP7_75t_L g4772 ( 
.A(n_4537),
.B(n_4378),
.Y(n_4772)
);

BUFx2_ASAP7_75t_L g4773 ( 
.A(n_4593),
.Y(n_4773)
);

NAND2x1_ASAP7_75t_L g4774 ( 
.A(n_4610),
.B(n_4367),
.Y(n_4774)
);

AND2x2_ASAP7_75t_L g4775 ( 
.A(n_4546),
.B(n_4364),
.Y(n_4775)
);

OR2x2_ASAP7_75t_L g4776 ( 
.A(n_4628),
.B(n_4378),
.Y(n_4776)
);

CKINVDCx5p33_ASAP7_75t_R g4777 ( 
.A(n_4619),
.Y(n_4777)
);

INVx2_ASAP7_75t_SL g4778 ( 
.A(n_4565),
.Y(n_4778)
);

O2A1O1Ixp33_ASAP7_75t_SL g4779 ( 
.A1(n_4623),
.A2(n_4651),
.B(n_4588),
.C(n_4607),
.Y(n_4779)
);

AND2x4_ASAP7_75t_L g4780 ( 
.A(n_4533),
.B(n_4404),
.Y(n_4780)
);

OAI22xp5_ASAP7_75t_L g4781 ( 
.A1(n_4545),
.A2(n_190),
.B1(n_187),
.B2(n_188),
.Y(n_4781)
);

INVx3_ASAP7_75t_SL g4782 ( 
.A(n_4610),
.Y(n_4782)
);

AOI21xp33_ASAP7_75t_L g4783 ( 
.A1(n_4659),
.A2(n_187),
.B(n_190),
.Y(n_4783)
);

AOI222xp33_ASAP7_75t_L g4784 ( 
.A1(n_4632),
.A2(n_4620),
.B1(n_4635),
.B2(n_4633),
.C1(n_4681),
.C2(n_4548),
.Y(n_4784)
);

AOI22xp33_ASAP7_75t_L g4785 ( 
.A1(n_4525),
.A2(n_1984),
.B1(n_2004),
.B2(n_1982),
.Y(n_4785)
);

AOI22xp33_ASAP7_75t_L g4786 ( 
.A1(n_4642),
.A2(n_1984),
.B1(n_2004),
.B2(n_1982),
.Y(n_4786)
);

AND2x2_ASAP7_75t_L g4787 ( 
.A(n_4546),
.B(n_4404),
.Y(n_4787)
);

INVx1_ASAP7_75t_L g4788 ( 
.A(n_4597),
.Y(n_4788)
);

INVx2_ASAP7_75t_SL g4789 ( 
.A(n_4681),
.Y(n_4789)
);

AOI22xp33_ASAP7_75t_L g4790 ( 
.A1(n_4589),
.A2(n_2004),
.B1(n_2035),
.B2(n_1991),
.Y(n_4790)
);

CKINVDCx6p67_ASAP7_75t_R g4791 ( 
.A(n_4674),
.Y(n_4791)
);

NAND2xp33_ASAP7_75t_R g4792 ( 
.A(n_4683),
.B(n_191),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_4597),
.Y(n_4793)
);

BUFx2_ASAP7_75t_L g4794 ( 
.A(n_4679),
.Y(n_4794)
);

NAND2xp5_ASAP7_75t_L g4795 ( 
.A(n_4577),
.B(n_4416),
.Y(n_4795)
);

INVx4_ASAP7_75t_L g4796 ( 
.A(n_4683),
.Y(n_4796)
);

INVx2_ASAP7_75t_L g4797 ( 
.A(n_4573),
.Y(n_4797)
);

OAI221xp5_ASAP7_75t_L g4798 ( 
.A1(n_4646),
.A2(n_4571),
.B1(n_4589),
.B2(n_4587),
.C(n_4648),
.Y(n_4798)
);

AND2x2_ASAP7_75t_L g4799 ( 
.A(n_4640),
.B(n_4416),
.Y(n_4799)
);

NAND3xp33_ASAP7_75t_SL g4800 ( 
.A(n_4655),
.B(n_191),
.C(n_192),
.Y(n_4800)
);

AND2x4_ASAP7_75t_L g4801 ( 
.A(n_4687),
.B(n_192),
.Y(n_4801)
);

NAND2xp5_ASAP7_75t_SL g4802 ( 
.A(n_4598),
.B(n_2004),
.Y(n_4802)
);

AOI21xp5_ASAP7_75t_L g4803 ( 
.A1(n_4554),
.A2(n_2035),
.B(n_193),
.Y(n_4803)
);

AOI22xp33_ASAP7_75t_L g4804 ( 
.A1(n_4648),
.A2(n_4604),
.B1(n_4602),
.B2(n_4543),
.Y(n_4804)
);

BUFx3_ASAP7_75t_L g4805 ( 
.A(n_4697),
.Y(n_4805)
);

INVx8_ASAP7_75t_L g4806 ( 
.A(n_4637),
.Y(n_4806)
);

BUFx3_ASAP7_75t_L g4807 ( 
.A(n_4697),
.Y(n_4807)
);

AO21x2_ASAP7_75t_L g4808 ( 
.A1(n_4702),
.A2(n_193),
.B(n_194),
.Y(n_4808)
);

INVx4_ASAP7_75t_L g4809 ( 
.A(n_4602),
.Y(n_4809)
);

AOI21xp5_ASAP7_75t_L g4810 ( 
.A1(n_4611),
.A2(n_2035),
.B(n_194),
.Y(n_4810)
);

OAI22xp5_ASAP7_75t_L g4811 ( 
.A1(n_4579),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.Y(n_4811)
);

INVx2_ASAP7_75t_L g4812 ( 
.A(n_4566),
.Y(n_4812)
);

INVx2_ASAP7_75t_L g4813 ( 
.A(n_4636),
.Y(n_4813)
);

INVx2_ASAP7_75t_L g4814 ( 
.A(n_4534),
.Y(n_4814)
);

AND2x4_ASAP7_75t_L g4815 ( 
.A(n_4673),
.B(n_198),
.Y(n_4815)
);

INVx1_ASAP7_75t_L g4816 ( 
.A(n_4599),
.Y(n_4816)
);

OAI22xp5_ASAP7_75t_L g4817 ( 
.A1(n_4531),
.A2(n_203),
.B1(n_199),
.B2(n_201),
.Y(n_4817)
);

NAND2xp5_ASAP7_75t_L g4818 ( 
.A(n_4559),
.B(n_203),
.Y(n_4818)
);

INVx1_ASAP7_75t_SL g4819 ( 
.A(n_4604),
.Y(n_4819)
);

AND2x2_ASAP7_75t_L g4820 ( 
.A(n_4679),
.B(n_204),
.Y(n_4820)
);

OAI22xp33_ASAP7_75t_L g4821 ( 
.A1(n_4598),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_4821)
);

BUFx2_ASAP7_75t_L g4822 ( 
.A(n_4691),
.Y(n_4822)
);

AOI22xp33_ASAP7_75t_L g4823 ( 
.A1(n_4621),
.A2(n_2035),
.B1(n_209),
.B2(n_205),
.Y(n_4823)
);

INVx1_ASAP7_75t_L g4824 ( 
.A(n_4599),
.Y(n_4824)
);

INVxp33_ASAP7_75t_L g4825 ( 
.A(n_4598),
.Y(n_4825)
);

OAI22xp5_ASAP7_75t_L g4826 ( 
.A1(n_4581),
.A2(n_210),
.B1(n_208),
.B2(n_209),
.Y(n_4826)
);

INVx2_ASAP7_75t_L g4827 ( 
.A(n_4534),
.Y(n_4827)
);

INVx2_ASAP7_75t_L g4828 ( 
.A(n_4530),
.Y(n_4828)
);

OAI22xp5_ASAP7_75t_L g4829 ( 
.A1(n_4581),
.A2(n_212),
.B1(n_208),
.B2(n_211),
.Y(n_4829)
);

AOI22xp33_ASAP7_75t_SL g4830 ( 
.A1(n_4603),
.A2(n_215),
.B1(n_213),
.B2(n_214),
.Y(n_4830)
);

OAI21x1_ASAP7_75t_L g4831 ( 
.A1(n_4522),
.A2(n_214),
.B(n_216),
.Y(n_4831)
);

INVx1_ASAP7_75t_L g4832 ( 
.A(n_4603),
.Y(n_4832)
);

INVx3_ASAP7_75t_L g4833 ( 
.A(n_4691),
.Y(n_4833)
);

NAND3xp33_ASAP7_75t_L g4834 ( 
.A(n_4568),
.B(n_4592),
.C(n_4583),
.Y(n_4834)
);

INVx2_ASAP7_75t_L g4835 ( 
.A(n_4552),
.Y(n_4835)
);

OAI22xp5_ASAP7_75t_L g4836 ( 
.A1(n_4644),
.A2(n_220),
.B1(n_216),
.B2(n_217),
.Y(n_4836)
);

OAI22xp33_ASAP7_75t_L g4837 ( 
.A1(n_4561),
.A2(n_221),
.B1(n_217),
.B2(n_220),
.Y(n_4837)
);

AO31x2_ASAP7_75t_L g4838 ( 
.A1(n_4616),
.A2(n_224),
.A3(n_222),
.B(n_223),
.Y(n_4838)
);

AOI22xp33_ASAP7_75t_L g4839 ( 
.A1(n_4616),
.A2(n_225),
.B1(n_222),
.B2(n_223),
.Y(n_4839)
);

INVx2_ASAP7_75t_L g4840 ( 
.A(n_4552),
.Y(n_4840)
);

OAI21x1_ASAP7_75t_L g4841 ( 
.A1(n_4521),
.A2(n_225),
.B(n_226),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_4622),
.Y(n_4842)
);

HB1xp67_ASAP7_75t_L g4843 ( 
.A(n_4569),
.Y(n_4843)
);

INVx1_ASAP7_75t_L g4844 ( 
.A(n_4622),
.Y(n_4844)
);

NOR2x1p5_ASAP7_75t_L g4845 ( 
.A(n_4676),
.B(n_227),
.Y(n_4845)
);

INVx3_ASAP7_75t_L g4846 ( 
.A(n_4691),
.Y(n_4846)
);

OAI21x1_ASAP7_75t_L g4847 ( 
.A1(n_4653),
.A2(n_227),
.B(n_228),
.Y(n_4847)
);

BUFx10_ASAP7_75t_L g4848 ( 
.A(n_4672),
.Y(n_4848)
);

AND2x2_ASAP7_75t_L g4849 ( 
.A(n_4686),
.B(n_228),
.Y(n_4849)
);

AO31x2_ASAP7_75t_L g4850 ( 
.A1(n_4625),
.A2(n_231),
.A3(n_229),
.B(n_230),
.Y(n_4850)
);

AOI22xp33_ASAP7_75t_L g4851 ( 
.A1(n_4625),
.A2(n_236),
.B1(n_232),
.B2(n_234),
.Y(n_4851)
);

OAI22xp5_ASAP7_75t_L g4852 ( 
.A1(n_4689),
.A2(n_237),
.B1(n_232),
.B2(n_236),
.Y(n_4852)
);

AND2x4_ASAP7_75t_L g4853 ( 
.A(n_4773),
.B(n_4686),
.Y(n_4853)
);

INVx2_ASAP7_75t_L g4854 ( 
.A(n_4772),
.Y(n_4854)
);

INVx4_ASAP7_75t_SL g4855 ( 
.A(n_4782),
.Y(n_4855)
);

AOI221xp5_ASAP7_75t_L g4856 ( 
.A1(n_4708),
.A2(n_4614),
.B1(n_4555),
.B2(n_4538),
.C(n_4549),
.Y(n_4856)
);

AOI22xp33_ASAP7_75t_SL g4857 ( 
.A1(n_4798),
.A2(n_4809),
.B1(n_4819),
.B2(n_4712),
.Y(n_4857)
);

OA21x2_ASAP7_75t_L g4858 ( 
.A1(n_4814),
.A2(n_4658),
.B(n_4647),
.Y(n_4858)
);

AOI21xp5_ASAP7_75t_L g4859 ( 
.A1(n_4768),
.A2(n_4611),
.B(n_4561),
.Y(n_4859)
);

OAI22xp5_ASAP7_75t_L g4860 ( 
.A1(n_4714),
.A2(n_4557),
.B1(n_4605),
.B2(n_4693),
.Y(n_4860)
);

AOI221xp5_ASAP7_75t_L g4861 ( 
.A1(n_4819),
.A2(n_4809),
.B1(n_4719),
.B2(n_4837),
.C(n_4829),
.Y(n_4861)
);

INVx3_ASAP7_75t_L g4862 ( 
.A(n_4806),
.Y(n_4862)
);

INVx1_ASAP7_75t_L g4863 ( 
.A(n_4728),
.Y(n_4863)
);

OAI22xp5_ASAP7_75t_L g4864 ( 
.A1(n_4752),
.A2(n_4557),
.B1(n_4693),
.B2(n_4613),
.Y(n_4864)
);

OAI22xp5_ASAP7_75t_L g4865 ( 
.A1(n_4752),
.A2(n_4693),
.B1(n_4606),
.B2(n_4664),
.Y(n_4865)
);

NAND2xp5_ASAP7_75t_L g4866 ( 
.A(n_4843),
.B(n_4618),
.Y(n_4866)
);

OR2x2_ASAP7_75t_L g4867 ( 
.A(n_4767),
.B(n_4618),
.Y(n_4867)
);

INVx2_ASAP7_75t_L g4868 ( 
.A(n_4827),
.Y(n_4868)
);

NAND2xp5_ASAP7_75t_L g4869 ( 
.A(n_4744),
.B(n_4600),
.Y(n_4869)
);

INVx1_ASAP7_75t_L g4870 ( 
.A(n_4729),
.Y(n_4870)
);

AND2x2_ASAP7_75t_L g4871 ( 
.A(n_4716),
.B(n_4606),
.Y(n_4871)
);

CKINVDCx5p33_ASAP7_75t_R g4872 ( 
.A(n_4710),
.Y(n_4872)
);

BUFx4f_ASAP7_75t_SL g4873 ( 
.A(n_4734),
.Y(n_4873)
);

INVx2_ASAP7_75t_L g4874 ( 
.A(n_4776),
.Y(n_4874)
);

INVx2_ASAP7_75t_L g4875 ( 
.A(n_4740),
.Y(n_4875)
);

AOI21xp33_ASAP7_75t_L g4876 ( 
.A1(n_4784),
.A2(n_4562),
.B(n_4634),
.Y(n_4876)
);

AOI21xp33_ASAP7_75t_L g4877 ( 
.A1(n_4784),
.A2(n_4664),
.B(n_4595),
.Y(n_4877)
);

OA21x2_ASAP7_75t_L g4878 ( 
.A1(n_4835),
.A2(n_4647),
.B(n_4629),
.Y(n_4878)
);

INVx2_ASAP7_75t_L g4879 ( 
.A(n_4799),
.Y(n_4879)
);

AND2x4_ASAP7_75t_L g4880 ( 
.A(n_4796),
.B(n_4520),
.Y(n_4880)
);

NAND2xp5_ASAP7_75t_L g4881 ( 
.A(n_4707),
.B(n_4600),
.Y(n_4881)
);

AOI21xp5_ASAP7_75t_L g4882 ( 
.A1(n_4748),
.A2(n_4595),
.B(n_4638),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4743),
.Y(n_4883)
);

OAI22xp5_ASAP7_75t_L g4884 ( 
.A1(n_4796),
.A2(n_4606),
.B1(n_4660),
.B2(n_4649),
.Y(n_4884)
);

OAI22xp33_ASAP7_75t_L g4885 ( 
.A1(n_4792),
.A2(n_4649),
.B1(n_4617),
.B2(n_4630),
.Y(n_4885)
);

AOI221xp5_ASAP7_75t_L g4886 ( 
.A1(n_4826),
.A2(n_4702),
.B1(n_4600),
.B2(n_4700),
.C(n_4662),
.Y(n_4886)
);

AOI22xp33_ASAP7_75t_L g4887 ( 
.A1(n_4715),
.A2(n_4615),
.B1(n_4661),
.B2(n_4672),
.Y(n_4887)
);

AOI22xp33_ASAP7_75t_L g4888 ( 
.A1(n_4804),
.A2(n_4615),
.B1(n_4672),
.B2(n_4656),
.Y(n_4888)
);

AOI22xp33_ASAP7_75t_SL g4889 ( 
.A1(n_4840),
.A2(n_4617),
.B1(n_4670),
.B2(n_4672),
.Y(n_4889)
);

HB1xp67_ASAP7_75t_L g4890 ( 
.A(n_4732),
.Y(n_4890)
);

NOR2x1_ASAP7_75t_L g4891 ( 
.A(n_4834),
.B(n_4630),
.Y(n_4891)
);

NAND2xp5_ASAP7_75t_L g4892 ( 
.A(n_4746),
.B(n_4747),
.Y(n_4892)
);

AOI21xp5_ASAP7_75t_L g4893 ( 
.A1(n_4779),
.A2(n_4570),
.B(n_4567),
.Y(n_4893)
);

AOI22xp33_ASAP7_75t_L g4894 ( 
.A1(n_4810),
.A2(n_4656),
.B1(n_4668),
.B2(n_4629),
.Y(n_4894)
);

AOI22xp33_ASAP7_75t_L g4895 ( 
.A1(n_4808),
.A2(n_4671),
.B1(n_4690),
.B2(n_4668),
.Y(n_4895)
);

AOI22xp33_ASAP7_75t_L g4896 ( 
.A1(n_4808),
.A2(n_4690),
.B1(n_4671),
.B2(n_4694),
.Y(n_4896)
);

AOI22xp33_ASAP7_75t_L g4897 ( 
.A1(n_4737),
.A2(n_4705),
.B1(n_4695),
.B2(n_4685),
.Y(n_4897)
);

OAI221xp5_ASAP7_75t_L g4898 ( 
.A1(n_4795),
.A2(n_4695),
.B1(n_4609),
.B2(n_4520),
.C(n_4675),
.Y(n_4898)
);

AOI22xp33_ASAP7_75t_L g4899 ( 
.A1(n_4720),
.A2(n_4717),
.B1(n_4722),
.B2(n_4757),
.Y(n_4899)
);

INVx2_ASAP7_75t_L g4900 ( 
.A(n_4751),
.Y(n_4900)
);

INVx2_ASAP7_75t_L g4901 ( 
.A(n_4828),
.Y(n_4901)
);

BUFx12f_ASAP7_75t_L g4902 ( 
.A(n_4723),
.Y(n_4902)
);

AOI21xp5_ASAP7_75t_L g4903 ( 
.A1(n_4738),
.A2(n_4558),
.B(n_4650),
.Y(n_4903)
);

AND2x2_ASAP7_75t_L g4904 ( 
.A(n_4716),
.B(n_4520),
.Y(n_4904)
);

OAI211xp5_ASAP7_75t_L g4905 ( 
.A1(n_4756),
.A2(n_4703),
.B(n_4698),
.C(n_4585),
.Y(n_4905)
);

OAI22xp33_ASAP7_75t_L g4906 ( 
.A1(n_4726),
.A2(n_4601),
.B1(n_4556),
.B2(n_4596),
.Y(n_4906)
);

AOI221xp5_ASAP7_75t_L g4907 ( 
.A1(n_4836),
.A2(n_239),
.B1(n_237),
.B2(n_238),
.C(n_240),
.Y(n_4907)
);

INVx1_ASAP7_75t_L g4908 ( 
.A(n_4788),
.Y(n_4908)
);

AND2x2_ASAP7_75t_L g4909 ( 
.A(n_4730),
.B(n_4578),
.Y(n_4909)
);

AOI21x1_ASAP7_75t_L g4910 ( 
.A1(n_4749),
.A2(n_4645),
.B(n_4654),
.Y(n_4910)
);

HB1xp67_ASAP7_75t_L g4911 ( 
.A(n_4736),
.Y(n_4911)
);

OAI22xp5_ASAP7_75t_L g4912 ( 
.A1(n_4791),
.A2(n_4777),
.B1(n_4789),
.B2(n_4834),
.Y(n_4912)
);

AOI222xp33_ASAP7_75t_L g4913 ( 
.A1(n_4800),
.A2(n_4677),
.B1(n_4680),
.B2(n_4594),
.C1(n_4684),
.C2(n_4669),
.Y(n_4913)
);

INVxp67_ASAP7_75t_L g4914 ( 
.A(n_4794),
.Y(n_4914)
);

AOI21xp5_ASAP7_75t_L g4915 ( 
.A1(n_4806),
.A2(n_4667),
.B(n_4665),
.Y(n_4915)
);

AOI22xp33_ASAP7_75t_L g4916 ( 
.A1(n_4722),
.A2(n_4704),
.B1(n_244),
.B2(n_240),
.Y(n_4916)
);

OAI22xp33_ASAP7_75t_L g4917 ( 
.A1(n_4726),
.A2(n_246),
.B1(n_241),
.B2(n_245),
.Y(n_4917)
);

OAI221xp5_ASAP7_75t_L g4918 ( 
.A1(n_4783),
.A2(n_249),
.B1(n_246),
.B2(n_247),
.C(n_250),
.Y(n_4918)
);

AO22x2_ASAP7_75t_L g4919 ( 
.A1(n_4793),
.A2(n_4824),
.B1(n_4832),
.B2(n_4816),
.Y(n_4919)
);

AOI21xp5_ASAP7_75t_L g4920 ( 
.A1(n_4806),
.A2(n_247),
.B(n_249),
.Y(n_4920)
);

OAI21x1_ASAP7_75t_L g4921 ( 
.A1(n_4758),
.A2(n_250),
.B(n_251),
.Y(n_4921)
);

OR2x6_ASAP7_75t_L g4922 ( 
.A(n_4726),
.B(n_251),
.Y(n_4922)
);

OR2x2_ASAP7_75t_L g4923 ( 
.A(n_4750),
.B(n_252),
.Y(n_4923)
);

AND2x2_ASAP7_75t_L g4924 ( 
.A(n_4730),
.B(n_252),
.Y(n_4924)
);

AND2x2_ASAP7_75t_L g4925 ( 
.A(n_4822),
.B(n_253),
.Y(n_4925)
);

OAI22xp5_ASAP7_75t_L g4926 ( 
.A1(n_4771),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_4926)
);

AOI21xp5_ASAP7_75t_L g4927 ( 
.A1(n_4731),
.A2(n_255),
.B(n_256),
.Y(n_4927)
);

AOI221xp5_ASAP7_75t_L g4928 ( 
.A1(n_4811),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.C(n_260),
.Y(n_4928)
);

NAND2xp5_ASAP7_75t_L g4929 ( 
.A(n_4787),
.B(n_4775),
.Y(n_4929)
);

AND2x4_ASAP7_75t_L g4930 ( 
.A(n_4735),
.B(n_4805),
.Y(n_4930)
);

AND2x4_ASAP7_75t_L g4931 ( 
.A(n_4735),
.B(n_260),
.Y(n_4931)
);

OR2x6_ASAP7_75t_L g4932 ( 
.A(n_4771),
.B(n_261),
.Y(n_4932)
);

INVx1_ASAP7_75t_L g4933 ( 
.A(n_4842),
.Y(n_4933)
);

INVx1_ASAP7_75t_L g4934 ( 
.A(n_4844),
.Y(n_4934)
);

AOI21xp33_ASAP7_75t_L g4935 ( 
.A1(n_4760),
.A2(n_262),
.B(n_263),
.Y(n_4935)
);

AOI22xp33_ASAP7_75t_L g4936 ( 
.A1(n_4845),
.A2(n_266),
.B1(n_264),
.B2(n_265),
.Y(n_4936)
);

AOI222xp33_ASAP7_75t_L g4937 ( 
.A1(n_4852),
.A2(n_264),
.B1(n_265),
.B2(n_267),
.C1(n_268),
.C2(n_269),
.Y(n_4937)
);

OAI22xp33_ASAP7_75t_L g4938 ( 
.A1(n_4727),
.A2(n_274),
.B1(n_270),
.B2(n_271),
.Y(n_4938)
);

OAI211xp5_ASAP7_75t_L g4939 ( 
.A1(n_4754),
.A2(n_277),
.B(n_270),
.C(n_274),
.Y(n_4939)
);

AOI21xp5_ASAP7_75t_L g4940 ( 
.A1(n_4802),
.A2(n_278),
.B(n_281),
.Y(n_4940)
);

AOI22xp33_ASAP7_75t_L g4941 ( 
.A1(n_4845),
.A2(n_282),
.B1(n_278),
.B2(n_281),
.Y(n_4941)
);

OAI22xp5_ASAP7_75t_L g4942 ( 
.A1(n_4727),
.A2(n_286),
.B1(n_283),
.B2(n_284),
.Y(n_4942)
);

OAI21x1_ASAP7_75t_L g4943 ( 
.A1(n_4711),
.A2(n_283),
.B(n_286),
.Y(n_4943)
);

AOI22xp33_ASAP7_75t_SL g4944 ( 
.A1(n_4781),
.A2(n_289),
.B1(n_287),
.B2(n_288),
.Y(n_4944)
);

NAND2xp5_ASAP7_75t_L g4945 ( 
.A(n_4741),
.B(n_287),
.Y(n_4945)
);

NAND3xp33_ASAP7_75t_L g4946 ( 
.A(n_4830),
.B(n_290),
.C(n_291),
.Y(n_4946)
);

OAI22xp5_ASAP7_75t_L g4947 ( 
.A1(n_4807),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.Y(n_4947)
);

AO221x2_ASAP7_75t_L g4948 ( 
.A1(n_4818),
.A2(n_295),
.B1(n_292),
.B2(n_294),
.C(n_296),
.Y(n_4948)
);

OAI211xp5_ASAP7_75t_SL g4949 ( 
.A1(n_4769),
.A2(n_297),
.B(n_294),
.C(n_296),
.Y(n_4949)
);

AOI222xp33_ASAP7_75t_L g4950 ( 
.A1(n_4839),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.C1(n_301),
.C2(n_302),
.Y(n_4950)
);

AOI222xp33_ASAP7_75t_L g4951 ( 
.A1(n_4851),
.A2(n_298),
.B1(n_301),
.B2(n_305),
.C1(n_306),
.C2(n_308),
.Y(n_4951)
);

AO21x2_ASAP7_75t_L g4952 ( 
.A1(n_4770),
.A2(n_306),
.B(n_309),
.Y(n_4952)
);

AOI221xp5_ASAP7_75t_L g4953 ( 
.A1(n_4821),
.A2(n_312),
.B1(n_310),
.B2(n_311),
.C(n_313),
.Y(n_4953)
);

AOI22xp5_ASAP7_75t_L g4954 ( 
.A1(n_4817),
.A2(n_314),
.B1(n_310),
.B2(n_311),
.Y(n_4954)
);

OAI22xp33_ASAP7_75t_L g4955 ( 
.A1(n_4733),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_4955)
);

NAND2xp5_ASAP7_75t_L g4956 ( 
.A(n_4745),
.B(n_315),
.Y(n_4956)
);

BUFx12f_ASAP7_75t_L g4957 ( 
.A(n_4765),
.Y(n_4957)
);

INVx2_ASAP7_75t_L g4958 ( 
.A(n_4764),
.Y(n_4958)
);

INVx2_ASAP7_75t_L g4959 ( 
.A(n_4797),
.Y(n_4959)
);

OAI221xp5_ASAP7_75t_SL g4960 ( 
.A1(n_4739),
.A2(n_4790),
.B1(n_4786),
.B2(n_4803),
.C(n_4849),
.Y(n_4960)
);

INVx1_ASAP7_75t_L g4961 ( 
.A(n_4838),
.Y(n_4961)
);

NAND2x1p5_ASAP7_75t_L g4962 ( 
.A(n_4815),
.B(n_316),
.Y(n_4962)
);

INVx2_ASAP7_75t_L g4963 ( 
.A(n_4763),
.Y(n_4963)
);

AOI21xp5_ASAP7_75t_L g4964 ( 
.A1(n_4759),
.A2(n_317),
.B(n_318),
.Y(n_4964)
);

AOI22xp33_ASAP7_75t_L g4965 ( 
.A1(n_4742),
.A2(n_321),
.B1(n_317),
.B2(n_320),
.Y(n_4965)
);

OAI221xp5_ASAP7_75t_L g4966 ( 
.A1(n_4724),
.A2(n_323),
.B1(n_320),
.B2(n_322),
.C(n_324),
.Y(n_4966)
);

INVx1_ASAP7_75t_SL g4967 ( 
.A(n_4718),
.Y(n_4967)
);

INVx3_ASAP7_75t_L g4968 ( 
.A(n_4721),
.Y(n_4968)
);

INVx1_ASAP7_75t_SL g4969 ( 
.A(n_4713),
.Y(n_4969)
);

BUFx3_ASAP7_75t_L g4970 ( 
.A(n_4721),
.Y(n_4970)
);

AOI22xp33_ASAP7_75t_L g4971 ( 
.A1(n_4785),
.A2(n_325),
.B1(n_322),
.B2(n_324),
.Y(n_4971)
);

OAI21xp5_ASAP7_75t_L g4972 ( 
.A1(n_4841),
.A2(n_325),
.B(n_326),
.Y(n_4972)
);

BUFx2_ASAP7_75t_L g4973 ( 
.A(n_4725),
.Y(n_4973)
);

INVx2_ASAP7_75t_L g4974 ( 
.A(n_4812),
.Y(n_4974)
);

AOI221xp5_ASAP7_75t_L g4975 ( 
.A1(n_4801),
.A2(n_328),
.B1(n_326),
.B2(n_327),
.C(n_329),
.Y(n_4975)
);

INVx2_ASAP7_75t_L g4976 ( 
.A(n_4813),
.Y(n_4976)
);

AND2x2_ASAP7_75t_L g4977 ( 
.A(n_4778),
.B(n_329),
.Y(n_4977)
);

AOI22xp33_ASAP7_75t_SL g4978 ( 
.A1(n_4801),
.A2(n_332),
.B1(n_330),
.B2(n_331),
.Y(n_4978)
);

INVx2_ASAP7_75t_L g4979 ( 
.A(n_4831),
.Y(n_4979)
);

INVx4_ASAP7_75t_L g4980 ( 
.A(n_4725),
.Y(n_4980)
);

OAI21xp33_ASAP7_75t_L g4981 ( 
.A1(n_4820),
.A2(n_330),
.B(n_331),
.Y(n_4981)
);

AO21x2_ASAP7_75t_L g4982 ( 
.A1(n_4762),
.A2(n_332),
.B(n_333),
.Y(n_4982)
);

OAI21x1_ASAP7_75t_L g4983 ( 
.A1(n_4774),
.A2(n_334),
.B(n_335),
.Y(n_4983)
);

AOI22xp33_ASAP7_75t_L g4984 ( 
.A1(n_4823),
.A2(n_337),
.B1(n_335),
.B2(n_336),
.Y(n_4984)
);

INVx1_ASAP7_75t_L g4985 ( 
.A(n_4838),
.Y(n_4985)
);

AO31x2_ASAP7_75t_L g4986 ( 
.A1(n_4838),
.A2(n_339),
.A3(n_336),
.B(n_338),
.Y(n_4986)
);

NAND2xp5_ASAP7_75t_L g4987 ( 
.A(n_4850),
.B(n_341),
.Y(n_4987)
);

AOI21xp5_ASAP7_75t_L g4988 ( 
.A1(n_4755),
.A2(n_341),
.B(n_342),
.Y(n_4988)
);

AOI22xp33_ASAP7_75t_L g4989 ( 
.A1(n_4825),
.A2(n_4780),
.B1(n_4761),
.B2(n_4848),
.Y(n_4989)
);

AOI21x1_ASAP7_75t_L g4990 ( 
.A1(n_4761),
.A2(n_345),
.B(n_346),
.Y(n_4990)
);

CKINVDCx8_ASAP7_75t_R g4991 ( 
.A(n_4855),
.Y(n_4991)
);

INVx1_ASAP7_75t_L g4992 ( 
.A(n_4863),
.Y(n_4992)
);

NAND2xp5_ASAP7_75t_L g4993 ( 
.A(n_4859),
.B(n_4945),
.Y(n_4993)
);

INVxp67_ASAP7_75t_L g4994 ( 
.A(n_4973),
.Y(n_4994)
);

NAND2xp33_ASAP7_75t_R g4995 ( 
.A(n_4862),
.B(n_4766),
.Y(n_4995)
);

NOR2xp33_ASAP7_75t_R g4996 ( 
.A(n_4902),
.B(n_4815),
.Y(n_4996)
);

NAND2xp33_ASAP7_75t_R g4997 ( 
.A(n_4862),
.B(n_4755),
.Y(n_4997)
);

BUFx3_ASAP7_75t_L g4998 ( 
.A(n_4873),
.Y(n_4998)
);

AND2x2_ASAP7_75t_L g4999 ( 
.A(n_4853),
.B(n_4930),
.Y(n_4999)
);

OR2x6_ASAP7_75t_L g5000 ( 
.A(n_4932),
.B(n_4847),
.Y(n_5000)
);

NAND2xp5_ASAP7_75t_L g5001 ( 
.A(n_4979),
.B(n_4850),
.Y(n_5001)
);

AND2x4_ASAP7_75t_L g5002 ( 
.A(n_4855),
.B(n_4833),
.Y(n_5002)
);

INVxp67_ASAP7_75t_L g5003 ( 
.A(n_4912),
.Y(n_5003)
);

NOR2xp33_ASAP7_75t_R g5004 ( 
.A(n_4872),
.B(n_4957),
.Y(n_5004)
);

AND2x4_ASAP7_75t_L g5005 ( 
.A(n_4970),
.B(n_4833),
.Y(n_5005)
);

XOR2xp5_ASAP7_75t_L g5006 ( 
.A(n_4857),
.B(n_4753),
.Y(n_5006)
);

INVx1_ASAP7_75t_L g5007 ( 
.A(n_4870),
.Y(n_5007)
);

BUFx10_ASAP7_75t_L g5008 ( 
.A(n_4931),
.Y(n_5008)
);

INVxp67_ASAP7_75t_L g5009 ( 
.A(n_4967),
.Y(n_5009)
);

AND2x4_ASAP7_75t_L g5010 ( 
.A(n_4930),
.B(n_4846),
.Y(n_5010)
);

CKINVDCx8_ASAP7_75t_R g5011 ( 
.A(n_4932),
.Y(n_5011)
);

INVx1_ASAP7_75t_L g5012 ( 
.A(n_4883),
.Y(n_5012)
);

NAND2xp5_ASAP7_75t_L g5013 ( 
.A(n_4865),
.B(n_4850),
.Y(n_5013)
);

NOR2xp33_ASAP7_75t_R g5014 ( 
.A(n_4968),
.B(n_4846),
.Y(n_5014)
);

INVx1_ASAP7_75t_L g5015 ( 
.A(n_4892),
.Y(n_5015)
);

NAND2xp33_ASAP7_75t_R g5016 ( 
.A(n_4932),
.B(n_4780),
.Y(n_5016)
);

AND2x2_ASAP7_75t_L g5017 ( 
.A(n_4853),
.B(n_4848),
.Y(n_5017)
);

AND2x4_ASAP7_75t_L g5018 ( 
.A(n_4968),
.B(n_4753),
.Y(n_5018)
);

NAND2xp33_ASAP7_75t_R g5019 ( 
.A(n_4922),
.B(n_345),
.Y(n_5019)
);

OR2x6_ASAP7_75t_L g5020 ( 
.A(n_4922),
.B(n_4709),
.Y(n_5020)
);

AND2x2_ASAP7_75t_L g5021 ( 
.A(n_4871),
.B(n_4709),
.Y(n_5021)
);

NOR2xp33_ASAP7_75t_L g5022 ( 
.A(n_4969),
.B(n_348),
.Y(n_5022)
);

AND2x2_ASAP7_75t_L g5023 ( 
.A(n_4909),
.B(n_4709),
.Y(n_5023)
);

AND2x2_ASAP7_75t_L g5024 ( 
.A(n_4914),
.B(n_350),
.Y(n_5024)
);

NAND2xp5_ASAP7_75t_L g5025 ( 
.A(n_4861),
.B(n_350),
.Y(n_5025)
);

NAND2x1p5_ASAP7_75t_L g5026 ( 
.A(n_4931),
.B(n_351),
.Y(n_5026)
);

AND2x4_ASAP7_75t_L g5027 ( 
.A(n_4880),
.B(n_352),
.Y(n_5027)
);

INVxp67_ASAP7_75t_L g5028 ( 
.A(n_4881),
.Y(n_5028)
);

BUFx10_ASAP7_75t_L g5029 ( 
.A(n_4922),
.Y(n_5029)
);

INVx1_ASAP7_75t_L g5030 ( 
.A(n_4961),
.Y(n_5030)
);

CKINVDCx5p33_ASAP7_75t_R g5031 ( 
.A(n_4980),
.Y(n_5031)
);

INVx2_ASAP7_75t_L g5032 ( 
.A(n_4919),
.Y(n_5032)
);

BUFx3_ASAP7_75t_L g5033 ( 
.A(n_4962),
.Y(n_5033)
);

NAND2xp33_ASAP7_75t_R g5034 ( 
.A(n_4880),
.B(n_4924),
.Y(n_5034)
);

NAND2xp5_ASAP7_75t_L g5035 ( 
.A(n_4891),
.B(n_353),
.Y(n_5035)
);

NOR2xp33_ASAP7_75t_R g5036 ( 
.A(n_4980),
.B(n_353),
.Y(n_5036)
);

BUFx3_ASAP7_75t_L g5037 ( 
.A(n_4977),
.Y(n_5037)
);

NAND2xp5_ASAP7_75t_SL g5038 ( 
.A(n_4885),
.B(n_354),
.Y(n_5038)
);

NOR2xp33_ASAP7_75t_R g5039 ( 
.A(n_4925),
.B(n_354),
.Y(n_5039)
);

AND2x4_ASAP7_75t_L g5040 ( 
.A(n_4923),
.B(n_355),
.Y(n_5040)
);

BUFx3_ASAP7_75t_L g5041 ( 
.A(n_4948),
.Y(n_5041)
);

NAND2xp33_ASAP7_75t_R g5042 ( 
.A(n_4920),
.B(n_356),
.Y(n_5042)
);

CKINVDCx16_ASAP7_75t_R g5043 ( 
.A(n_4860),
.Y(n_5043)
);

AND2x4_ASAP7_75t_L g5044 ( 
.A(n_4911),
.B(n_357),
.Y(n_5044)
);

NOR2xp33_ASAP7_75t_R g5045 ( 
.A(n_4990),
.B(n_4936),
.Y(n_5045)
);

NOR2xp33_ASAP7_75t_R g5046 ( 
.A(n_4941),
.B(n_357),
.Y(n_5046)
);

NAND2xp33_ASAP7_75t_SL g5047 ( 
.A(n_4884),
.B(n_4899),
.Y(n_5047)
);

NOR2xp33_ASAP7_75t_R g5048 ( 
.A(n_4910),
.B(n_359),
.Y(n_5048)
);

AND2x4_ASAP7_75t_L g5049 ( 
.A(n_4915),
.B(n_359),
.Y(n_5049)
);

NAND2xp33_ASAP7_75t_R g5050 ( 
.A(n_4893),
.B(n_360),
.Y(n_5050)
);

BUFx3_ASAP7_75t_L g5051 ( 
.A(n_4948),
.Y(n_5051)
);

BUFx5_ASAP7_75t_L g5052 ( 
.A(n_4985),
.Y(n_5052)
);

NAND2xp33_ASAP7_75t_R g5053 ( 
.A(n_4987),
.B(n_361),
.Y(n_5053)
);

BUFx10_ASAP7_75t_L g5054 ( 
.A(n_4981),
.Y(n_5054)
);

AND2x2_ASAP7_75t_L g5055 ( 
.A(n_4891),
.B(n_362),
.Y(n_5055)
);

NAND2xp5_ASAP7_75t_L g5056 ( 
.A(n_4943),
.B(n_362),
.Y(n_5056)
);

NAND2xp33_ASAP7_75t_R g5057 ( 
.A(n_4904),
.B(n_363),
.Y(n_5057)
);

INVx1_ASAP7_75t_L g5058 ( 
.A(n_4908),
.Y(n_5058)
);

OR2x6_ASAP7_75t_L g5059 ( 
.A(n_4988),
.B(n_363),
.Y(n_5059)
);

AND2x4_ASAP7_75t_L g5060 ( 
.A(n_4929),
.B(n_365),
.Y(n_5060)
);

NAND2xp5_ASAP7_75t_L g5061 ( 
.A(n_4876),
.B(n_367),
.Y(n_5061)
);

AND2x4_ASAP7_75t_L g5062 ( 
.A(n_4921),
.B(n_369),
.Y(n_5062)
);

CKINVDCx5p33_ASAP7_75t_R g5063 ( 
.A(n_4956),
.Y(n_5063)
);

CKINVDCx5p33_ASAP7_75t_R g5064 ( 
.A(n_4942),
.Y(n_5064)
);

INVx1_ASAP7_75t_L g5065 ( 
.A(n_4933),
.Y(n_5065)
);

NAND2xp33_ASAP7_75t_R g5066 ( 
.A(n_4927),
.B(n_369),
.Y(n_5066)
);

CKINVDCx11_ASAP7_75t_R g5067 ( 
.A(n_4926),
.Y(n_5067)
);

AND2x2_ASAP7_75t_L g5068 ( 
.A(n_4989),
.B(n_371),
.Y(n_5068)
);

AND2x4_ASAP7_75t_L g5069 ( 
.A(n_4890),
.B(n_371),
.Y(n_5069)
);

NAND2xp33_ASAP7_75t_R g5070 ( 
.A(n_4983),
.B(n_372),
.Y(n_5070)
);

AND2x4_ASAP7_75t_L g5071 ( 
.A(n_4900),
.B(n_372),
.Y(n_5071)
);

NAND2xp33_ASAP7_75t_R g5072 ( 
.A(n_4869),
.B(n_375),
.Y(n_5072)
);

AND2x4_ASAP7_75t_L g5073 ( 
.A(n_4934),
.B(n_375),
.Y(n_5073)
);

OR2x2_ASAP7_75t_L g5074 ( 
.A(n_4866),
.B(n_376),
.Y(n_5074)
);

NOR2xp33_ASAP7_75t_R g5075 ( 
.A(n_4965),
.B(n_376),
.Y(n_5075)
);

NAND2xp33_ASAP7_75t_R g5076 ( 
.A(n_4882),
.B(n_4903),
.Y(n_5076)
);

INVxp67_ASAP7_75t_L g5077 ( 
.A(n_4952),
.Y(n_5077)
);

AND2x2_ASAP7_75t_L g5078 ( 
.A(n_4919),
.B(n_377),
.Y(n_5078)
);

XNOR2xp5_ASAP7_75t_L g5079 ( 
.A(n_4856),
.B(n_377),
.Y(n_5079)
);

CKINVDCx8_ASAP7_75t_R g5080 ( 
.A(n_4981),
.Y(n_5080)
);

INVxp67_ASAP7_75t_L g5081 ( 
.A(n_4952),
.Y(n_5081)
);

INVxp67_ASAP7_75t_L g5082 ( 
.A(n_4877),
.Y(n_5082)
);

BUFx3_ASAP7_75t_L g5083 ( 
.A(n_4954),
.Y(n_5083)
);

NOR2xp33_ASAP7_75t_R g5084 ( 
.A(n_4916),
.B(n_378),
.Y(n_5084)
);

CKINVDCx5p33_ASAP7_75t_R g5085 ( 
.A(n_4947),
.Y(n_5085)
);

CKINVDCx5p33_ASAP7_75t_R g5086 ( 
.A(n_4978),
.Y(n_5086)
);

NOR2xp33_ASAP7_75t_R g5087 ( 
.A(n_4939),
.B(n_378),
.Y(n_5087)
);

NAND2xp5_ASAP7_75t_SL g5088 ( 
.A(n_4906),
.B(n_379),
.Y(n_5088)
);

NAND2xp5_ASAP7_75t_L g5089 ( 
.A(n_4886),
.B(n_379),
.Y(n_5089)
);

NAND2xp33_ASAP7_75t_R g5090 ( 
.A(n_4972),
.B(n_381),
.Y(n_5090)
);

INVxp67_ASAP7_75t_L g5091 ( 
.A(n_4905),
.Y(n_5091)
);

NAND2xp5_ASAP7_75t_L g5092 ( 
.A(n_4982),
.B(n_381),
.Y(n_5092)
);

AND2x4_ASAP7_75t_L g5093 ( 
.A(n_4982),
.B(n_382),
.Y(n_5093)
);

BUFx3_ASAP7_75t_L g5094 ( 
.A(n_4954),
.Y(n_5094)
);

NOR2xp33_ASAP7_75t_R g5095 ( 
.A(n_4938),
.B(n_382),
.Y(n_5095)
);

CKINVDCx5p33_ASAP7_75t_R g5096 ( 
.A(n_4864),
.Y(n_5096)
);

AND2x4_ASAP7_75t_L g5097 ( 
.A(n_4879),
.B(n_383),
.Y(n_5097)
);

XNOR2xp5_ASAP7_75t_L g5098 ( 
.A(n_4946),
.B(n_383),
.Y(n_5098)
);

NAND2xp5_ASAP7_75t_L g5099 ( 
.A(n_5055),
.B(n_4897),
.Y(n_5099)
);

AND2x2_ASAP7_75t_L g5100 ( 
.A(n_4999),
.B(n_4867),
.Y(n_5100)
);

NAND2xp33_ASAP7_75t_SL g5101 ( 
.A(n_5048),
.B(n_4887),
.Y(n_5101)
);

INVx1_ASAP7_75t_L g5102 ( 
.A(n_5030),
.Y(n_5102)
);

BUFx3_ASAP7_75t_L g5103 ( 
.A(n_4991),
.Y(n_5103)
);

OR2x2_ASAP7_75t_L g5104 ( 
.A(n_5015),
.B(n_4960),
.Y(n_5104)
);

INVx1_ASAP7_75t_L g5105 ( 
.A(n_4992),
.Y(n_5105)
);

AND2x2_ASAP7_75t_L g5106 ( 
.A(n_5002),
.B(n_4854),
.Y(n_5106)
);

NOR2xp33_ASAP7_75t_L g5107 ( 
.A(n_4998),
.B(n_4949),
.Y(n_5107)
);

AND2x2_ASAP7_75t_L g5108 ( 
.A(n_5018),
.B(n_4889),
.Y(n_5108)
);

AOI22xp33_ASAP7_75t_SL g5109 ( 
.A1(n_5043),
.A2(n_5013),
.B1(n_5091),
.B2(n_5051),
.Y(n_5109)
);

AND2x2_ASAP7_75t_L g5110 ( 
.A(n_4994),
.B(n_4874),
.Y(n_5110)
);

AND2x4_ASAP7_75t_L g5111 ( 
.A(n_5032),
.B(n_4986),
.Y(n_5111)
);

INVx2_ASAP7_75t_L g5112 ( 
.A(n_5054),
.Y(n_5112)
);

NAND2xp5_ASAP7_75t_L g5113 ( 
.A(n_5083),
.B(n_4888),
.Y(n_5113)
);

HB1xp67_ASAP7_75t_L g5114 ( 
.A(n_5009),
.Y(n_5114)
);

AND2x2_ASAP7_75t_L g5115 ( 
.A(n_5010),
.B(n_4868),
.Y(n_5115)
);

INVx2_ASAP7_75t_SL g5116 ( 
.A(n_5008),
.Y(n_5116)
);

INVx1_ASAP7_75t_L g5117 ( 
.A(n_5007),
.Y(n_5117)
);

INVx1_ASAP7_75t_L g5118 ( 
.A(n_5012),
.Y(n_5118)
);

BUFx2_ASAP7_75t_L g5119 ( 
.A(n_4996),
.Y(n_5119)
);

INVx2_ASAP7_75t_L g5120 ( 
.A(n_5078),
.Y(n_5120)
);

INVx2_ASAP7_75t_L g5121 ( 
.A(n_5041),
.Y(n_5121)
);

INVx2_ASAP7_75t_L g5122 ( 
.A(n_5052),
.Y(n_5122)
);

INVx2_ASAP7_75t_L g5123 ( 
.A(n_5052),
.Y(n_5123)
);

AND2x2_ASAP7_75t_L g5124 ( 
.A(n_5017),
.B(n_4875),
.Y(n_5124)
);

AND2x2_ASAP7_75t_L g5125 ( 
.A(n_5003),
.B(n_4901),
.Y(n_5125)
);

NAND2xp5_ASAP7_75t_L g5126 ( 
.A(n_5094),
.B(n_5035),
.Y(n_5126)
);

OR2x2_ASAP7_75t_L g5127 ( 
.A(n_5058),
.B(n_4986),
.Y(n_5127)
);

INVx1_ASAP7_75t_L g5128 ( 
.A(n_5065),
.Y(n_5128)
);

BUFx3_ASAP7_75t_L g5129 ( 
.A(n_5069),
.Y(n_5129)
);

AND2x2_ASAP7_75t_L g5130 ( 
.A(n_5014),
.B(n_4913),
.Y(n_5130)
);

AND2x2_ASAP7_75t_L g5131 ( 
.A(n_5005),
.B(n_4894),
.Y(n_5131)
);

AND2x2_ASAP7_75t_L g5132 ( 
.A(n_5037),
.B(n_4878),
.Y(n_5132)
);

OR2x2_ASAP7_75t_L g5133 ( 
.A(n_5028),
.B(n_4986),
.Y(n_5133)
);

INVx2_ASAP7_75t_L g5134 ( 
.A(n_5052),
.Y(n_5134)
);

INVx2_ASAP7_75t_L g5135 ( 
.A(n_5052),
.Y(n_5135)
);

INVx1_ASAP7_75t_L g5136 ( 
.A(n_5092),
.Y(n_5136)
);

INVxp67_ASAP7_75t_L g5137 ( 
.A(n_5050),
.Y(n_5137)
);

INVx1_ASAP7_75t_L g5138 ( 
.A(n_5089),
.Y(n_5138)
);

INVx2_ASAP7_75t_L g5139 ( 
.A(n_5080),
.Y(n_5139)
);

NAND2xp5_ASAP7_75t_L g5140 ( 
.A(n_4993),
.B(n_5021),
.Y(n_5140)
);

AND2x4_ASAP7_75t_SL g5141 ( 
.A(n_5029),
.B(n_4958),
.Y(n_5141)
);

BUFx3_ASAP7_75t_L g5142 ( 
.A(n_5069),
.Y(n_5142)
);

AOI22xp33_ASAP7_75t_L g5143 ( 
.A1(n_5006),
.A2(n_4964),
.B1(n_4946),
.B2(n_4898),
.Y(n_5143)
);

INVx2_ASAP7_75t_L g5144 ( 
.A(n_5093),
.Y(n_5144)
);

BUFx3_ASAP7_75t_L g5145 ( 
.A(n_5011),
.Y(n_5145)
);

INVx2_ASAP7_75t_L g5146 ( 
.A(n_5077),
.Y(n_5146)
);

AND2x2_ASAP7_75t_L g5147 ( 
.A(n_5027),
.B(n_4878),
.Y(n_5147)
);

AND2x2_ASAP7_75t_L g5148 ( 
.A(n_5027),
.B(n_4959),
.Y(n_5148)
);

AND2x2_ASAP7_75t_L g5149 ( 
.A(n_5044),
.B(n_4963),
.Y(n_5149)
);

OAI221xp5_ASAP7_75t_L g5150 ( 
.A1(n_5081),
.A2(n_5082),
.B1(n_5076),
.B2(n_5047),
.C(n_5072),
.Y(n_5150)
);

CKINVDCx6p67_ASAP7_75t_R g5151 ( 
.A(n_5033),
.Y(n_5151)
);

INVx1_ASAP7_75t_L g5152 ( 
.A(n_5001),
.Y(n_5152)
);

INVx1_ASAP7_75t_L g5153 ( 
.A(n_5025),
.Y(n_5153)
);

INVx1_ASAP7_75t_L g5154 ( 
.A(n_5061),
.Y(n_5154)
);

INVx2_ASAP7_75t_L g5155 ( 
.A(n_5044),
.Y(n_5155)
);

OR2x2_ASAP7_75t_L g5156 ( 
.A(n_5074),
.B(n_5020),
.Y(n_5156)
);

OR2x2_ASAP7_75t_L g5157 ( 
.A(n_5020),
.B(n_4966),
.Y(n_5157)
);

BUFx3_ASAP7_75t_L g5158 ( 
.A(n_5040),
.Y(n_5158)
);

AND2x2_ASAP7_75t_L g5159 ( 
.A(n_5023),
.B(n_4974),
.Y(n_5159)
);

INVx1_ASAP7_75t_L g5160 ( 
.A(n_5056),
.Y(n_5160)
);

NAND2xp5_ASAP7_75t_L g5161 ( 
.A(n_5049),
.B(n_4955),
.Y(n_5161)
);

INVxp67_ASAP7_75t_L g5162 ( 
.A(n_5053),
.Y(n_5162)
);

INVx3_ASAP7_75t_L g5163 ( 
.A(n_5031),
.Y(n_5163)
);

INVx1_ASAP7_75t_SL g5164 ( 
.A(n_5067),
.Y(n_5164)
);

NAND2xp5_ASAP7_75t_L g5165 ( 
.A(n_5060),
.B(n_4935),
.Y(n_5165)
);

INVx1_ASAP7_75t_L g5166 ( 
.A(n_5024),
.Y(n_5166)
);

INVxp67_ASAP7_75t_L g5167 ( 
.A(n_5019),
.Y(n_5167)
);

AND2x2_ASAP7_75t_L g5168 ( 
.A(n_5073),
.B(n_4976),
.Y(n_5168)
);

OAI221xp5_ASAP7_75t_SL g5169 ( 
.A1(n_5079),
.A2(n_4907),
.B1(n_4975),
.B2(n_4928),
.C(n_4953),
.Y(n_5169)
);

INVx1_ASAP7_75t_L g5170 ( 
.A(n_5098),
.Y(n_5170)
);

NAND2xp5_ASAP7_75t_L g5171 ( 
.A(n_5114),
.B(n_5064),
.Y(n_5171)
);

AND2x2_ASAP7_75t_L g5172 ( 
.A(n_5119),
.B(n_5004),
.Y(n_5172)
);

NAND2xp33_ASAP7_75t_SL g5173 ( 
.A(n_5119),
.B(n_5036),
.Y(n_5173)
);

OR2x2_ASAP7_75t_L g5174 ( 
.A(n_5140),
.B(n_5038),
.Y(n_5174)
);

NOR3xp33_ASAP7_75t_L g5175 ( 
.A(n_5150),
.B(n_5088),
.C(n_5022),
.Y(n_5175)
);

NAND2xp5_ASAP7_75t_L g5176 ( 
.A(n_5166),
.B(n_5153),
.Y(n_5176)
);

NAND2xp5_ASAP7_75t_L g5177 ( 
.A(n_5166),
.B(n_5079),
.Y(n_5177)
);

AND2x2_ASAP7_75t_L g5178 ( 
.A(n_5151),
.B(n_5026),
.Y(n_5178)
);

NOR3xp33_ASAP7_75t_L g5179 ( 
.A(n_5109),
.B(n_4918),
.C(n_4944),
.Y(n_5179)
);

OAI21xp5_ASAP7_75t_SL g5180 ( 
.A1(n_5164),
.A2(n_5098),
.B(n_4937),
.Y(n_5180)
);

NAND2xp5_ASAP7_75t_L g5181 ( 
.A(n_5153),
.B(n_5085),
.Y(n_5181)
);

NAND2xp5_ASAP7_75t_L g5182 ( 
.A(n_5138),
.B(n_5045),
.Y(n_5182)
);

AND2x2_ASAP7_75t_L g5183 ( 
.A(n_5151),
.B(n_5068),
.Y(n_5183)
);

NAND3xp33_ASAP7_75t_L g5184 ( 
.A(n_5143),
.B(n_5066),
.C(n_5090),
.Y(n_5184)
);

NAND2xp5_ASAP7_75t_L g5185 ( 
.A(n_5138),
.B(n_5063),
.Y(n_5185)
);

NAND2xp5_ASAP7_75t_L g5186 ( 
.A(n_5125),
.B(n_5062),
.Y(n_5186)
);

OAI221xp5_ASAP7_75t_SL g5187 ( 
.A1(n_5130),
.A2(n_5059),
.B1(n_4917),
.B2(n_5087),
.C(n_4940),
.Y(n_5187)
);

NAND3xp33_ASAP7_75t_L g5188 ( 
.A(n_5104),
.B(n_5042),
.C(n_5057),
.Y(n_5188)
);

OAI221xp5_ASAP7_75t_L g5189 ( 
.A1(n_5101),
.A2(n_5070),
.B1(n_5034),
.B2(n_5016),
.C(n_5086),
.Y(n_5189)
);

AND2x2_ASAP7_75t_L g5190 ( 
.A(n_5164),
.B(n_5039),
.Y(n_5190)
);

NAND3xp33_ASAP7_75t_L g5191 ( 
.A(n_5104),
.B(n_5059),
.C(n_4951),
.Y(n_5191)
);

AND2x2_ASAP7_75t_L g5192 ( 
.A(n_5121),
.B(n_5000),
.Y(n_5192)
);

AND2x2_ASAP7_75t_L g5193 ( 
.A(n_5121),
.B(n_5000),
.Y(n_5193)
);

NAND2xp5_ASAP7_75t_L g5194 ( 
.A(n_5125),
.B(n_5095),
.Y(n_5194)
);

NAND2xp5_ASAP7_75t_L g5195 ( 
.A(n_5160),
.B(n_5071),
.Y(n_5195)
);

NOR3xp33_ASAP7_75t_L g5196 ( 
.A(n_5146),
.B(n_5096),
.C(n_5084),
.Y(n_5196)
);

NAND2xp5_ASAP7_75t_L g5197 ( 
.A(n_5160),
.B(n_5097),
.Y(n_5197)
);

NAND3xp33_ASAP7_75t_L g5198 ( 
.A(n_5169),
.B(n_4950),
.C(n_4984),
.Y(n_5198)
);

AOI22xp33_ASAP7_75t_SL g5199 ( 
.A1(n_5108),
.A2(n_5046),
.B1(n_5075),
.B2(n_4858),
.Y(n_5199)
);

NAND2xp5_ASAP7_75t_L g5200 ( 
.A(n_5126),
.B(n_4895),
.Y(n_5200)
);

NAND3xp33_ASAP7_75t_L g5201 ( 
.A(n_5157),
.B(n_4971),
.C(n_4995),
.Y(n_5201)
);

OAI221xp5_ASAP7_75t_SL g5202 ( 
.A1(n_5130),
.A2(n_4896),
.B1(n_4997),
.B2(n_387),
.C(n_388),
.Y(n_5202)
);

AND2x2_ASAP7_75t_L g5203 ( 
.A(n_5116),
.B(n_4858),
.Y(n_5203)
);

NAND2xp5_ASAP7_75t_L g5204 ( 
.A(n_5136),
.B(n_384),
.Y(n_5204)
);

AND2x2_ASAP7_75t_L g5205 ( 
.A(n_5116),
.B(n_385),
.Y(n_5205)
);

NAND2xp5_ASAP7_75t_L g5206 ( 
.A(n_5136),
.B(n_389),
.Y(n_5206)
);

NAND2xp5_ASAP7_75t_L g5207 ( 
.A(n_5139),
.B(n_389),
.Y(n_5207)
);

AND2x2_ASAP7_75t_L g5208 ( 
.A(n_5100),
.B(n_391),
.Y(n_5208)
);

NAND3xp33_ASAP7_75t_L g5209 ( 
.A(n_5157),
.B(n_391),
.C(n_392),
.Y(n_5209)
);

AOI221xp5_ASAP7_75t_L g5210 ( 
.A1(n_5146),
.A2(n_392),
.B1(n_393),
.B2(n_394),
.C(n_395),
.Y(n_5210)
);

NAND4xp25_ASAP7_75t_L g5211 ( 
.A(n_5103),
.B(n_396),
.C(n_393),
.D(n_394),
.Y(n_5211)
);

NAND3xp33_ASAP7_75t_L g5212 ( 
.A(n_5139),
.B(n_5162),
.C(n_5112),
.Y(n_5212)
);

AOI221xp5_ASAP7_75t_L g5213 ( 
.A1(n_5099),
.A2(n_396),
.B1(n_397),
.B2(n_398),
.C(n_400),
.Y(n_5213)
);

NAND2xp5_ASAP7_75t_L g5214 ( 
.A(n_5155),
.B(n_398),
.Y(n_5214)
);

AOI22xp33_ASAP7_75t_L g5215 ( 
.A1(n_5137),
.A2(n_402),
.B1(n_400),
.B2(n_401),
.Y(n_5215)
);

OAI22xp5_ASAP7_75t_L g5216 ( 
.A1(n_5108),
.A2(n_404),
.B1(n_401),
.B2(n_403),
.Y(n_5216)
);

INVx2_ASAP7_75t_L g5217 ( 
.A(n_5190),
.Y(n_5217)
);

OR2x2_ASAP7_75t_L g5218 ( 
.A(n_5176),
.B(n_5105),
.Y(n_5218)
);

HB1xp67_ASAP7_75t_L g5219 ( 
.A(n_5171),
.Y(n_5219)
);

INVx1_ASAP7_75t_L g5220 ( 
.A(n_5198),
.Y(n_5220)
);

AOI22xp33_ASAP7_75t_SL g5221 ( 
.A1(n_5189),
.A2(n_5132),
.B1(n_5113),
.B2(n_5120),
.Y(n_5221)
);

OR2x2_ASAP7_75t_L g5222 ( 
.A(n_5177),
.B(n_5105),
.Y(n_5222)
);

HB1xp67_ASAP7_75t_L g5223 ( 
.A(n_5208),
.Y(n_5223)
);

INVx1_ASAP7_75t_L g5224 ( 
.A(n_5204),
.Y(n_5224)
);

AND2x4_ASAP7_75t_L g5225 ( 
.A(n_5172),
.B(n_5103),
.Y(n_5225)
);

INVx2_ASAP7_75t_L g5226 ( 
.A(n_5184),
.Y(n_5226)
);

AND2x2_ASAP7_75t_L g5227 ( 
.A(n_5183),
.B(n_5103),
.Y(n_5227)
);

NOR2x1_ASAP7_75t_L g5228 ( 
.A(n_5212),
.B(n_5163),
.Y(n_5228)
);

OR2x2_ASAP7_75t_L g5229 ( 
.A(n_5174),
.B(n_5117),
.Y(n_5229)
);

HB1xp67_ASAP7_75t_L g5230 ( 
.A(n_5205),
.Y(n_5230)
);

AOI33xp33_ASAP7_75t_L g5231 ( 
.A1(n_5199),
.A2(n_5112),
.A3(n_5152),
.B1(n_5154),
.B2(n_5120),
.B3(n_5110),
.Y(n_5231)
);

INVx1_ASAP7_75t_L g5232 ( 
.A(n_5206),
.Y(n_5232)
);

HB1xp67_ASAP7_75t_L g5233 ( 
.A(n_5207),
.Y(n_5233)
);

NAND2xp5_ASAP7_75t_L g5234 ( 
.A(n_5180),
.B(n_5145),
.Y(n_5234)
);

AND2x2_ASAP7_75t_L g5235 ( 
.A(n_5178),
.B(n_5163),
.Y(n_5235)
);

AND2x2_ASAP7_75t_L g5236 ( 
.A(n_5203),
.B(n_5163),
.Y(n_5236)
);

INVx2_ASAP7_75t_L g5237 ( 
.A(n_5188),
.Y(n_5237)
);

HB1xp67_ASAP7_75t_L g5238 ( 
.A(n_5186),
.Y(n_5238)
);

INVx1_ASAP7_75t_L g5239 ( 
.A(n_5191),
.Y(n_5239)
);

NAND2xp5_ASAP7_75t_L g5240 ( 
.A(n_5216),
.B(n_5145),
.Y(n_5240)
);

AND2x2_ASAP7_75t_L g5241 ( 
.A(n_5185),
.B(n_5100),
.Y(n_5241)
);

INVx2_ASAP7_75t_L g5242 ( 
.A(n_5194),
.Y(n_5242)
);

INVx2_ASAP7_75t_L g5243 ( 
.A(n_5209),
.Y(n_5243)
);

AND2x2_ASAP7_75t_L g5244 ( 
.A(n_5181),
.B(n_5110),
.Y(n_5244)
);

INVx3_ASAP7_75t_L g5245 ( 
.A(n_5192),
.Y(n_5245)
);

INVx2_ASAP7_75t_L g5246 ( 
.A(n_5182),
.Y(n_5246)
);

NAND2xp5_ASAP7_75t_L g5247 ( 
.A(n_5179),
.B(n_5155),
.Y(n_5247)
);

INVx4_ASAP7_75t_L g5248 ( 
.A(n_5193),
.Y(n_5248)
);

BUFx2_ASAP7_75t_L g5249 ( 
.A(n_5173),
.Y(n_5249)
);

INVx2_ASAP7_75t_L g5250 ( 
.A(n_5228),
.Y(n_5250)
);

AND2x2_ASAP7_75t_L g5251 ( 
.A(n_5225),
.B(n_5106),
.Y(n_5251)
);

INVx2_ASAP7_75t_L g5252 ( 
.A(n_5228),
.Y(n_5252)
);

AND2x4_ASAP7_75t_L g5253 ( 
.A(n_5225),
.B(n_5129),
.Y(n_5253)
);

HB1xp67_ASAP7_75t_L g5254 ( 
.A(n_5223),
.Y(n_5254)
);

AND2x2_ASAP7_75t_L g5255 ( 
.A(n_5225),
.B(n_5106),
.Y(n_5255)
);

NAND2xp5_ASAP7_75t_L g5256 ( 
.A(n_5230),
.B(n_5179),
.Y(n_5256)
);

HB1xp67_ASAP7_75t_L g5257 ( 
.A(n_5217),
.Y(n_5257)
);

INVx1_ASAP7_75t_L g5258 ( 
.A(n_5237),
.Y(n_5258)
);

INVx1_ASAP7_75t_L g5259 ( 
.A(n_5237),
.Y(n_5259)
);

INVx1_ASAP7_75t_L g5260 ( 
.A(n_5237),
.Y(n_5260)
);

NAND2xp5_ASAP7_75t_SL g5261 ( 
.A(n_5225),
.B(n_5199),
.Y(n_5261)
);

HB1xp67_ASAP7_75t_L g5262 ( 
.A(n_5217),
.Y(n_5262)
);

INVx1_ASAP7_75t_L g5263 ( 
.A(n_5226),
.Y(n_5263)
);

INVxp67_ASAP7_75t_L g5264 ( 
.A(n_5227),
.Y(n_5264)
);

NAND2xp5_ASAP7_75t_L g5265 ( 
.A(n_5233),
.B(n_5129),
.Y(n_5265)
);

INVx3_ASAP7_75t_L g5266 ( 
.A(n_5248),
.Y(n_5266)
);

AND2x2_ASAP7_75t_L g5267 ( 
.A(n_5227),
.B(n_5142),
.Y(n_5267)
);

AND2x2_ASAP7_75t_L g5268 ( 
.A(n_5249),
.B(n_5142),
.Y(n_5268)
);

AND2x4_ASAP7_75t_L g5269 ( 
.A(n_5235),
.B(n_5158),
.Y(n_5269)
);

AND2x4_ASAP7_75t_L g5270 ( 
.A(n_5235),
.B(n_5248),
.Y(n_5270)
);

INVx1_ASAP7_75t_L g5271 ( 
.A(n_5226),
.Y(n_5271)
);

NAND2xp5_ASAP7_75t_L g5272 ( 
.A(n_5234),
.B(n_5167),
.Y(n_5272)
);

OR2x2_ASAP7_75t_L g5273 ( 
.A(n_5263),
.B(n_5226),
.Y(n_5273)
);

INVx1_ASAP7_75t_L g5274 ( 
.A(n_5257),
.Y(n_5274)
);

OR2x2_ASAP7_75t_L g5275 ( 
.A(n_5262),
.B(n_5229),
.Y(n_5275)
);

INVx2_ASAP7_75t_SL g5276 ( 
.A(n_5251),
.Y(n_5276)
);

NAND2xp5_ASAP7_75t_L g5277 ( 
.A(n_5264),
.B(n_5244),
.Y(n_5277)
);

BUFx2_ASAP7_75t_L g5278 ( 
.A(n_5253),
.Y(n_5278)
);

AND2x2_ASAP7_75t_L g5279 ( 
.A(n_5251),
.B(n_5249),
.Y(n_5279)
);

NOR2x1_ASAP7_75t_L g5280 ( 
.A(n_5250),
.B(n_5248),
.Y(n_5280)
);

INVx1_ASAP7_75t_L g5281 ( 
.A(n_5254),
.Y(n_5281)
);

INVx1_ASAP7_75t_L g5282 ( 
.A(n_5268),
.Y(n_5282)
);

OR2x2_ASAP7_75t_L g5283 ( 
.A(n_5263),
.B(n_5271),
.Y(n_5283)
);

AND2x2_ASAP7_75t_L g5284 ( 
.A(n_5255),
.B(n_5244),
.Y(n_5284)
);

NAND2xp5_ASAP7_75t_L g5285 ( 
.A(n_5270),
.B(n_5241),
.Y(n_5285)
);

INVx1_ASAP7_75t_L g5286 ( 
.A(n_5268),
.Y(n_5286)
);

INVx1_ASAP7_75t_L g5287 ( 
.A(n_5267),
.Y(n_5287)
);

INVx1_ASAP7_75t_L g5288 ( 
.A(n_5267),
.Y(n_5288)
);

AND2x2_ASAP7_75t_L g5289 ( 
.A(n_5255),
.B(n_5236),
.Y(n_5289)
);

BUFx2_ASAP7_75t_L g5290 ( 
.A(n_5253),
.Y(n_5290)
);

INVx2_ASAP7_75t_L g5291 ( 
.A(n_5250),
.Y(n_5291)
);

INVx1_ASAP7_75t_L g5292 ( 
.A(n_5266),
.Y(n_5292)
);

INVx2_ASAP7_75t_L g5293 ( 
.A(n_5252),
.Y(n_5293)
);

INVx1_ASAP7_75t_L g5294 ( 
.A(n_5266),
.Y(n_5294)
);

NAND2xp5_ASAP7_75t_L g5295 ( 
.A(n_5270),
.B(n_5241),
.Y(n_5295)
);

OAI22xp33_ASAP7_75t_L g5296 ( 
.A1(n_5273),
.A2(n_5271),
.B1(n_5259),
.B2(n_5260),
.Y(n_5296)
);

NOR4xp25_ASAP7_75t_SL g5297 ( 
.A(n_5278),
.B(n_5261),
.C(n_5290),
.D(n_5286),
.Y(n_5297)
);

NOR2xp33_ASAP7_75t_L g5298 ( 
.A(n_5285),
.B(n_5248),
.Y(n_5298)
);

CKINVDCx8_ASAP7_75t_R g5299 ( 
.A(n_5280),
.Y(n_5299)
);

BUFx3_ASAP7_75t_L g5300 ( 
.A(n_5287),
.Y(n_5300)
);

NAND2xp5_ASAP7_75t_L g5301 ( 
.A(n_5279),
.B(n_5270),
.Y(n_5301)
);

CKINVDCx5p33_ASAP7_75t_R g5302 ( 
.A(n_5288),
.Y(n_5302)
);

NAND2xp5_ASAP7_75t_L g5303 ( 
.A(n_5279),
.B(n_5253),
.Y(n_5303)
);

NAND2xp5_ASAP7_75t_L g5304 ( 
.A(n_5284),
.B(n_5269),
.Y(n_5304)
);

NOR2xp33_ASAP7_75t_L g5305 ( 
.A(n_5295),
.B(n_5269),
.Y(n_5305)
);

AO221x2_ASAP7_75t_L g5306 ( 
.A1(n_5282),
.A2(n_5252),
.B1(n_5258),
.B2(n_5260),
.C(n_5259),
.Y(n_5306)
);

CKINVDCx20_ASAP7_75t_R g5307 ( 
.A(n_5284),
.Y(n_5307)
);

NAND2xp5_ASAP7_75t_L g5308 ( 
.A(n_5289),
.B(n_5269),
.Y(n_5308)
);

NOR2x1_ASAP7_75t_L g5309 ( 
.A(n_5273),
.B(n_5258),
.Y(n_5309)
);

OAI221xp5_ASAP7_75t_L g5310 ( 
.A1(n_5283),
.A2(n_5187),
.B1(n_5202),
.B2(n_5239),
.C(n_5221),
.Y(n_5310)
);

NAND2xp5_ASAP7_75t_L g5311 ( 
.A(n_5289),
.B(n_5266),
.Y(n_5311)
);

NAND2xp5_ASAP7_75t_L g5312 ( 
.A(n_5276),
.B(n_5245),
.Y(n_5312)
);

INVx1_ASAP7_75t_SL g5313 ( 
.A(n_5307),
.Y(n_5313)
);

INVx1_ASAP7_75t_L g5314 ( 
.A(n_5309),
.Y(n_5314)
);

AND2x2_ASAP7_75t_L g5315 ( 
.A(n_5297),
.B(n_5276),
.Y(n_5315)
);

AND2x4_ASAP7_75t_L g5316 ( 
.A(n_5300),
.B(n_5274),
.Y(n_5316)
);

INVx2_ASAP7_75t_SL g5317 ( 
.A(n_5304),
.Y(n_5317)
);

NAND2xp5_ASAP7_75t_L g5318 ( 
.A(n_5306),
.B(n_5231),
.Y(n_5318)
);

INVx1_ASAP7_75t_L g5319 ( 
.A(n_5312),
.Y(n_5319)
);

INVx2_ASAP7_75t_L g5320 ( 
.A(n_5303),
.Y(n_5320)
);

AOI22xp33_ASAP7_75t_L g5321 ( 
.A1(n_5306),
.A2(n_5239),
.B1(n_5220),
.B2(n_5246),
.Y(n_5321)
);

AND2x2_ASAP7_75t_L g5322 ( 
.A(n_5305),
.B(n_5236),
.Y(n_5322)
);

AND2x2_ASAP7_75t_L g5323 ( 
.A(n_5308),
.B(n_5219),
.Y(n_5323)
);

OR2x2_ASAP7_75t_L g5324 ( 
.A(n_5301),
.B(n_5275),
.Y(n_5324)
);

AND2x2_ASAP7_75t_L g5325 ( 
.A(n_5313),
.B(n_5238),
.Y(n_5325)
);

AOI22xp5_ASAP7_75t_L g5326 ( 
.A1(n_5321),
.A2(n_5242),
.B1(n_5220),
.B2(n_5310),
.Y(n_5326)
);

INVxp67_ASAP7_75t_L g5327 ( 
.A(n_5315),
.Y(n_5327)
);

OAI21xp33_ASAP7_75t_L g5328 ( 
.A1(n_5313),
.A2(n_5272),
.B(n_5256),
.Y(n_5328)
);

AND2x2_ASAP7_75t_L g5329 ( 
.A(n_5322),
.B(n_5298),
.Y(n_5329)
);

NOR2xp33_ASAP7_75t_L g5330 ( 
.A(n_5317),
.B(n_5245),
.Y(n_5330)
);

NOR2x1p5_ASAP7_75t_SL g5331 ( 
.A(n_5324),
.B(n_5314),
.Y(n_5331)
);

AND2x2_ASAP7_75t_L g5332 ( 
.A(n_5323),
.B(n_5277),
.Y(n_5332)
);

OAI21xp5_ASAP7_75t_L g5333 ( 
.A1(n_5321),
.A2(n_5296),
.B(n_5311),
.Y(n_5333)
);

AOI22xp33_ASAP7_75t_L g5334 ( 
.A1(n_5318),
.A2(n_5200),
.B1(n_5242),
.B2(n_5246),
.Y(n_5334)
);

INVx1_ASAP7_75t_L g5335 ( 
.A(n_5316),
.Y(n_5335)
);

AND2x2_ASAP7_75t_L g5336 ( 
.A(n_5320),
.B(n_5302),
.Y(n_5336)
);

AND2x2_ASAP7_75t_L g5337 ( 
.A(n_5316),
.B(n_5281),
.Y(n_5337)
);

INVx1_ASAP7_75t_L g5338 ( 
.A(n_5319),
.Y(n_5338)
);

NAND2xp5_ASAP7_75t_SL g5339 ( 
.A(n_5318),
.B(n_5245),
.Y(n_5339)
);

INVx1_ASAP7_75t_L g5340 ( 
.A(n_5325),
.Y(n_5340)
);

AND2x2_ASAP7_75t_L g5341 ( 
.A(n_5332),
.B(n_5265),
.Y(n_5341)
);

NAND2xp5_ASAP7_75t_L g5342 ( 
.A(n_5331),
.B(n_5245),
.Y(n_5342)
);

OAI21xp5_ASAP7_75t_L g5343 ( 
.A1(n_5327),
.A2(n_5246),
.B(n_5242),
.Y(n_5343)
);

INVx1_ASAP7_75t_L g5344 ( 
.A(n_5330),
.Y(n_5344)
);

OAI21xp33_ASAP7_75t_L g5345 ( 
.A1(n_5328),
.A2(n_5247),
.B(n_5240),
.Y(n_5345)
);

INVx1_ASAP7_75t_L g5346 ( 
.A(n_5337),
.Y(n_5346)
);

OAI21xp33_ASAP7_75t_L g5347 ( 
.A1(n_5329),
.A2(n_5222),
.B(n_5229),
.Y(n_5347)
);

OAI22xp33_ASAP7_75t_L g5348 ( 
.A1(n_5326),
.A2(n_5201),
.B1(n_5222),
.B2(n_5243),
.Y(n_5348)
);

NOR2xp67_ASAP7_75t_SL g5349 ( 
.A(n_5335),
.B(n_5299),
.Y(n_5349)
);

OR2x2_ASAP7_75t_L g5350 ( 
.A(n_5339),
.B(n_5218),
.Y(n_5350)
);

AOI22xp5_ASAP7_75t_L g5351 ( 
.A1(n_5334),
.A2(n_5224),
.B1(n_5232),
.B2(n_5243),
.Y(n_5351)
);

INVxp67_ASAP7_75t_L g5352 ( 
.A(n_5342),
.Y(n_5352)
);

INVx1_ASAP7_75t_L g5353 ( 
.A(n_5347),
.Y(n_5353)
);

NOR2xp33_ASAP7_75t_L g5354 ( 
.A(n_5345),
.B(n_5327),
.Y(n_5354)
);

NAND2xp5_ASAP7_75t_L g5355 ( 
.A(n_5341),
.B(n_5336),
.Y(n_5355)
);

INVx1_ASAP7_75t_L g5356 ( 
.A(n_5343),
.Y(n_5356)
);

INVx1_ASAP7_75t_L g5357 ( 
.A(n_5350),
.Y(n_5357)
);

NOR2xp33_ASAP7_75t_L g5358 ( 
.A(n_5340),
.B(n_5243),
.Y(n_5358)
);

NAND2xp5_ASAP7_75t_L g5359 ( 
.A(n_5346),
.B(n_5291),
.Y(n_5359)
);

NAND2xp5_ASAP7_75t_L g5360 ( 
.A(n_5349),
.B(n_5291),
.Y(n_5360)
);

NAND2xp5_ASAP7_75t_SL g5361 ( 
.A(n_5348),
.B(n_5333),
.Y(n_5361)
);

INVx1_ASAP7_75t_L g5362 ( 
.A(n_5351),
.Y(n_5362)
);

NAND2xp5_ASAP7_75t_L g5363 ( 
.A(n_5358),
.B(n_5293),
.Y(n_5363)
);

AOI22xp5_ASAP7_75t_L g5364 ( 
.A1(n_5352),
.A2(n_5293),
.B1(n_5333),
.B2(n_5232),
.Y(n_5364)
);

NAND2xp5_ASAP7_75t_L g5365 ( 
.A(n_5355),
.B(n_5224),
.Y(n_5365)
);

HB1xp67_ASAP7_75t_L g5366 ( 
.A(n_5360),
.Y(n_5366)
);

AOI222xp33_ASAP7_75t_L g5367 ( 
.A1(n_5361),
.A2(n_5356),
.B1(n_5362),
.B2(n_5359),
.C1(n_5354),
.C2(n_5357),
.Y(n_5367)
);

INVx1_ASAP7_75t_L g5368 ( 
.A(n_5353),
.Y(n_5368)
);

OAI21xp5_ASAP7_75t_L g5369 ( 
.A1(n_5361),
.A2(n_5338),
.B(n_5344),
.Y(n_5369)
);

AOI22xp5_ASAP7_75t_L g5370 ( 
.A1(n_5352),
.A2(n_5175),
.B1(n_5294),
.B2(n_5292),
.Y(n_5370)
);

INVx1_ASAP7_75t_L g5371 ( 
.A(n_5360),
.Y(n_5371)
);

NAND2xp5_ASAP7_75t_L g5372 ( 
.A(n_5358),
.B(n_5175),
.Y(n_5372)
);

NOR2x1_ASAP7_75t_L g5373 ( 
.A(n_5360),
.B(n_5218),
.Y(n_5373)
);

INVxp67_ASAP7_75t_SL g5374 ( 
.A(n_5361),
.Y(n_5374)
);

INVx1_ASAP7_75t_L g5375 ( 
.A(n_5360),
.Y(n_5375)
);

AND2x2_ASAP7_75t_L g5376 ( 
.A(n_5357),
.B(n_5158),
.Y(n_5376)
);

INVx1_ASAP7_75t_L g5377 ( 
.A(n_5360),
.Y(n_5377)
);

INVx1_ASAP7_75t_L g5378 ( 
.A(n_5360),
.Y(n_5378)
);

NAND2xp5_ASAP7_75t_L g5379 ( 
.A(n_5358),
.B(n_5170),
.Y(n_5379)
);

NAND2xp33_ASAP7_75t_SL g5380 ( 
.A(n_5355),
.B(n_5214),
.Y(n_5380)
);

AOI22xp33_ASAP7_75t_L g5381 ( 
.A1(n_5352),
.A2(n_5152),
.B1(n_5111),
.B2(n_5132),
.Y(n_5381)
);

HB1xp67_ASAP7_75t_L g5382 ( 
.A(n_5373),
.Y(n_5382)
);

INVx1_ASAP7_75t_L g5383 ( 
.A(n_5374),
.Y(n_5383)
);

INVx2_ASAP7_75t_L g5384 ( 
.A(n_5376),
.Y(n_5384)
);

INVx3_ASAP7_75t_L g5385 ( 
.A(n_5368),
.Y(n_5385)
);

INVx1_ASAP7_75t_L g5386 ( 
.A(n_5363),
.Y(n_5386)
);

INVx1_ASAP7_75t_SL g5387 ( 
.A(n_5365),
.Y(n_5387)
);

INVx2_ASAP7_75t_L g5388 ( 
.A(n_5366),
.Y(n_5388)
);

NAND2xp5_ASAP7_75t_L g5389 ( 
.A(n_5364),
.B(n_5170),
.Y(n_5389)
);

INVx1_ASAP7_75t_L g5390 ( 
.A(n_5372),
.Y(n_5390)
);

INVx1_ASAP7_75t_L g5391 ( 
.A(n_5379),
.Y(n_5391)
);

INVx2_ASAP7_75t_L g5392 ( 
.A(n_5371),
.Y(n_5392)
);

HB1xp67_ASAP7_75t_L g5393 ( 
.A(n_5369),
.Y(n_5393)
);

INVx1_ASAP7_75t_SL g5394 ( 
.A(n_5375),
.Y(n_5394)
);

INVx2_ASAP7_75t_L g5395 ( 
.A(n_5377),
.Y(n_5395)
);

BUFx4f_ASAP7_75t_SL g5396 ( 
.A(n_5378),
.Y(n_5396)
);

INVx2_ASAP7_75t_L g5397 ( 
.A(n_5370),
.Y(n_5397)
);

INVx1_ASAP7_75t_L g5398 ( 
.A(n_5367),
.Y(n_5398)
);

INVx1_ASAP7_75t_L g5399 ( 
.A(n_5380),
.Y(n_5399)
);

INVx1_ASAP7_75t_L g5400 ( 
.A(n_5381),
.Y(n_5400)
);

INVx1_ASAP7_75t_L g5401 ( 
.A(n_5374),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_5374),
.Y(n_5402)
);

BUFx2_ASAP7_75t_L g5403 ( 
.A(n_5374),
.Y(n_5403)
);

OR2x2_ASAP7_75t_L g5404 ( 
.A(n_5374),
.B(n_5156),
.Y(n_5404)
);

INVx1_ASAP7_75t_L g5405 ( 
.A(n_5374),
.Y(n_5405)
);

INVx1_ASAP7_75t_L g5406 ( 
.A(n_5374),
.Y(n_5406)
);

OAI22xp5_ASAP7_75t_L g5407 ( 
.A1(n_5394),
.A2(n_5156),
.B1(n_5102),
.B2(n_5154),
.Y(n_5407)
);

AOI21xp33_ASAP7_75t_L g5408 ( 
.A1(n_5382),
.A2(n_5111),
.B(n_5133),
.Y(n_5408)
);

AOI221x1_ASAP7_75t_SL g5409 ( 
.A1(n_5398),
.A2(n_5197),
.B1(n_5195),
.B2(n_5211),
.C(n_5107),
.Y(n_5409)
);

XNOR2x1_ASAP7_75t_L g5410 ( 
.A(n_5404),
.B(n_5111),
.Y(n_5410)
);

AOI221xp5_ASAP7_75t_L g5411 ( 
.A1(n_5382),
.A2(n_5187),
.B1(n_5202),
.B2(n_5213),
.C(n_5196),
.Y(n_5411)
);

O2A1O1Ixp33_ASAP7_75t_L g5412 ( 
.A1(n_5393),
.A2(n_5196),
.B(n_5122),
.C(n_5134),
.Y(n_5412)
);

INVx2_ASAP7_75t_L g5413 ( 
.A(n_5403),
.Y(n_5413)
);

NAND2xp5_ASAP7_75t_L g5414 ( 
.A(n_5387),
.B(n_5144),
.Y(n_5414)
);

XOR2xp5_ASAP7_75t_L g5415 ( 
.A(n_5383),
.B(n_5215),
.Y(n_5415)
);

AOI221xp5_ASAP7_75t_L g5416 ( 
.A1(n_5394),
.A2(n_5210),
.B1(n_5111),
.B2(n_5122),
.C(n_5123),
.Y(n_5416)
);

AOI21xp5_ASAP7_75t_L g5417 ( 
.A1(n_5401),
.A2(n_5102),
.B(n_5123),
.Y(n_5417)
);

INVx1_ASAP7_75t_SL g5418 ( 
.A(n_5387),
.Y(n_5418)
);

AOI22xp5_ASAP7_75t_L g5419 ( 
.A1(n_5385),
.A2(n_5134),
.B1(n_5135),
.B2(n_5141),
.Y(n_5419)
);

OAI321xp33_ASAP7_75t_L g5420 ( 
.A1(n_5402),
.A2(n_5133),
.A3(n_5135),
.B1(n_5144),
.B2(n_5127),
.C(n_5118),
.Y(n_5420)
);

AOI221xp5_ASAP7_75t_L g5421 ( 
.A1(n_5385),
.A2(n_5118),
.B1(n_5128),
.B2(n_5117),
.C(n_5161),
.Y(n_5421)
);

NOR4xp25_ASAP7_75t_L g5422 ( 
.A(n_5405),
.B(n_5127),
.C(n_5128),
.D(n_5147),
.Y(n_5422)
);

INVx1_ASAP7_75t_L g5423 ( 
.A(n_5406),
.Y(n_5423)
);

AOI22xp5_ASAP7_75t_L g5424 ( 
.A1(n_5388),
.A2(n_5141),
.B1(n_5147),
.B2(n_5131),
.Y(n_5424)
);

INVx1_ASAP7_75t_SL g5425 ( 
.A(n_5396),
.Y(n_5425)
);

NOR4xp25_ASAP7_75t_L g5426 ( 
.A(n_5399),
.B(n_5395),
.C(n_5392),
.D(n_5400),
.Y(n_5426)
);

NOR3xp33_ASAP7_75t_L g5427 ( 
.A(n_5386),
.B(n_5165),
.C(n_5131),
.Y(n_5427)
);

AOI221xp5_ASAP7_75t_L g5428 ( 
.A1(n_5389),
.A2(n_5391),
.B1(n_5390),
.B2(n_5397),
.C(n_5384),
.Y(n_5428)
);

AND2x2_ASAP7_75t_L g5429 ( 
.A(n_5389),
.B(n_5124),
.Y(n_5429)
);

INVx1_ASAP7_75t_SL g5430 ( 
.A(n_5403),
.Y(n_5430)
);

AOI21xp5_ASAP7_75t_L g5431 ( 
.A1(n_5382),
.A2(n_5115),
.B(n_5149),
.Y(n_5431)
);

AOI21xp5_ASAP7_75t_L g5432 ( 
.A1(n_5382),
.A2(n_5115),
.B(n_5149),
.Y(n_5432)
);

AOI22xp5_ASAP7_75t_L g5433 ( 
.A1(n_5393),
.A2(n_5159),
.B1(n_5124),
.B2(n_5168),
.Y(n_5433)
);

OR2x2_ASAP7_75t_L g5434 ( 
.A(n_5403),
.B(n_5159),
.Y(n_5434)
);

OAI321xp33_ASAP7_75t_L g5435 ( 
.A1(n_5414),
.A2(n_5148),
.A3(n_5168),
.B1(n_406),
.B2(n_407),
.C(n_408),
.Y(n_5435)
);

OAI211xp5_ASAP7_75t_L g5436 ( 
.A1(n_5430),
.A2(n_408),
.B(n_403),
.C(n_405),
.Y(n_5436)
);

NAND2xp5_ASAP7_75t_L g5437 ( 
.A(n_5431),
.B(n_5148),
.Y(n_5437)
);

AOI221xp5_ASAP7_75t_L g5438 ( 
.A1(n_5426),
.A2(n_409),
.B1(n_410),
.B2(n_411),
.C(n_412),
.Y(n_5438)
);

OAI211xp5_ASAP7_75t_SL g5439 ( 
.A1(n_5418),
.A2(n_412),
.B(n_409),
.C(n_411),
.Y(n_5439)
);

AOI22xp5_ASAP7_75t_L g5440 ( 
.A1(n_5413),
.A2(n_413),
.B1(n_415),
.B2(n_416),
.Y(n_5440)
);

AOI221xp5_ASAP7_75t_L g5441 ( 
.A1(n_5408),
.A2(n_418),
.B1(n_419),
.B2(n_420),
.C(n_421),
.Y(n_5441)
);

NAND4xp25_ASAP7_75t_SL g5442 ( 
.A(n_5425),
.B(n_418),
.C(n_422),
.D(n_423),
.Y(n_5442)
);

OAI211xp5_ASAP7_75t_SL g5443 ( 
.A1(n_5428),
.A2(n_422),
.B(n_423),
.C(n_424),
.Y(n_5443)
);

OAI221xp5_ASAP7_75t_SL g5444 ( 
.A1(n_5434),
.A2(n_425),
.B1(n_426),
.B2(n_427),
.C(n_428),
.Y(n_5444)
);

AOI22xp5_ASAP7_75t_L g5445 ( 
.A1(n_5423),
.A2(n_425),
.B1(n_426),
.B2(n_427),
.Y(n_5445)
);

AOI22xp33_ASAP7_75t_L g5446 ( 
.A1(n_5410),
.A2(n_428),
.B1(n_429),
.B2(n_430),
.Y(n_5446)
);

AOI221x1_ASAP7_75t_L g5447 ( 
.A1(n_5417),
.A2(n_430),
.B1(n_431),
.B2(n_432),
.C(n_433),
.Y(n_5447)
);

INVx1_ASAP7_75t_SL g5448 ( 
.A(n_5429),
.Y(n_5448)
);

OAI21xp5_ASAP7_75t_SL g5449 ( 
.A1(n_5415),
.A2(n_431),
.B(n_432),
.Y(n_5449)
);

AOI221x1_ASAP7_75t_L g5450 ( 
.A1(n_5407),
.A2(n_433),
.B1(n_436),
.B2(n_438),
.C(n_439),
.Y(n_5450)
);

OAI222xp33_ASAP7_75t_L g5451 ( 
.A1(n_5424),
.A2(n_436),
.B1(n_438),
.B2(n_440),
.C1(n_442),
.C2(n_443),
.Y(n_5451)
);

NAND2xp5_ASAP7_75t_SL g5452 ( 
.A(n_5427),
.B(n_443),
.Y(n_5452)
);

AOI211xp5_ASAP7_75t_L g5453 ( 
.A1(n_5412),
.A2(n_445),
.B(n_446),
.C(n_449),
.Y(n_5453)
);

NAND3xp33_ASAP7_75t_SL g5454 ( 
.A(n_5411),
.B(n_445),
.C(n_446),
.Y(n_5454)
);

OAI22xp33_ASAP7_75t_L g5455 ( 
.A1(n_5419),
.A2(n_449),
.B1(n_453),
.B2(n_454),
.Y(n_5455)
);

NOR2xp33_ASAP7_75t_L g5456 ( 
.A(n_5432),
.B(n_453),
.Y(n_5456)
);

AOI221xp5_ASAP7_75t_L g5457 ( 
.A1(n_5422),
.A2(n_456),
.B1(n_457),
.B2(n_460),
.C(n_461),
.Y(n_5457)
);

AOI211xp5_ASAP7_75t_L g5458 ( 
.A1(n_5420),
.A2(n_460),
.B(n_461),
.C(n_462),
.Y(n_5458)
);

AND2x2_ASAP7_75t_L g5459 ( 
.A(n_5448),
.B(n_5433),
.Y(n_5459)
);

NOR2xp33_ASAP7_75t_L g5460 ( 
.A(n_5435),
.B(n_5421),
.Y(n_5460)
);

AOI221xp5_ASAP7_75t_L g5461 ( 
.A1(n_5456),
.A2(n_5416),
.B1(n_5409),
.B2(n_464),
.C(n_465),
.Y(n_5461)
);

OAI211xp5_ASAP7_75t_L g5462 ( 
.A1(n_5438),
.A2(n_462),
.B(n_463),
.C(n_464),
.Y(n_5462)
);

INVx1_ASAP7_75t_SL g5463 ( 
.A(n_5452),
.Y(n_5463)
);

AOI22xp5_ASAP7_75t_L g5464 ( 
.A1(n_5437),
.A2(n_465),
.B1(n_468),
.B2(n_469),
.Y(n_5464)
);

OAI21xp5_ASAP7_75t_SL g5465 ( 
.A1(n_5439),
.A2(n_468),
.B(n_469),
.Y(n_5465)
);

NOR3xp33_ASAP7_75t_L g5466 ( 
.A(n_5451),
.B(n_471),
.C(n_472),
.Y(n_5466)
);

OAI211xp5_ASAP7_75t_SL g5467 ( 
.A1(n_5458),
.A2(n_471),
.B(n_473),
.C(n_476),
.Y(n_5467)
);

AOI21xp5_ASAP7_75t_L g5468 ( 
.A1(n_5457),
.A2(n_473),
.B(n_476),
.Y(n_5468)
);

AOI22xp33_ASAP7_75t_L g5469 ( 
.A1(n_5443),
.A2(n_477),
.B1(n_478),
.B2(n_479),
.Y(n_5469)
);

AO22x2_ASAP7_75t_L g5470 ( 
.A1(n_5454),
.A2(n_478),
.B1(n_480),
.B2(n_481),
.Y(n_5470)
);

OAI211xp5_ASAP7_75t_L g5471 ( 
.A1(n_5450),
.A2(n_480),
.B(n_482),
.C(n_484),
.Y(n_5471)
);

AOI22xp5_ASAP7_75t_L g5472 ( 
.A1(n_5446),
.A2(n_482),
.B1(n_485),
.B2(n_488),
.Y(n_5472)
);

AOI221xp5_ASAP7_75t_L g5473 ( 
.A1(n_5449),
.A2(n_485),
.B1(n_489),
.B2(n_490),
.C(n_492),
.Y(n_5473)
);

NAND3xp33_ASAP7_75t_L g5474 ( 
.A(n_5441),
.B(n_489),
.C(n_490),
.Y(n_5474)
);

NOR3xp33_ASAP7_75t_L g5475 ( 
.A(n_5436),
.B(n_5442),
.C(n_5444),
.Y(n_5475)
);

OA22x2_ASAP7_75t_L g5476 ( 
.A1(n_5447),
.A2(n_492),
.B1(n_493),
.B2(n_494),
.Y(n_5476)
);

OR2x2_ASAP7_75t_L g5477 ( 
.A(n_5465),
.B(n_5463),
.Y(n_5477)
);

AOI22xp5_ASAP7_75t_L g5478 ( 
.A1(n_5460),
.A2(n_5453),
.B1(n_5440),
.B2(n_5455),
.Y(n_5478)
);

INVx1_ASAP7_75t_L g5479 ( 
.A(n_5476),
.Y(n_5479)
);

AOI22xp5_ASAP7_75t_L g5480 ( 
.A1(n_5475),
.A2(n_5445),
.B1(n_495),
.B2(n_496),
.Y(n_5480)
);

INVx1_ASAP7_75t_L g5481 ( 
.A(n_5470),
.Y(n_5481)
);

NOR2x2_ASAP7_75t_L g5482 ( 
.A(n_5470),
.B(n_5471),
.Y(n_5482)
);

NAND2xp5_ASAP7_75t_L g5483 ( 
.A(n_5459),
.B(n_5461),
.Y(n_5483)
);

INVx1_ASAP7_75t_L g5484 ( 
.A(n_5467),
.Y(n_5484)
);

INVx1_ASAP7_75t_L g5485 ( 
.A(n_5466),
.Y(n_5485)
);

INVx1_ASAP7_75t_L g5486 ( 
.A(n_5472),
.Y(n_5486)
);

INVx1_ASAP7_75t_L g5487 ( 
.A(n_5464),
.Y(n_5487)
);

INVx1_ASAP7_75t_L g5488 ( 
.A(n_5462),
.Y(n_5488)
);

INVx1_ASAP7_75t_L g5489 ( 
.A(n_5474),
.Y(n_5489)
);

AOI22xp5_ASAP7_75t_L g5490 ( 
.A1(n_5469),
.A2(n_494),
.B1(n_498),
.B2(n_499),
.Y(n_5490)
);

AOI22xp5_ASAP7_75t_L g5491 ( 
.A1(n_5473),
.A2(n_5468),
.B1(n_499),
.B2(n_500),
.Y(n_5491)
);

NOR2xp33_ASAP7_75t_L g5492 ( 
.A(n_5459),
.B(n_498),
.Y(n_5492)
);

OAI21xp5_ASAP7_75t_SL g5493 ( 
.A1(n_5479),
.A2(n_500),
.B(n_501),
.Y(n_5493)
);

AND2x2_ASAP7_75t_L g5494 ( 
.A(n_5481),
.B(n_501),
.Y(n_5494)
);

OR5x1_ASAP7_75t_L g5495 ( 
.A(n_5482),
.B(n_502),
.C(n_503),
.D(n_504),
.E(n_506),
.Y(n_5495)
);

AOI221xp5_ASAP7_75t_L g5496 ( 
.A1(n_5484),
.A2(n_502),
.B1(n_506),
.B2(n_508),
.C(n_509),
.Y(n_5496)
);

AND2x2_ASAP7_75t_L g5497 ( 
.A(n_5492),
.B(n_508),
.Y(n_5497)
);

OR2x2_ASAP7_75t_L g5498 ( 
.A(n_5477),
.B(n_509),
.Y(n_5498)
);

XNOR2xp5_ASAP7_75t_L g5499 ( 
.A(n_5478),
.B(n_5483),
.Y(n_5499)
);

NAND2xp5_ASAP7_75t_L g5500 ( 
.A(n_5485),
.B(n_511),
.Y(n_5500)
);

NOR2x1_ASAP7_75t_L g5501 ( 
.A(n_5488),
.B(n_511),
.Y(n_5501)
);

NAND2xp33_ASAP7_75t_R g5502 ( 
.A(n_5489),
.B(n_512),
.Y(n_5502)
);

AOI22xp5_ASAP7_75t_L g5503 ( 
.A1(n_5480),
.A2(n_512),
.B1(n_513),
.B2(n_514),
.Y(n_5503)
);

NAND3xp33_ASAP7_75t_L g5504 ( 
.A(n_5486),
.B(n_513),
.C(n_515),
.Y(n_5504)
);

NOR3xp33_ASAP7_75t_L g5505 ( 
.A(n_5487),
.B(n_515),
.C(n_516),
.Y(n_5505)
);

AND2x4_ASAP7_75t_L g5506 ( 
.A(n_5491),
.B(n_5490),
.Y(n_5506)
);

INVxp67_ASAP7_75t_L g5507 ( 
.A(n_5492),
.Y(n_5507)
);

INVx1_ASAP7_75t_L g5508 ( 
.A(n_5481),
.Y(n_5508)
);

NAND3xp33_ASAP7_75t_L g5509 ( 
.A(n_5481),
.B(n_516),
.C(n_518),
.Y(n_5509)
);

NAND4xp25_ASAP7_75t_SL g5510 ( 
.A(n_5483),
.B(n_518),
.C(n_519),
.D(n_521),
.Y(n_5510)
);

XNOR2xp5_ASAP7_75t_L g5511 ( 
.A(n_5499),
.B(n_5495),
.Y(n_5511)
);

NOR2xp33_ASAP7_75t_R g5512 ( 
.A(n_5502),
.B(n_519),
.Y(n_5512)
);

NOR2xp33_ASAP7_75t_R g5513 ( 
.A(n_5508),
.B(n_521),
.Y(n_5513)
);

NOR2xp33_ASAP7_75t_R g5514 ( 
.A(n_5510),
.B(n_5500),
.Y(n_5514)
);

NOR3xp33_ASAP7_75t_SL g5515 ( 
.A(n_5493),
.B(n_523),
.C(n_525),
.Y(n_5515)
);

NAND2xp33_ASAP7_75t_SL g5516 ( 
.A(n_5498),
.B(n_523),
.Y(n_5516)
);

NOR2xp33_ASAP7_75t_R g5517 ( 
.A(n_5494),
.B(n_5497),
.Y(n_5517)
);

NOR2xp33_ASAP7_75t_R g5518 ( 
.A(n_5507),
.B(n_525),
.Y(n_5518)
);

NAND2xp5_ASAP7_75t_L g5519 ( 
.A(n_5501),
.B(n_526),
.Y(n_5519)
);

NAND2xp5_ASAP7_75t_SL g5520 ( 
.A(n_5505),
.B(n_526),
.Y(n_5520)
);

NOR2xp33_ASAP7_75t_R g5521 ( 
.A(n_5506),
.B(n_527),
.Y(n_5521)
);

NOR2xp33_ASAP7_75t_R g5522 ( 
.A(n_5506),
.B(n_527),
.Y(n_5522)
);

NAND2xp5_ASAP7_75t_SL g5523 ( 
.A(n_5509),
.B(n_530),
.Y(n_5523)
);

AOI22xp5_ASAP7_75t_L g5524 ( 
.A1(n_5511),
.A2(n_5503),
.B1(n_5504),
.B2(n_5496),
.Y(n_5524)
);

NOR3xp33_ASAP7_75t_L g5525 ( 
.A(n_5516),
.B(n_531),
.C(n_532),
.Y(n_5525)
);

AOI21xp5_ASAP7_75t_L g5526 ( 
.A1(n_5519),
.A2(n_532),
.B(n_533),
.Y(n_5526)
);

OR2x6_ASAP7_75t_L g5527 ( 
.A(n_5517),
.B(n_533),
.Y(n_5527)
);

AND4x1_ASAP7_75t_L g5528 ( 
.A(n_5515),
.B(n_534),
.C(n_535),
.D(n_536),
.Y(n_5528)
);

NAND2xp5_ASAP7_75t_L g5529 ( 
.A(n_5512),
.B(n_535),
.Y(n_5529)
);

NOR3xp33_ASAP7_75t_L g5530 ( 
.A(n_5520),
.B(n_536),
.C(n_537),
.Y(n_5530)
);

BUFx2_ASAP7_75t_L g5531 ( 
.A(n_5527),
.Y(n_5531)
);

BUFx2_ASAP7_75t_L g5532 ( 
.A(n_5529),
.Y(n_5532)
);

OAI222xp33_ASAP7_75t_L g5533 ( 
.A1(n_5524),
.A2(n_5523),
.B1(n_5514),
.B2(n_5513),
.C1(n_5522),
.C2(n_5521),
.Y(n_5533)
);

XOR2xp5_ASAP7_75t_L g5534 ( 
.A(n_5526),
.B(n_5518),
.Y(n_5534)
);

CKINVDCx5p33_ASAP7_75t_R g5535 ( 
.A(n_5528),
.Y(n_5535)
);

INVx1_ASAP7_75t_L g5536 ( 
.A(n_5525),
.Y(n_5536)
);

HB1xp67_ASAP7_75t_L g5537 ( 
.A(n_5530),
.Y(n_5537)
);

INVx1_ASAP7_75t_L g5538 ( 
.A(n_5531),
.Y(n_5538)
);

INVx2_ASAP7_75t_L g5539 ( 
.A(n_5535),
.Y(n_5539)
);

OAI21xp5_ASAP7_75t_L g5540 ( 
.A1(n_5533),
.A2(n_5534),
.B(n_5532),
.Y(n_5540)
);

NAND2xp5_ASAP7_75t_SL g5541 ( 
.A(n_5536),
.B(n_538),
.Y(n_5541)
);

NAND3xp33_ASAP7_75t_L g5542 ( 
.A(n_5537),
.B(n_538),
.C(n_539),
.Y(n_5542)
);

XNOR2xp5_ASAP7_75t_L g5543 ( 
.A(n_5534),
.B(n_541),
.Y(n_5543)
);

XOR2x1_ASAP7_75t_L g5544 ( 
.A(n_5538),
.B(n_541),
.Y(n_5544)
);

AOI21xp5_ASAP7_75t_L g5545 ( 
.A1(n_5540),
.A2(n_542),
.B(n_543),
.Y(n_5545)
);

INVx2_ASAP7_75t_L g5546 ( 
.A(n_5539),
.Y(n_5546)
);

OA22x2_ASAP7_75t_L g5547 ( 
.A1(n_5543),
.A2(n_544),
.B1(n_545),
.B2(n_546),
.Y(n_5547)
);

INVx1_ASAP7_75t_L g5548 ( 
.A(n_5541),
.Y(n_5548)
);

NAND2xp5_ASAP7_75t_L g5549 ( 
.A(n_5546),
.B(n_5542),
.Y(n_5549)
);

INVxp67_ASAP7_75t_SL g5550 ( 
.A(n_5548),
.Y(n_5550)
);

INVx4_ASAP7_75t_L g5551 ( 
.A(n_5544),
.Y(n_5551)
);

AOI22x1_ASAP7_75t_L g5552 ( 
.A1(n_5545),
.A2(n_5547),
.B1(n_549),
.B2(n_550),
.Y(n_5552)
);

AOI31xp33_ASAP7_75t_L g5553 ( 
.A1(n_5550),
.A2(n_548),
.A3(n_549),
.B(n_550),
.Y(n_5553)
);

AOI22xp33_ASAP7_75t_L g5554 ( 
.A1(n_5551),
.A2(n_548),
.B1(n_551),
.B2(n_552),
.Y(n_5554)
);

AOI22xp33_ASAP7_75t_L g5555 ( 
.A1(n_5552),
.A2(n_551),
.B1(n_552),
.B2(n_553),
.Y(n_5555)
);

AOI22xp33_ASAP7_75t_L g5556 ( 
.A1(n_5549),
.A2(n_554),
.B1(n_555),
.B2(n_556),
.Y(n_5556)
);

AOI22xp33_ASAP7_75t_L g5557 ( 
.A1(n_5550),
.A2(n_554),
.B1(n_555),
.B2(n_556),
.Y(n_5557)
);

INVx1_ASAP7_75t_SL g5558 ( 
.A(n_5555),
.Y(n_5558)
);

INVx1_ASAP7_75t_L g5559 ( 
.A(n_5553),
.Y(n_5559)
);

OAI22x1_ASAP7_75t_L g5560 ( 
.A1(n_5554),
.A2(n_558),
.B1(n_559),
.B2(n_560),
.Y(n_5560)
);

INVx1_ASAP7_75t_L g5561 ( 
.A(n_5557),
.Y(n_5561)
);

OR2x6_ASAP7_75t_L g5562 ( 
.A(n_5556),
.B(n_559),
.Y(n_5562)
);

INVx3_ASAP7_75t_L g5563 ( 
.A(n_5553),
.Y(n_5563)
);

INVxp67_ASAP7_75t_L g5564 ( 
.A(n_5555),
.Y(n_5564)
);

XNOR2xp5_ASAP7_75t_L g5565 ( 
.A(n_5555),
.B(n_563),
.Y(n_5565)
);

AOI22xp5_ASAP7_75t_L g5566 ( 
.A1(n_5555),
.A2(n_563),
.B1(n_564),
.B2(n_565),
.Y(n_5566)
);

AOI22xp5_ASAP7_75t_L g5567 ( 
.A1(n_5555),
.A2(n_565),
.B1(n_567),
.B2(n_569),
.Y(n_5567)
);

NAND3xp33_ASAP7_75t_L g5568 ( 
.A(n_5559),
.B(n_567),
.C(n_569),
.Y(n_5568)
);

AOI21xp5_ASAP7_75t_SL g5569 ( 
.A1(n_5564),
.A2(n_570),
.B(n_571),
.Y(n_5569)
);

A2O1A1O1Ixp25_ASAP7_75t_L g5570 ( 
.A1(n_5561),
.A2(n_570),
.B(n_572),
.C(n_573),
.D(n_574),
.Y(n_5570)
);

INVx1_ASAP7_75t_L g5571 ( 
.A(n_5563),
.Y(n_5571)
);

OR2x6_ASAP7_75t_L g5572 ( 
.A(n_5562),
.B(n_573),
.Y(n_5572)
);

AOI22xp5_ASAP7_75t_SL g5573 ( 
.A1(n_5558),
.A2(n_574),
.B1(n_576),
.B2(n_577),
.Y(n_5573)
);

OR2x2_ASAP7_75t_L g5574 ( 
.A(n_5560),
.B(n_576),
.Y(n_5574)
);

OAI21xp5_ASAP7_75t_SL g5575 ( 
.A1(n_5565),
.A2(n_578),
.B(n_579),
.Y(n_5575)
);

OR2x6_ASAP7_75t_L g5576 ( 
.A(n_5566),
.B(n_578),
.Y(n_5576)
);

AOI22xp33_ASAP7_75t_L g5577 ( 
.A1(n_5567),
.A2(n_580),
.B1(n_581),
.B2(n_582),
.Y(n_5577)
);

AOI22xp33_ASAP7_75t_L g5578 ( 
.A1(n_5571),
.A2(n_580),
.B1(n_581),
.B2(n_582),
.Y(n_5578)
);

AOI21xp5_ASAP7_75t_L g5579 ( 
.A1(n_5572),
.A2(n_5575),
.B(n_5569),
.Y(n_5579)
);

AOI222xp33_ASAP7_75t_SL g5580 ( 
.A1(n_5570),
.A2(n_583),
.B1(n_584),
.B2(n_586),
.C1(n_587),
.C2(n_588),
.Y(n_5580)
);

OAI22xp33_ASAP7_75t_SL g5581 ( 
.A1(n_5574),
.A2(n_584),
.B1(n_586),
.B2(n_587),
.Y(n_5581)
);

AOI22xp5_ASAP7_75t_SL g5582 ( 
.A1(n_5576),
.A2(n_5573),
.B1(n_5568),
.B2(n_5577),
.Y(n_5582)
);

INVx1_ASAP7_75t_L g5583 ( 
.A(n_5571),
.Y(n_5583)
);

AOI22xp5_ASAP7_75t_L g5584 ( 
.A1(n_5571),
.A2(n_589),
.B1(n_590),
.B2(n_591),
.Y(n_5584)
);

INVx1_ASAP7_75t_L g5585 ( 
.A(n_5571),
.Y(n_5585)
);

AOI21xp33_ASAP7_75t_L g5586 ( 
.A1(n_5583),
.A2(n_589),
.B(n_592),
.Y(n_5586)
);

AOI21xp33_ASAP7_75t_L g5587 ( 
.A1(n_5585),
.A2(n_594),
.B(n_595),
.Y(n_5587)
);

OR2x2_ASAP7_75t_L g5588 ( 
.A(n_5579),
.B(n_596),
.Y(n_5588)
);

FAx1_ASAP7_75t_L g5589 ( 
.A(n_5584),
.B(n_5582),
.CI(n_5580),
.CON(n_5589),
.SN(n_5589)
);

OR2x2_ASAP7_75t_L g5590 ( 
.A(n_5578),
.B(n_597),
.Y(n_5590)
);

OA331x2_ASAP7_75t_L g5591 ( 
.A1(n_5589),
.A2(n_5581),
.A3(n_600),
.B1(n_601),
.B2(n_602),
.B3(n_603),
.C1(n_604),
.Y(n_5591)
);

HB1xp67_ASAP7_75t_L g5592 ( 
.A(n_5588),
.Y(n_5592)
);

OAI221xp5_ASAP7_75t_R g5593 ( 
.A1(n_5592),
.A2(n_5590),
.B1(n_5587),
.B2(n_5586),
.C(n_602),
.Y(n_5593)
);

AOI22xp33_ASAP7_75t_SL g5594 ( 
.A1(n_5593),
.A2(n_5591),
.B1(n_600),
.B2(n_601),
.Y(n_5594)
);

AOI211xp5_ASAP7_75t_L g5595 ( 
.A1(n_5594),
.A2(n_598),
.B(n_603),
.C(n_606),
.Y(n_5595)
);


endmodule