module fake_netlist_5_821_n_1000 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1000);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1000;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_380;
wire n_419;
wire n_318;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_916;
wire n_452;
wire n_885;
wire n_397;
wire n_525;
wire n_493;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_998;
wire n_841;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_951;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_932;
wire n_417;
wire n_946;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_640;
wire n_275;
wire n_559;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_820;
wire n_757;
wire n_947;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_325;
wire n_449;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_271;
wire n_934;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_654;
wire n_370;
wire n_607;
wire n_976;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_783;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_670;
wire n_486;
wire n_816;
wire n_584;
wire n_681;
wire n_336;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_727;
wire n_553;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_517;
wire n_482;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_903;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_699;
wire n_632;
wire n_979;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_963;
wire n_745;
wire n_954;
wire n_627;
wire n_767;
wire n_206;
wire n_993;
wire n_217;
wire n_440;
wire n_726;
wire n_793;
wire n_478;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_970;
wire n_911;
wire n_557;
wire n_354;
wire n_575;
wire n_647;
wire n_480;
wire n_679;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_710;
wire n_707;
wire n_795;
wire n_832;
wire n_695;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_931;
wire n_870;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_666;
wire n_538;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_890;
wire n_960;
wire n_759;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_904;
wire n_985;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_401;
wire n_348;
wire n_626;
wire n_925;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_191),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_56),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_117),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_40),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_165),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_179),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_134),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_131),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_43),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_126),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_128),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_194),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_138),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_192),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_57),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_60),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_177),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_116),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_10),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_72),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_154),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_30),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_66),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_130),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_176),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_81),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_187),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_51),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_168),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_23),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_183),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_188),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_10),
.Y(n_229)
);

BUFx8_ASAP7_75t_SL g230 ( 
.A(n_59),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_148),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_45),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_53),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_190),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_65),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_122),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_14),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_193),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_129),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_100),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_106),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_28),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_62),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_47),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_71),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_76),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_92),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_114),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_149),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_82),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_87),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_19),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_147),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_68),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_36),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_112),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_22),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_105),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_4),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_46),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_41),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_74),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_96),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_163),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_77),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_182),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_73),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_78),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_67),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g270 ( 
.A(n_48),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_150),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_30),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_20),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_5),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_159),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_13),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_189),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_111),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_173),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_31),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_102),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_11),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_0),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_232),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_232),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_226),
.Y(n_286)
);

BUFx8_ASAP7_75t_SL g287 ( 
.A(n_230),
.Y(n_287)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_232),
.Y(n_288)
);

BUFx12f_ASAP7_75t_L g289 ( 
.A(n_282),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_226),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_196),
.B(n_0),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_232),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_1),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_237),
.Y(n_294)
);

AND2x4_ASAP7_75t_L g295 ( 
.A(n_246),
.B(n_38),
.Y(n_295)
);

AND2x4_ASAP7_75t_L g296 ( 
.A(n_246),
.B(n_248),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_226),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_212),
.B(n_1),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_248),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_209),
.B(n_2),
.Y(n_300)
);

NAND2xp33_ASAP7_75t_L g301 ( 
.A(n_226),
.B(n_2),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_206),
.Y(n_302)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_205),
.Y(n_303)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_205),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_272),
.B(n_242),
.Y(n_305)
);

AND2x4_ASAP7_75t_L g306 ( 
.A(n_206),
.B(n_39),
.Y(n_306)
);

AND2x4_ASAP7_75t_L g307 ( 
.A(n_221),
.B(n_42),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_257),
.Y(n_308)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_205),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_3),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_221),
.B(n_3),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_208),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_207),
.Y(n_313)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_207),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_257),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_207),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_257),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_257),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_211),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_214),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_216),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_229),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_239),
.Y(n_323)
);

AND2x6_ASAP7_75t_L g324 ( 
.A(n_241),
.B(n_44),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_244),
.B(n_49),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_255),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_234),
.B(n_4),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_250),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_273),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_276),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_268),
.B(n_5),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_258),
.B(n_6),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_274),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_280),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_260),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_261),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_294),
.B(n_210),
.Y(n_337)
);

OAI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_331),
.A2(n_217),
.B1(n_252),
.B2(n_265),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_223),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_333),
.B(n_227),
.Y(n_340)
);

AO22x2_ASAP7_75t_L g341 ( 
.A1(n_307),
.A2(n_266),
.B1(n_267),
.B2(n_282),
.Y(n_341)
);

OAI22xp33_ASAP7_75t_L g342 ( 
.A1(n_291),
.A2(n_259),
.B1(n_279),
.B2(n_200),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_334),
.B(n_282),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_305),
.B(n_195),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_305),
.B(n_197),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_297),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_300),
.B(n_198),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_327),
.A2(n_200),
.B1(n_279),
.B2(n_262),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_283),
.A2(n_262),
.B1(n_219),
.B2(n_259),
.Y(n_349)
);

OAI22xp33_ASAP7_75t_L g350 ( 
.A1(n_293),
.A2(n_281),
.B1(n_278),
.B2(n_277),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_313),
.B(n_199),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_329),
.A2(n_275),
.B1(n_271),
.B2(n_269),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_303),
.A2(n_264),
.B1(n_263),
.B2(n_256),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_313),
.B(n_201),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_329),
.A2(n_254),
.B1(n_253),
.B2(n_251),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_298),
.B(n_202),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_297),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_289),
.A2(n_203),
.B1(n_247),
.B2(n_245),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_316),
.B(n_204),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_285),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_316),
.B(n_213),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_289),
.A2(n_249),
.B1(n_243),
.B2(n_240),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_296),
.B(n_215),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_295),
.A2(n_238),
.B1(n_236),
.B2(n_235),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_308),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_296),
.B(n_218),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_296),
.B(n_220),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_308),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_295),
.A2(n_231),
.B1(n_228),
.B2(n_225),
.Y(n_369)
);

OAI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_303),
.A2(n_233),
.B1(n_224),
.B2(n_222),
.Y(n_370)
);

OA22x2_ASAP7_75t_L g371 ( 
.A1(n_296),
.A2(n_230),
.B1(n_7),
.B2(n_8),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_295),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_303),
.B(n_50),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_302),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_295),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_303),
.B(n_52),
.Y(n_376)
);

OAI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_303),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_377)
);

XNOR2x2_ASAP7_75t_SL g378 ( 
.A(n_310),
.B(n_14),
.Y(n_378)
);

OAI22xp33_ASAP7_75t_L g379 ( 
.A1(n_332),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_325),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_380)
);

OAI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_303),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_286),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_325),
.A2(n_18),
.B1(n_21),
.B2(n_22),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_302),
.Y(n_384)
);

AO22x2_ASAP7_75t_L g385 ( 
.A1(n_307),
.A2(n_306),
.B1(n_325),
.B2(n_310),
.Y(n_385)
);

BUFx6f_ASAP7_75t_SL g386 ( 
.A(n_287),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_304),
.B(n_21),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_302),
.Y(n_388)
);

OAI22xp33_ASAP7_75t_L g389 ( 
.A1(n_304),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_335),
.B(n_24),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_311),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_302),
.Y(n_392)
);

OR2x6_ASAP7_75t_L g393 ( 
.A(n_306),
.B(n_26),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_382),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_365),
.Y(n_395)
);

INVxp33_ASAP7_75t_L g396 ( 
.A(n_343),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_350),
.B(n_304),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_350),
.B(n_307),
.Y(n_398)
);

AO21x1_ASAP7_75t_L g399 ( 
.A1(n_387),
.A2(n_307),
.B(n_306),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_346),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_337),
.B(n_339),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_346),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_347),
.B(n_304),
.Y(n_403)
);

NOR2xp67_ASAP7_75t_L g404 ( 
.A(n_352),
.B(n_304),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_356),
.B(n_304),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_357),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_357),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_368),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_368),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_374),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_348),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_374),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_349),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_384),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_384),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_388),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_388),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_392),
.Y(n_418)
);

NAND2x1p5_ASAP7_75t_L g419 ( 
.A(n_387),
.B(n_299),
.Y(n_419)
);

AND2x2_ASAP7_75t_SL g420 ( 
.A(n_372),
.B(n_301),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_392),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_363),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_366),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_367),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_356),
.A2(n_324),
.B(n_335),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_360),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_360),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_358),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_360),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_362),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_347),
.B(n_309),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_378),
.B(n_54),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_340),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_344),
.B(n_309),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_355),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_385),
.A2(n_284),
.B(n_286),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_345),
.B(n_309),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_360),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_351),
.B(n_309),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_385),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_386),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_354),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_378),
.B(n_27),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_385),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_390),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_393),
.Y(n_446)
);

INVxp33_ASAP7_75t_SL g447 ( 
.A(n_364),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_393),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_393),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_373),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_359),
.B(n_361),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_369),
.B(n_338),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_341),
.B(n_309),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_380),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_376),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_383),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_342),
.B(n_28),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_375),
.Y(n_458)
);

INVxp33_ASAP7_75t_L g459 ( 
.A(n_341),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_391),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_341),
.B(n_309),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_377),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_381),
.Y(n_463)
);

AOI21x1_ASAP7_75t_L g464 ( 
.A1(n_371),
.A2(n_290),
.B(n_320),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_371),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_353),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_342),
.B(n_314),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_450),
.B(n_314),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_401),
.B(n_322),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_444),
.B(n_322),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_444),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_440),
.B(n_324),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_400),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_465),
.B(n_330),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_402),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_445),
.B(n_330),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_422),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_450),
.B(n_314),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_396),
.B(n_320),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_396),
.B(n_442),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_406),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_455),
.B(n_314),
.Y(n_482)
);

AND2x2_ASAP7_75t_SL g483 ( 
.A(n_397),
.B(n_324),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_419),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_464),
.B(n_324),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_423),
.B(n_314),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_407),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_419),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_455),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_447),
.B(n_370),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_424),
.B(n_314),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_442),
.B(n_299),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_425),
.A2(n_324),
.B(n_290),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_446),
.B(n_324),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_408),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_451),
.B(n_299),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g497 ( 
.A(n_433),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_448),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_462),
.B(n_299),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_463),
.B(n_299),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_467),
.B(n_302),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_441),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_398),
.B(n_453),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_409),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_398),
.B(n_315),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_461),
.B(n_315),
.Y(n_506)
);

AND2x6_ASAP7_75t_L g507 ( 
.A(n_466),
.B(n_324),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_412),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_449),
.B(n_55),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_458),
.B(n_315),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_394),
.B(n_58),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_412),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_460),
.B(n_318),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_454),
.B(n_318),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_399),
.B(n_312),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_403),
.B(n_431),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_447),
.B(n_389),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_395),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_410),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_433),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_420),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_397),
.B(n_389),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_436),
.A2(n_288),
.B(n_284),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_456),
.B(n_452),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_414),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_452),
.B(n_379),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_420),
.B(n_318),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_403),
.B(n_312),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_431),
.B(n_312),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_415),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_459),
.B(n_439),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_434),
.A2(n_288),
.B(n_284),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_426),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_434),
.B(n_312),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_413),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_437),
.B(n_312),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_459),
.B(n_317),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_416),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_417),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_418),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_437),
.B(n_319),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_404),
.B(n_317),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g543 ( 
.A(n_427),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_405),
.B(n_319),
.Y(n_544)
);

NAND2x1p5_ASAP7_75t_L g545 ( 
.A(n_421),
.B(n_317),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_429),
.Y(n_546)
);

AND2x6_ASAP7_75t_L g547 ( 
.A(n_438),
.B(n_285),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_435),
.B(n_379),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_457),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_435),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_428),
.B(n_61),
.Y(n_551)
);

INVxp67_ASAP7_75t_SL g552 ( 
.A(n_489),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_489),
.B(n_319),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_489),
.B(n_319),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_489),
.B(n_319),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_509),
.B(n_428),
.Y(n_556)
);

NAND2x1p5_ASAP7_75t_L g557 ( 
.A(n_471),
.B(n_285),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_503),
.B(n_443),
.Y(n_558)
);

NOR2x1_ASAP7_75t_R g559 ( 
.A(n_502),
.B(n_441),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_503),
.B(n_432),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_496),
.B(n_321),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_497),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_521),
.B(n_411),
.Y(n_563)
);

AND2x6_ASAP7_75t_L g564 ( 
.A(n_472),
.B(n_285),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_479),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_496),
.B(n_321),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_499),
.B(n_321),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_SL g568 ( 
.A(n_497),
.B(n_386),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_509),
.B(n_430),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_471),
.Y(n_570)
);

INVx4_ASAP7_75t_L g571 ( 
.A(n_471),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_499),
.B(n_321),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_521),
.B(n_411),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_479),
.B(n_430),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_522),
.B(n_29),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_524),
.B(n_321),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_512),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_471),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_512),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_471),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_520),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_512),
.Y(n_582)
);

OR2x6_ASAP7_75t_L g583 ( 
.A(n_551),
.B(n_323),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_509),
.B(n_63),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_509),
.B(n_64),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_500),
.B(n_323),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_508),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_508),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_477),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_470),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_525),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_527),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_535),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_527),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_511),
.B(n_69),
.Y(n_595)
);

BUFx12f_ASAP7_75t_L g596 ( 
.A(n_551),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_525),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_533),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_492),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_470),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_500),
.B(n_323),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_511),
.B(n_70),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_519),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_525),
.Y(n_604)
);

AND2x2_ASAP7_75t_SL g605 ( 
.A(n_483),
.B(n_323),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_539),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_501),
.B(n_323),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_519),
.Y(n_608)
);

NOR2x1_ASAP7_75t_L g609 ( 
.A(n_477),
.B(n_288),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_501),
.B(n_328),
.Y(n_610)
);

INVx6_ASAP7_75t_L g611 ( 
.A(n_511),
.Y(n_611)
);

NAND2x1p5_ASAP7_75t_L g612 ( 
.A(n_511),
.B(n_285),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_492),
.B(n_328),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_533),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_531),
.B(n_75),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_539),
.Y(n_616)
);

BUFx8_ASAP7_75t_L g617 ( 
.A(n_524),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_530),
.Y(n_618)
);

INVx3_ASAP7_75t_SL g619 ( 
.A(n_583),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_576),
.B(n_531),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_575),
.A2(n_526),
.B1(n_517),
.B2(n_548),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_591),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_591),
.Y(n_623)
);

CKINVDCx16_ASAP7_75t_R g624 ( 
.A(n_568),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_597),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_598),
.Y(n_626)
);

INVx4_ASAP7_75t_L g627 ( 
.A(n_578),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_598),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_597),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_598),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_617),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_578),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_565),
.B(n_469),
.Y(n_633)
);

INVx4_ASAP7_75t_L g634 ( 
.A(n_578),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_605),
.A2(n_483),
.B1(n_516),
.B2(n_488),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_578),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_617),
.Y(n_637)
);

BUFx5_ASAP7_75t_L g638 ( 
.A(n_605),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_589),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_562),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_617),
.Y(n_641)
);

CKINVDCx20_ASAP7_75t_R g642 ( 
.A(n_563),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_581),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_604),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_614),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_576),
.B(n_537),
.Y(n_646)
);

BUFx12f_ASAP7_75t_L g647 ( 
.A(n_596),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_571),
.Y(n_648)
);

INVxp67_ASAP7_75t_SL g649 ( 
.A(n_552),
.Y(n_649)
);

OAI22xp33_ASAP7_75t_L g650 ( 
.A1(n_583),
.A2(n_550),
.B1(n_477),
.B2(n_549),
.Y(n_650)
);

INVx1_ASAP7_75t_SL g651 ( 
.A(n_574),
.Y(n_651)
);

INVx3_ASAP7_75t_SL g652 ( 
.A(n_583),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_590),
.B(n_469),
.Y(n_653)
);

INVx5_ASAP7_75t_L g654 ( 
.A(n_614),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_604),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_606),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_614),
.Y(n_657)
);

INVx3_ASAP7_75t_SL g658 ( 
.A(n_556),
.Y(n_658)
);

INVx6_ASAP7_75t_L g659 ( 
.A(n_571),
.Y(n_659)
);

BUFx12f_ASAP7_75t_L g660 ( 
.A(n_596),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_592),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_614),
.Y(n_662)
);

BUFx4_ASAP7_75t_SL g663 ( 
.A(n_573),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_606),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_571),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_558),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_611),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_616),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_593),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_600),
.B(n_537),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_616),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_594),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_577),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_SL g674 ( 
.A1(n_651),
.A2(n_551),
.B1(n_575),
.B2(n_490),
.Y(n_674)
);

BUFx8_ASAP7_75t_L g675 ( 
.A(n_647),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_622),
.Y(n_676)
);

INVx6_ASAP7_75t_L g677 ( 
.A(n_647),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_642),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_629),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_622),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_621),
.A2(n_483),
.B1(n_551),
.B2(n_595),
.Y(n_681)
);

BUFx8_ASAP7_75t_L g682 ( 
.A(n_660),
.Y(n_682)
);

INVx6_ASAP7_75t_L g683 ( 
.A(n_660),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_620),
.A2(n_595),
.B1(n_602),
.B2(n_558),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_620),
.B(n_589),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_623),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_646),
.A2(n_602),
.B1(n_595),
.B2(n_505),
.Y(n_687)
);

INVx6_ASAP7_75t_L g688 ( 
.A(n_667),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_623),
.Y(n_689)
);

INVx4_ASAP7_75t_L g690 ( 
.A(n_654),
.Y(n_690)
);

BUFx10_ASAP7_75t_L g691 ( 
.A(n_669),
.Y(n_691)
);

OAI22xp33_ASAP7_75t_R g692 ( 
.A1(n_666),
.A2(n_549),
.B1(n_550),
.B2(n_498),
.Y(n_692)
);

HB1xp67_ASAP7_75t_L g693 ( 
.A(n_661),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_625),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_629),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_646),
.A2(n_602),
.B1(n_505),
.B2(n_615),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_625),
.Y(n_697)
);

OAI21xp33_ASAP7_75t_L g698 ( 
.A1(n_651),
.A2(n_550),
.B(n_560),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_670),
.A2(n_615),
.B1(n_618),
.B2(n_603),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_655),
.Y(n_700)
);

CKINVDCx11_ASAP7_75t_R g701 ( 
.A(n_624),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_644),
.Y(n_702)
);

INVx4_ASAP7_75t_SL g703 ( 
.A(n_619),
.Y(n_703)
);

BUFx4_ASAP7_75t_SL g704 ( 
.A(n_631),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_669),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_631),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_655),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_644),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_653),
.A2(n_615),
.B1(n_608),
.B2(n_513),
.Y(n_709)
);

BUFx4f_ASAP7_75t_L g710 ( 
.A(n_658),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_656),
.Y(n_711)
);

BUFx12f_ASAP7_75t_L g712 ( 
.A(n_637),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_656),
.Y(n_713)
);

BUFx2_ASAP7_75t_L g714 ( 
.A(n_661),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_643),
.A2(n_569),
.B1(n_556),
.B2(n_560),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_672),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_671),
.Y(n_717)
);

CKINVDCx11_ASAP7_75t_R g718 ( 
.A(n_624),
.Y(n_718)
);

OAI22xp33_ASAP7_75t_L g719 ( 
.A1(n_633),
.A2(n_611),
.B1(n_556),
.B2(n_569),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_SL g720 ( 
.A1(n_637),
.A2(n_569),
.B1(n_584),
.B2(n_585),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_650),
.A2(n_513),
.B1(n_585),
.B2(n_584),
.Y(n_721)
);

CKINVDCx11_ASAP7_75t_R g722 ( 
.A(n_640),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_671),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_635),
.A2(n_584),
.B1(n_585),
.B2(n_510),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_641),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_664),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_638),
.A2(n_510),
.B1(n_514),
.B2(n_599),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_681),
.A2(n_611),
.B1(n_619),
.B2(n_652),
.Y(n_728)
);

OAI21xp5_ASAP7_75t_SL g729 ( 
.A1(n_674),
.A2(n_681),
.B(n_720),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_721),
.A2(n_652),
.B1(n_619),
.B2(n_649),
.Y(n_730)
);

OAI222xp33_ASAP7_75t_L g731 ( 
.A1(n_684),
.A2(n_599),
.B1(n_480),
.B2(n_672),
.C1(n_498),
.C2(n_639),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_676),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_698),
.A2(n_658),
.B1(n_518),
.B2(n_514),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_692),
.A2(n_658),
.B1(n_641),
.B2(n_476),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_684),
.A2(n_476),
.B1(n_652),
.B2(n_506),
.Y(n_735)
);

INVx5_ASAP7_75t_SL g736 ( 
.A(n_704),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_721),
.A2(n_639),
.B1(n_488),
.B2(n_484),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_679),
.Y(n_738)
);

INVx5_ASAP7_75t_SL g739 ( 
.A(n_704),
.Y(n_739)
);

INVx4_ASAP7_75t_L g740 ( 
.A(n_710),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_680),
.Y(n_741)
);

OAI22xp33_ASAP7_75t_L g742 ( 
.A1(n_715),
.A2(n_667),
.B1(n_484),
.B2(n_518),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_719),
.A2(n_506),
.B1(n_486),
.B2(n_491),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_710),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_686),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_689),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_699),
.A2(n_612),
.B1(n_667),
.B2(n_659),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_719),
.A2(n_518),
.B1(n_507),
.B2(n_638),
.Y(n_748)
);

BUFx12f_ASAP7_75t_L g749 ( 
.A(n_722),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_709),
.A2(n_507),
.B1(n_638),
.B2(n_495),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_699),
.A2(n_612),
.B1(n_667),
.B2(n_659),
.Y(n_751)
);

OAI22xp5_ASAP7_75t_L g752 ( 
.A1(n_724),
.A2(n_696),
.B1(n_709),
.B2(n_687),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_694),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_724),
.A2(n_507),
.B1(n_638),
.B2(n_495),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_697),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_702),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_SL g757 ( 
.A1(n_678),
.A2(n_638),
.B1(n_659),
.B2(n_663),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_SL g758 ( 
.A1(n_677),
.A2(n_638),
.B1(n_659),
.B2(n_630),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_696),
.A2(n_507),
.B1(n_638),
.B2(n_481),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_SL g760 ( 
.A1(n_677),
.A2(n_638),
.B1(n_626),
.B2(n_628),
.Y(n_760)
);

INVx4_ASAP7_75t_L g761 ( 
.A(n_688),
.Y(n_761)
);

OAI222xp33_ASAP7_75t_L g762 ( 
.A1(n_687),
.A2(n_570),
.B1(n_601),
.B2(n_567),
.C1(n_572),
.C2(n_586),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_727),
.A2(n_507),
.B1(n_504),
.B2(n_473),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_691),
.Y(n_764)
);

BUFx5_ASAP7_75t_L g765 ( 
.A(n_708),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_L g766 ( 
.A1(n_727),
.A2(n_580),
.B1(n_542),
.B2(n_630),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_693),
.A2(n_580),
.B1(n_542),
.B2(n_630),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_695),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_693),
.A2(n_580),
.B1(n_628),
.B2(n_626),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_701),
.A2(n_507),
.B1(n_487),
.B2(n_504),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_718),
.A2(n_507),
.B1(n_473),
.B2(n_475),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_705),
.A2(n_481),
.B1(n_475),
.B2(n_487),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_685),
.A2(n_609),
.B1(n_491),
.B2(n_486),
.Y(n_773)
);

AOI211xp5_ASAP7_75t_SL g774 ( 
.A1(n_716),
.A2(n_530),
.B(n_610),
.C(n_607),
.Y(n_774)
);

OAI21xp5_ASAP7_75t_SL g775 ( 
.A1(n_714),
.A2(n_493),
.B(n_474),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_711),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_716),
.B(n_474),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_SL g778 ( 
.A1(n_677),
.A2(n_626),
.B1(n_628),
.B2(n_648),
.Y(n_778)
);

OAI222xp33_ASAP7_75t_L g779 ( 
.A1(n_713),
.A2(n_515),
.B1(n_588),
.B2(n_587),
.C1(n_668),
.C2(n_664),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_SL g780 ( 
.A1(n_683),
.A2(n_682),
.B1(n_675),
.B2(n_712),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_683),
.A2(n_538),
.B1(n_546),
.B2(n_588),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_706),
.Y(n_782)
);

BUFx8_ASAP7_75t_SL g783 ( 
.A(n_725),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_700),
.B(n_668),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_688),
.A2(n_654),
.B1(n_648),
.B2(n_665),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_703),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_683),
.A2(n_538),
.B1(n_546),
.B2(n_587),
.Y(n_787)
);

AOI221xp5_ASAP7_75t_L g788 ( 
.A1(n_752),
.A2(n_336),
.B1(n_328),
.B2(n_717),
.C(n_723),
.Y(n_788)
);

OAI221xp5_ASAP7_75t_L g789 ( 
.A1(n_729),
.A2(n_534),
.B1(n_536),
.B2(n_541),
.C(n_544),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_732),
.Y(n_790)
);

OAI22xp33_ASAP7_75t_L g791 ( 
.A1(n_734),
.A2(n_688),
.B1(n_665),
.B2(n_648),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_783),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_777),
.B(n_703),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_738),
.B(n_768),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_741),
.B(n_726),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_772),
.A2(n_654),
.B1(n_657),
.B2(n_665),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_745),
.B(n_707),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_735),
.A2(n_691),
.B1(n_682),
.B2(n_675),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_730),
.A2(n_538),
.B1(n_546),
.B2(n_613),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_735),
.A2(n_703),
.B1(n_539),
.B2(n_540),
.Y(n_800)
);

NAND3xp33_ASAP7_75t_L g801 ( 
.A(n_774),
.B(n_336),
.C(n_328),
.Y(n_801)
);

NAND3xp33_ASAP7_75t_L g802 ( 
.A(n_775),
.B(n_336),
.C(n_328),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_SL g803 ( 
.A1(n_728),
.A2(n_690),
.B1(n_665),
.B2(n_654),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_757),
.A2(n_743),
.B1(n_742),
.B2(n_780),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_746),
.B(n_673),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_SL g806 ( 
.A1(n_736),
.A2(n_690),
.B1(n_665),
.B2(n_654),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_733),
.A2(n_540),
.B1(n_561),
.B2(n_566),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_740),
.A2(n_540),
.B1(n_533),
.B2(n_494),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_SL g809 ( 
.A1(n_736),
.A2(n_654),
.B1(n_657),
.B2(n_662),
.Y(n_809)
);

NAND3xp33_ASAP7_75t_L g810 ( 
.A(n_770),
.B(n_336),
.C(n_529),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_740),
.A2(n_533),
.B1(n_494),
.B2(n_468),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_744),
.B(n_645),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_753),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_771),
.A2(n_657),
.B1(n_636),
.B2(n_634),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_744),
.B(n_645),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_755),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_743),
.A2(n_494),
.B1(n_657),
.B2(n_564),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_756),
.B(n_673),
.Y(n_818)
);

NAND2xp33_ASAP7_75t_L g819 ( 
.A(n_744),
.B(n_559),
.Y(n_819)
);

OA21x2_ASAP7_75t_L g820 ( 
.A1(n_762),
.A2(n_779),
.B(n_731),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_782),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_754),
.A2(n_636),
.B1(n_634),
.B2(n_632),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_750),
.A2(n_336),
.B1(n_532),
.B2(n_579),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_776),
.B(n_662),
.Y(n_824)
);

AOI221xp5_ASAP7_75t_L g825 ( 
.A1(n_737),
.A2(n_528),
.B1(n_543),
.B2(n_494),
.C(n_482),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_SL g826 ( 
.A1(n_739),
.A2(n_747),
.B1(n_751),
.B2(n_786),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_749),
.A2(n_577),
.B1(n_579),
.B2(n_582),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_748),
.A2(n_582),
.B1(n_554),
.B2(n_555),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_784),
.B(n_645),
.Y(n_829)
);

OAI222xp33_ASAP7_75t_L g830 ( 
.A1(n_758),
.A2(n_634),
.B1(n_627),
.B2(n_632),
.C1(n_557),
.C2(n_553),
.Y(n_830)
);

OAI21xp5_ASAP7_75t_SL g831 ( 
.A1(n_760),
.A2(n_472),
.B(n_485),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_759),
.A2(n_627),
.B1(n_634),
.B2(n_632),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_773),
.A2(n_632),
.B1(n_627),
.B2(n_472),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_SL g834 ( 
.A1(n_739),
.A2(n_645),
.B1(n_662),
.B2(n_627),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_763),
.A2(n_472),
.B1(n_645),
.B2(n_662),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_790),
.B(n_765),
.Y(n_836)
);

NAND3xp33_ASAP7_75t_L g837 ( 
.A(n_798),
.B(n_826),
.C(n_804),
.Y(n_837)
);

NOR3xp33_ASAP7_75t_L g838 ( 
.A(n_802),
.B(n_764),
.C(n_761),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_813),
.B(n_765),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_816),
.B(n_765),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_794),
.B(n_765),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_800),
.A2(n_781),
.B1(n_787),
.B2(n_778),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_795),
.B(n_765),
.Y(n_843)
);

NAND3xp33_ASAP7_75t_L g844 ( 
.A(n_788),
.B(n_827),
.C(n_801),
.Y(n_844)
);

NAND2xp33_ASAP7_75t_SL g845 ( 
.A(n_792),
.B(n_761),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_830),
.A2(n_785),
.B(n_766),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_805),
.B(n_797),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_821),
.B(n_769),
.Y(n_848)
);

NAND3xp33_ASAP7_75t_L g849 ( 
.A(n_827),
.B(n_767),
.C(n_533),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_824),
.B(n_29),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_818),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_829),
.B(n_31),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_793),
.B(n_32),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_820),
.B(n_32),
.Y(n_854)
);

OA21x2_ASAP7_75t_L g855 ( 
.A1(n_831),
.A2(n_810),
.B(n_817),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_803),
.A2(n_791),
.B1(n_820),
.B2(n_833),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_820),
.B(n_828),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_833),
.B(n_33),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_812),
.B(n_33),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_815),
.B(n_828),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_834),
.B(n_34),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_835),
.B(n_34),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_SL g863 ( 
.A1(n_796),
.A2(n_662),
.B1(n_564),
.B2(n_485),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_835),
.B(n_35),
.Y(n_864)
);

OAI21xp33_ASAP7_75t_L g865 ( 
.A1(n_819),
.A2(n_35),
.B(n_36),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_806),
.B(n_37),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_832),
.B(n_37),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_799),
.B(n_79),
.Y(n_868)
);

NAND2x1p5_ASAP7_75t_L g869 ( 
.A(n_809),
.B(n_485),
.Y(n_869)
);

OAI221xp5_ASAP7_75t_L g870 ( 
.A1(n_811),
.A2(n_478),
.B1(n_557),
.B2(n_523),
.C(n_545),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_832),
.B(n_292),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_837),
.B(n_789),
.Y(n_872)
);

NOR3xp33_ASAP7_75t_L g873 ( 
.A(n_865),
.B(n_814),
.C(n_822),
.Y(n_873)
);

AO21x2_ASAP7_75t_L g874 ( 
.A1(n_838),
.A2(n_485),
.B(n_823),
.Y(n_874)
);

NAND3xp33_ASAP7_75t_L g875 ( 
.A(n_865),
.B(n_808),
.C(n_825),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_847),
.B(n_807),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_839),
.B(n_823),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_851),
.B(n_80),
.Y(n_878)
);

OA211x2_ASAP7_75t_L g879 ( 
.A1(n_866),
.A2(n_83),
.B(n_84),
.C(n_85),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_839),
.B(n_840),
.Y(n_880)
);

NAND3xp33_ASAP7_75t_L g881 ( 
.A(n_854),
.B(n_292),
.C(n_284),
.Y(n_881)
);

INVx1_ASAP7_75t_SL g882 ( 
.A(n_845),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_836),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_840),
.B(n_86),
.Y(n_884)
);

NAND3xp33_ASAP7_75t_L g885 ( 
.A(n_854),
.B(n_852),
.C(n_858),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_843),
.B(n_292),
.Y(n_886)
);

AO21x2_ASAP7_75t_L g887 ( 
.A1(n_857),
.A2(n_564),
.B(n_89),
.Y(n_887)
);

NAND3xp33_ASAP7_75t_L g888 ( 
.A(n_860),
.B(n_292),
.C(n_284),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_845),
.A2(n_842),
.B1(n_855),
.B2(n_867),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_853),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_855),
.A2(n_564),
.B1(n_545),
.B2(n_547),
.Y(n_891)
);

AO21x2_ASAP7_75t_L g892 ( 
.A1(n_857),
.A2(n_564),
.B(n_90),
.Y(n_892)
);

NAND3xp33_ASAP7_75t_L g893 ( 
.A(n_862),
.B(n_292),
.C(n_284),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_867),
.A2(n_545),
.B1(n_547),
.B2(n_93),
.Y(n_894)
);

XOR2x2_ASAP7_75t_L g895 ( 
.A(n_872),
.B(n_861),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_883),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_880),
.Y(n_897)
);

NOR4xp25_ASAP7_75t_L g898 ( 
.A(n_872),
.B(n_864),
.C(n_859),
.D(n_850),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_873),
.A2(n_856),
.B1(n_855),
.B2(n_844),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_886),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_877),
.B(n_850),
.Y(n_901)
);

NOR4xp25_ASAP7_75t_L g902 ( 
.A(n_885),
.B(n_848),
.C(n_849),
.D(n_868),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_877),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_887),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_876),
.Y(n_905)
);

INVxp67_ASAP7_75t_SL g906 ( 
.A(n_889),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_884),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_884),
.B(n_851),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_878),
.Y(n_909)
);

XNOR2xp5_ASAP7_75t_L g910 ( 
.A(n_890),
.B(n_869),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_903),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_896),
.Y(n_912)
);

AO22x2_ASAP7_75t_L g913 ( 
.A1(n_906),
.A2(n_882),
.B1(n_875),
.B2(n_881),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_901),
.Y(n_914)
);

INVx1_ASAP7_75t_SL g915 ( 
.A(n_901),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_900),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_900),
.Y(n_917)
);

INVx1_ASAP7_75t_SL g918 ( 
.A(n_908),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_905),
.Y(n_919)
);

OA22x2_ASAP7_75t_L g920 ( 
.A1(n_914),
.A2(n_899),
.B1(n_910),
.B2(n_905),
.Y(n_920)
);

XNOR2xp5_ASAP7_75t_L g921 ( 
.A(n_915),
.B(n_895),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_918),
.B(n_890),
.Y(n_922)
);

AOI22x1_ASAP7_75t_L g923 ( 
.A1(n_913),
.A2(n_910),
.B1(n_904),
.B2(n_909),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_912),
.Y(n_924)
);

XNOR2x1_ASAP7_75t_L g925 ( 
.A(n_913),
.B(n_895),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_913),
.A2(n_898),
.B1(n_902),
.B2(n_919),
.Y(n_926)
);

OAI22xp33_ASAP7_75t_SL g927 ( 
.A1(n_911),
.A2(n_904),
.B1(n_907),
.B2(n_897),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_924),
.Y(n_928)
);

AOI322xp5_ASAP7_75t_L g929 ( 
.A1(n_926),
.A2(n_911),
.A3(n_917),
.B1(n_916),
.B2(n_894),
.C1(n_891),
.C2(n_871),
.Y(n_929)
);

INVxp67_ASAP7_75t_SL g930 ( 
.A(n_925),
.Y(n_930)
);

AO22x2_ASAP7_75t_L g931 ( 
.A1(n_923),
.A2(n_916),
.B1(n_888),
.B2(n_893),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_921),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_930),
.A2(n_920),
.B1(n_922),
.B2(n_927),
.Y(n_933)
);

AND4x1_ASAP7_75t_L g934 ( 
.A(n_932),
.B(n_929),
.C(n_931),
.D(n_894),
.Y(n_934)
);

AO22x2_ASAP7_75t_L g935 ( 
.A1(n_928),
.A2(n_846),
.B1(n_841),
.B2(n_871),
.Y(n_935)
);

CKINVDCx20_ASAP7_75t_R g936 ( 
.A(n_933),
.Y(n_936)
);

OAI22x1_ASAP7_75t_L g937 ( 
.A1(n_934),
.A2(n_929),
.B1(n_931),
.B2(n_869),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_935),
.A2(n_879),
.B1(n_869),
.B2(n_863),
.Y(n_938)
);

OAI22xp33_ASAP7_75t_L g939 ( 
.A1(n_933),
.A2(n_892),
.B1(n_887),
.B2(n_874),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_936),
.B(n_892),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_937),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_938),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_939),
.Y(n_943)
);

AOI22xp33_ASAP7_75t_SL g944 ( 
.A1(n_936),
.A2(n_874),
.B1(n_870),
.B2(n_94),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_936),
.B(n_88),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_936),
.B(n_91),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_941),
.B(n_95),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_942),
.A2(n_943),
.B1(n_940),
.B2(n_946),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_945),
.B(n_97),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_944),
.Y(n_950)
);

OAI22xp33_ASAP7_75t_L g951 ( 
.A1(n_941),
.A2(n_98),
.B1(n_99),
.B2(n_101),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_941),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_941),
.A2(n_547),
.B1(n_104),
.B2(n_107),
.Y(n_953)
);

NOR4xp25_ASAP7_75t_L g954 ( 
.A(n_952),
.B(n_103),
.C(n_108),
.D(n_109),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_948),
.A2(n_547),
.B1(n_115),
.B2(n_118),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_950),
.A2(n_547),
.B1(n_119),
.B2(n_120),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_947),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_951),
.A2(n_547),
.B1(n_121),
.B2(n_123),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_949),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_953),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_959),
.B(n_110),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_957),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_960),
.Y(n_963)
);

OR2x2_ASAP7_75t_L g964 ( 
.A(n_954),
.B(n_124),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_958),
.Y(n_965)
);

AO22x2_ASAP7_75t_L g966 ( 
.A1(n_955),
.A2(n_956),
.B1(n_127),
.B2(n_132),
.Y(n_966)
);

INVxp67_ASAP7_75t_SL g967 ( 
.A(n_959),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_957),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_957),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_957),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_963),
.A2(n_125),
.B1(n_133),
.B2(n_135),
.Y(n_971)
);

AO22x2_ASAP7_75t_L g972 ( 
.A1(n_967),
.A2(n_964),
.B1(n_969),
.B2(n_968),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_970),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_967),
.A2(n_547),
.B1(n_137),
.B2(n_139),
.Y(n_974)
);

AO22x2_ASAP7_75t_L g975 ( 
.A1(n_962),
.A2(n_136),
.B1(n_140),
.B2(n_141),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_SL g976 ( 
.A1(n_970),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_965),
.A2(n_145),
.B1(n_146),
.B2(n_151),
.Y(n_977)
);

AOI22xp5_ASAP7_75t_L g978 ( 
.A1(n_961),
.A2(n_152),
.B1(n_153),
.B2(n_155),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_966),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_966),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_966),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_973),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_972),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_980),
.Y(n_984)
);

INVxp33_ASAP7_75t_SL g985 ( 
.A(n_976),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_975),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_979),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_981),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_L g989 ( 
.A1(n_985),
.A2(n_971),
.B1(n_974),
.B2(n_977),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_982),
.A2(n_978),
.B1(n_166),
.B2(n_167),
.Y(n_990)
);

AOI22xp33_ASAP7_75t_L g991 ( 
.A1(n_983),
.A2(n_164),
.B1(n_169),
.B2(n_170),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_989),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_990),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_SL g994 ( 
.A1(n_992),
.A2(n_984),
.B1(n_986),
.B2(n_987),
.Y(n_994)
);

AO22x2_ASAP7_75t_L g995 ( 
.A1(n_993),
.A2(n_988),
.B1(n_991),
.B2(n_174),
.Y(n_995)
);

OA22x2_ASAP7_75t_L g996 ( 
.A1(n_992),
.A2(n_171),
.B1(n_172),
.B2(n_175),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_994),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_995),
.Y(n_998)
);

AOI221xp5_ASAP7_75t_L g999 ( 
.A1(n_997),
.A2(n_996),
.B1(n_178),
.B2(n_180),
.C(n_181),
.Y(n_999)
);

AOI211xp5_ASAP7_75t_L g1000 ( 
.A1(n_999),
.A2(n_998),
.B(n_184),
.C(n_185),
.Y(n_1000)
);


endmodule