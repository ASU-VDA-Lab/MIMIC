module fake_jpeg_11230_n_116 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_116);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_116;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_22),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_25),
.B(n_17),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_53),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_47),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_3),
.Y(n_65)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_49),
.B(n_1),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_58),
.B(n_44),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_2),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_42),
.Y(n_67)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_55),
.C(n_51),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_7),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_7),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_SL g66 ( 
.A1(n_59),
.A2(n_48),
.B(n_42),
.C(n_47),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_70),
.B(n_6),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_5),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_69),
.B(n_3),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_40),
.B1(n_46),
.B2(n_48),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_40),
.B1(n_38),
.B2(n_41),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_73),
.A2(n_47),
.B1(n_24),
.B2(n_26),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_81),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_76),
.B(n_78),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_4),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_86),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_4),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_62),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_82),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_5),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_28),
.B(n_29),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_14),
.Y(n_93)
);

BUFx24_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_88),
.Y(n_101)
);

AOI32xp33_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_13),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_93),
.B(n_94),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_70),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_86),
.A2(n_20),
.B1(n_21),
.B2(n_27),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_37),
.B1(n_98),
.B2(n_101),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_74),
.B(n_33),
.Y(n_102)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_31),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_100),
.B(n_32),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_104),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_74),
.B(n_35),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_89),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_106),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_96),
.B(n_90),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_110),
.Y(n_113)
);

BUFx24_ASAP7_75t_SL g114 ( 
.A(n_113),
.Y(n_114)
);

AOI322xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_108),
.A3(n_109),
.B1(n_105),
.B2(n_92),
.C1(n_103),
.C2(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_115),
.B(n_91),
.Y(n_116)
);


endmodule