module fake_jpeg_24033_n_220 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_220);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_220;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_25),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_25),
.Y(n_68)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_25),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_17),
.B(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_44),
.Y(n_46)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_48),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_49),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_26),
.B1(n_25),
.B2(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_52),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_26),
.B1(n_33),
.B2(n_30),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_33),
.B1(n_32),
.B2(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_58),
.Y(n_76)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_64),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_18),
.B1(n_31),
.B2(n_22),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_66),
.Y(n_78)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_18),
.B1(n_31),
.B2(n_22),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_45),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_36),
.A2(n_32),
.B1(n_29),
.B2(n_27),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_27),
.B(n_29),
.C(n_20),
.Y(n_100)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_86),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_82),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_45),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_65),
.B(n_43),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_83),
.B(n_97),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_65),
.B(n_43),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_84),
.B(n_87),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_42),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_92),
.Y(n_114)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_46),
.B(n_16),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_19),
.Y(n_89)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_42),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

BUFx16f_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_46),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_96),
.B(n_99),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_62),
.B(n_19),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_69),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_100),
.A2(n_16),
.B(n_23),
.Y(n_120)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_41),
.B1(n_34),
.B2(n_39),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_103),
.A2(n_123),
.B1(n_124),
.B2(n_127),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_51),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_121),
.C(n_88),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_78),
.A2(n_34),
.B1(n_39),
.B2(n_47),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_116),
.B1(n_117),
.B2(n_122),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_20),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_110),
.B(n_120),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_59),
.B1(n_67),
.B2(n_58),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_99),
.A2(n_55),
.B1(n_37),
.B2(n_35),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_82),
.B(n_37),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_92),
.A2(n_37),
.B1(n_57),
.B2(n_24),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_85),
.A2(n_37),
.B1(n_24),
.B2(n_23),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_96),
.A2(n_15),
.B1(n_14),
.B2(n_2),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_79),
.B(n_77),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_97),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_75),
.A2(n_15),
.B1(n_1),
.B2(n_3),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_75),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_128),
.A2(n_81),
.B1(n_91),
.B2(n_71),
.Y(n_140)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_131),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_81),
.B(n_91),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_132),
.B(n_133),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_115),
.A2(n_93),
.B1(n_80),
.B2(n_86),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_115),
.A2(n_101),
.B1(n_95),
.B2(n_94),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_98),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_134),
.A2(n_146),
.B(n_119),
.Y(n_167)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_136),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_83),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_142),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_103),
.A2(n_114),
.B1(n_121),
.B2(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_72),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_149),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_121),
.B(n_122),
.Y(n_146)
);

NOR3xp33_ASAP7_75t_SL g147 ( 
.A(n_107),
.B(n_90),
.C(n_4),
.Y(n_147)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_106),
.C(n_124),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_117),
.Y(n_148)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

AOI322xp5_ASAP7_75t_L g151 ( 
.A1(n_134),
.A2(n_137),
.A3(n_139),
.B1(n_150),
.B2(n_142),
.C1(n_149),
.C2(n_146),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_167),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_156),
.Y(n_176)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_126),
.C(n_106),
.Y(n_156)
);

A2O1A1O1Ixp25_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_144),
.B(n_130),
.C(n_145),
.D(n_141),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_161),
.B(n_138),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_165),
.B(n_4),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_166),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_165),
.A2(n_141),
.B1(n_137),
.B2(n_132),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_169),
.B1(n_173),
.B2(n_174),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_138),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_161),
.C(n_154),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_162),
.A2(n_143),
.B(n_118),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_160),
.A2(n_147),
.B1(n_110),
.B2(n_128),
.Y(n_172)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

OA22x2_ASAP7_75t_L g173 ( 
.A1(n_162),
.A2(n_127),
.B1(n_111),
.B2(n_118),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_119),
.B1(n_111),
.B2(n_125),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_158),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_177)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_177),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_157),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_125),
.B(n_7),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_166),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_190),
.Y(n_197)
);

FAx1_ASAP7_75t_SL g184 ( 
.A(n_170),
.B(n_155),
.CI(n_164),
.CON(n_184),
.SN(n_184)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_184),
.B(n_186),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_153),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_189),
.B(n_172),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_179),
.B(n_159),
.Y(n_191)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_155),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_181),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_200),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_182),
.A2(n_154),
.B1(n_173),
.B2(n_171),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_194),
.A2(n_199),
.B1(n_187),
.B2(n_185),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_L g195 ( 
.A1(n_182),
.A2(n_180),
.B(n_159),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_198),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_188),
.A2(n_173),
.B1(n_177),
.B2(n_175),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_202),
.B(n_207),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_183),
.C(n_190),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_205),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_184),
.C(n_192),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_195),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_194),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_210),
.Y(n_213)
);

AOI322xp5_ASAP7_75t_L g210 ( 
.A1(n_206),
.A2(n_201),
.A3(n_203),
.B1(n_189),
.B2(n_205),
.C1(n_6),
.C2(n_10),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_211),
.A2(n_6),
.B(n_8),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_208),
.A2(n_8),
.B(n_9),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_214),
.A2(n_9),
.B(n_10),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_215),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_217),
.A2(n_218),
.B(n_12),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_215),
.A2(n_213),
.B(n_209),
.Y(n_218)
);

BUFx24_ASAP7_75t_SL g220 ( 
.A(n_219),
.Y(n_220)
);


endmodule