module fake_netlist_5_1586_n_5372 (n_924, n_977, n_611, n_1126, n_1166, n_469, n_82, n_785, n_549, n_532, n_1161, n_1150, n_226, n_667, n_790, n_1055, n_111, n_880, n_544, n_1007, n_155, n_552, n_1198, n_1099, n_956, n_564, n_423, n_21, n_105, n_1021, n_4, n_551, n_688, n_800, n_671, n_819, n_1022, n_915, n_864, n_173, n_859, n_951, n_447, n_247, n_292, n_625, n_854, n_674, n_417, n_516, n_933, n_1152, n_497, n_606, n_275, n_26, n_877, n_2, n_755, n_1118, n_6, n_947, n_373, n_307, n_530, n_87, n_150, n_1107, n_556, n_1230, n_668, n_375, n_301, n_929, n_1124, n_902, n_191, n_1104, n_659, n_51, n_171, n_1182, n_579, n_938, n_1098, n_320, n_1154, n_1242, n_1135, n_24, n_406, n_519, n_1016, n_1243, n_546, n_101, n_281, n_240, n_291, n_231, n_257, n_731, n_371, n_709, n_317, n_1236, n_569, n_227, n_920, n_94, n_335, n_370, n_976, n_343, n_308, n_297, n_156, n_1078, n_775, n_219, n_157, n_600, n_223, n_264, n_955, n_163, n_339, n_1146, n_882, n_183, n_243, n_1036, n_1097, n_347, n_59, n_550, n_696, n_897, n_215, n_350, n_196, n_798, n_646, n_436, n_1216, n_290, n_580, n_1040, n_578, n_926, n_344, n_1218, n_422, n_475, n_777, n_1070, n_1030, n_72, n_415, n_1071, n_485, n_1165, n_496, n_958, n_1034, n_670, n_48, n_521, n_663, n_845, n_673, n_837, n_1239, n_528, n_680, n_395, n_164, n_553, n_901, n_813, n_214, n_675, n_888, n_1167, n_637, n_184, n_446, n_1064, n_144, n_858, n_114, n_96, n_923, n_691, n_1151, n_881, n_468, n_213, n_129, n_342, n_464, n_363, n_197, n_1069, n_1075, n_460, n_889, n_973, n_477, n_571, n_461, n_1211, n_1197, n_907, n_190, n_989, n_1039, n_34, n_228, n_283, n_488, n_736, n_892, n_1000, n_1202, n_1002, n_49, n_310, n_54, n_593, n_12, n_748, n_586, n_1058, n_838, n_332, n_1053, n_1224, n_349, n_1248, n_230, n_953, n_279, n_1014, n_1241, n_70, n_289, n_963, n_1052, n_954, n_627, n_440, n_793, n_478, n_476, n_534, n_884, n_345, n_944, n_91, n_182, n_143, n_647, n_237, n_407, n_1072, n_832, n_857, n_207, n_561, n_18, n_1027, n_971, n_1156, n_117, n_326, n_794, n_404, n_686, n_847, n_596, n_558, n_702, n_822, n_728, n_266, n_1162, n_272, n_1199, n_352, n_53, n_1038, n_520, n_409, n_887, n_154, n_71, n_300, n_809, n_870, n_931, n_599, n_434, n_868, n_639, n_914, n_411, n_414, n_965, n_935, n_121, n_1175, n_817, n_360, n_36, n_64, n_759, n_28, n_806, n_324, n_187, n_1189, n_103, n_97, n_11, n_7, n_706, n_746, n_747, n_52, n_784, n_110, n_1244, n_431, n_1194, n_615, n_851, n_843, n_523, n_913, n_705, n_865, n_61, n_678, n_697, n_127, n_1222, n_75, n_776, n_367, n_452, n_525, n_649, n_547, n_43, n_1191, n_116, n_284, n_1128, n_139, n_744, n_590, n_629, n_254, n_1233, n_23, n_526, n_293, n_372, n_677, n_244, n_47, n_1121, n_314, n_368, n_433, n_604, n_8, n_949, n_100, n_1008, n_946, n_1001, n_498, n_689, n_738, n_640, n_252, n_624, n_295, n_133, n_1010, n_1231, n_739, n_1195, n_610, n_936, n_568, n_39, n_1090, n_757, n_633, n_439, n_106, n_259, n_448, n_758, n_999, n_93, n_1158, n_563, n_1145, n_878, n_524, n_204, n_394, n_1049, n_1153, n_741, n_1068, n_122, n_331, n_10, n_906, n_1163, n_1207, n_919, n_908, n_90, n_724, n_658, n_456, n_959, n_535, n_152, n_940, n_9, n_592, n_1169, n_45, n_1017, n_123, n_978, n_1054, n_1095, n_267, n_514, n_457, n_1079, n_1045, n_1208, n_603, n_484, n_1033, n_442, n_131, n_636, n_660, n_1009, n_1148, n_109, n_742, n_750, n_995, n_454, n_374, n_185, n_396, n_1073, n_255, n_662, n_459, n_218, n_962, n_1215, n_1171, n_723, n_1065, n_473, n_1043, n_355, n_486, n_614, n_337, n_88, n_1177, n_168, n_974, n_727, n_1159, n_957, n_773, n_208, n_142, n_743, n_299, n_303, n_296, n_613, n_1119, n_1240, n_65, n_829, n_361, n_700, n_1237, n_573, n_69, n_1132, n_388, n_1127, n_761, n_1006, n_329, n_274, n_582, n_73, n_19, n_309, n_30, n_512, n_84, n_130, n_322, n_652, n_1111, n_25, n_1093, n_288, n_1031, n_263, n_609, n_1041, n_44, n_224, n_383, n_834, n_112, n_765, n_893, n_1015, n_1140, n_891, n_239, n_630, n_55, n_504, n_511, n_874, n_358, n_1101, n_77, n_102, n_1106, n_987, n_261, n_174, n_767, n_993, n_545, n_441, n_860, n_450, n_429, n_948, n_1217, n_628, n_365, n_729, n_1131, n_1084, n_970, n_911, n_83, n_513, n_1094, n_560, n_340, n_1044, n_1205, n_346, n_1209, n_495, n_602, n_574, n_879, n_16, n_58, n_623, n_405, n_824, n_359, n_490, n_996, n_921, n_233, n_572, n_366, n_815, n_128, n_120, n_327, n_135, n_1037, n_1080, n_426, n_1082, n_589, n_716, n_562, n_62, n_952, n_1229, n_391, n_701, n_1023, n_645, n_539, n_803, n_1092, n_238, n_531, n_890, n_764, n_1056, n_162, n_960, n_222, n_1123, n_1047, n_634, n_199, n_32, n_348, n_1029, n_925, n_1206, n_424, n_256, n_950, n_380, n_419, n_444, n_1060, n_1141, n_316, n_389, n_418, n_248, n_136, n_86, n_146, n_912, n_315, n_968, n_451, n_619, n_408, n_376, n_967, n_74, n_1139, n_515, n_57, n_351, n_885, n_397, n_483, n_683, n_1057, n_1051, n_1085, n_1066, n_721, n_1157, n_841, n_1050, n_22, n_802, n_46, n_983, n_38, n_280, n_873, n_378, n_1112, n_762, n_17, n_690, n_33, n_583, n_302, n_1203, n_821, n_321, n_1179, n_621, n_753, n_455, n_1048, n_212, n_385, n_507, n_330, n_1228, n_972, n_692, n_820, n_1200, n_1185, n_991, n_828, n_779, n_576, n_1143, n_804, n_537, n_945, n_492, n_153, n_943, n_341, n_250, n_992, n_543, n_260, n_842, n_650, n_984, n_694, n_286, n_883, n_470, n_325, n_449, n_132, n_1214, n_900, n_856, n_918, n_942, n_189, n_1147, n_13, n_1077, n_540, n_618, n_896, n_323, n_195, n_356, n_894, n_831, n_964, n_1096, n_234, n_833, n_5, n_225, n_988, n_814, n_192, n_1201, n_1114, n_655, n_669, n_472, n_1176, n_387, n_1149, n_398, n_635, n_763, n_1020, n_1062, n_211, n_1219, n_3, n_1204, n_178, n_1035, n_287, n_555, n_783, n_1188, n_661, n_41, n_849, n_15, n_336, n_584, n_681, n_50, n_430, n_510, n_216, n_311, n_830, n_801, n_241, n_875, n_357, n_1110, n_445, n_749, n_1134, n_717, n_165, n_939, n_482, n_1088, n_588, n_1173, n_789, n_1232, n_734, n_638, n_866, n_107, n_969, n_1019, n_1105, n_249, n_304, n_577, n_338, n_149, n_693, n_14, n_836, n_990, n_975, n_567, n_778, n_1122, n_151, n_306, n_458, n_770, n_1102, n_711, n_85, n_1187, n_1164, n_489, n_1174, n_617, n_876, n_1190, n_118, n_601, n_917, n_966, n_253, n_1116, n_1212, n_172, n_206, n_217, n_726, n_982, n_818, n_861, n_1183, n_899, n_210, n_774, n_1059, n_176, n_1133, n_557, n_1005, n_607, n_1003, n_679, n_710, n_527, n_1168, n_707, n_937, n_393, n_108, n_487, n_665, n_66, n_177, n_421, n_910, n_768, n_205, n_1136, n_754, n_179, n_1125, n_125, n_410, n_708, n_529, n_735, n_232, n_1109, n_126, n_895, n_202, n_427, n_791, n_732, n_193, n_808, n_797, n_1025, n_500, n_1067, n_148, n_435, n_159, n_766, n_541, n_538, n_1117, n_799, n_687, n_715, n_1213, n_536, n_872, n_594, n_200, n_1155, n_89, n_115, n_1011, n_1184, n_985, n_869, n_810, n_416, n_827, n_401, n_626, n_1144, n_1137, n_1170, n_305, n_137, n_676, n_294, n_318, n_653, n_642, n_194, n_855, n_1178, n_850, n_684, n_124, n_268, n_664, n_503, n_235, n_605, n_353, n_620, n_643, n_916, n_1081, n_493, n_1235, n_703, n_698, n_980, n_1115, n_780, n_998, n_467, n_1227, n_840, n_501, n_823, n_245, n_725, n_672, n_581, n_382, n_554, n_898, n_1013, n_718, n_265, n_1120, n_719, n_443, n_198, n_714, n_909, n_997, n_932, n_612, n_788, n_119, n_559, n_825, n_508, n_506, n_737, n_986, n_509, n_147, n_67, n_1192, n_1024, n_1063, n_209, n_733, n_941, n_981, n_68, n_867, n_186, n_134, n_587, n_63, n_792, n_756, n_399, n_1238, n_548, n_812, n_298, n_518, n_505, n_282, n_752, n_905, n_1108, n_782, n_1100, n_862, n_760, n_381, n_220, n_390, n_31, n_481, n_769, n_42, n_1046, n_271, n_934, n_826, n_886, n_1221, n_654, n_1172, n_167, n_379, n_428, n_570, n_853, n_377, n_751, n_786, n_1083, n_1142, n_1129, n_392, n_158, n_704, n_787, n_138, n_961, n_771, n_276, n_95, n_1225, n_169, n_522, n_400, n_930, n_181, n_221, n_622, n_1087, n_386, n_994, n_848, n_1223, n_104, n_682, n_56, n_141, n_1247, n_922, n_816, n_591, n_145, n_313, n_631, n_479, n_1246, n_432, n_839, n_1210, n_328, n_140, n_369, n_871, n_598, n_685, n_928, n_608, n_78, n_772, n_499, n_517, n_98, n_402, n_413, n_1086, n_796, n_236, n_1012, n_1, n_903, n_740, n_203, n_384, n_80, n_35, n_277, n_1061, n_92, n_333, n_462, n_1193, n_258, n_1113, n_29, n_79, n_1226, n_722, n_188, n_844, n_201, n_471, n_852, n_40, n_1028, n_781, n_474, n_542, n_463, n_595, n_502, n_466, n_420, n_632, n_699, n_979, n_1245, n_846, n_465, n_76, n_362, n_170, n_27, n_161, n_273, n_585, n_270, n_616, n_81, n_745, n_1103, n_648, n_312, n_1076, n_1091, n_494, n_641, n_730, n_354, n_575, n_480, n_425, n_795, n_695, n_180, n_656, n_1220, n_37, n_229, n_437, n_60, n_403, n_453, n_1130, n_720, n_0, n_863, n_805, n_113, n_712, n_246, n_1042, n_269, n_285, n_412, n_657, n_644, n_1160, n_491, n_1074, n_251, n_160, n_566, n_565, n_597, n_1181, n_1196, n_651, n_334, n_811, n_807, n_835, n_175, n_666, n_262, n_99, n_1026, n_1234, n_319, n_364, n_1138, n_927, n_20, n_1089, n_1004, n_1186, n_1032, n_242, n_1018, n_438, n_713, n_904, n_166, n_1180, n_533, n_278, n_5372);

input n_924;
input n_977;
input n_611;
input n_1126;
input n_1166;
input n_469;
input n_82;
input n_785;
input n_549;
input n_532;
input n_1161;
input n_1150;
input n_226;
input n_667;
input n_790;
input n_1055;
input n_111;
input n_880;
input n_544;
input n_1007;
input n_155;
input n_552;
input n_1198;
input n_1099;
input n_956;
input n_564;
input n_423;
input n_21;
input n_105;
input n_1021;
input n_4;
input n_551;
input n_688;
input n_800;
input n_671;
input n_819;
input n_1022;
input n_915;
input n_864;
input n_173;
input n_859;
input n_951;
input n_447;
input n_247;
input n_292;
input n_625;
input n_854;
input n_674;
input n_417;
input n_516;
input n_933;
input n_1152;
input n_497;
input n_606;
input n_275;
input n_26;
input n_877;
input n_2;
input n_755;
input n_1118;
input n_6;
input n_947;
input n_373;
input n_307;
input n_530;
input n_87;
input n_150;
input n_1107;
input n_556;
input n_1230;
input n_668;
input n_375;
input n_301;
input n_929;
input n_1124;
input n_902;
input n_191;
input n_1104;
input n_659;
input n_51;
input n_171;
input n_1182;
input n_579;
input n_938;
input n_1098;
input n_320;
input n_1154;
input n_1242;
input n_1135;
input n_24;
input n_406;
input n_519;
input n_1016;
input n_1243;
input n_546;
input n_101;
input n_281;
input n_240;
input n_291;
input n_231;
input n_257;
input n_731;
input n_371;
input n_709;
input n_317;
input n_1236;
input n_569;
input n_227;
input n_920;
input n_94;
input n_335;
input n_370;
input n_976;
input n_343;
input n_308;
input n_297;
input n_156;
input n_1078;
input n_775;
input n_219;
input n_157;
input n_600;
input n_223;
input n_264;
input n_955;
input n_163;
input n_339;
input n_1146;
input n_882;
input n_183;
input n_243;
input n_1036;
input n_1097;
input n_347;
input n_59;
input n_550;
input n_696;
input n_897;
input n_215;
input n_350;
input n_196;
input n_798;
input n_646;
input n_436;
input n_1216;
input n_290;
input n_580;
input n_1040;
input n_578;
input n_926;
input n_344;
input n_1218;
input n_422;
input n_475;
input n_777;
input n_1070;
input n_1030;
input n_72;
input n_415;
input n_1071;
input n_485;
input n_1165;
input n_496;
input n_958;
input n_1034;
input n_670;
input n_48;
input n_521;
input n_663;
input n_845;
input n_673;
input n_837;
input n_1239;
input n_528;
input n_680;
input n_395;
input n_164;
input n_553;
input n_901;
input n_813;
input n_214;
input n_675;
input n_888;
input n_1167;
input n_637;
input n_184;
input n_446;
input n_1064;
input n_144;
input n_858;
input n_114;
input n_96;
input n_923;
input n_691;
input n_1151;
input n_881;
input n_468;
input n_213;
input n_129;
input n_342;
input n_464;
input n_363;
input n_197;
input n_1069;
input n_1075;
input n_460;
input n_889;
input n_973;
input n_477;
input n_571;
input n_461;
input n_1211;
input n_1197;
input n_907;
input n_190;
input n_989;
input n_1039;
input n_34;
input n_228;
input n_283;
input n_488;
input n_736;
input n_892;
input n_1000;
input n_1202;
input n_1002;
input n_49;
input n_310;
input n_54;
input n_593;
input n_12;
input n_748;
input n_586;
input n_1058;
input n_838;
input n_332;
input n_1053;
input n_1224;
input n_349;
input n_1248;
input n_230;
input n_953;
input n_279;
input n_1014;
input n_1241;
input n_70;
input n_289;
input n_963;
input n_1052;
input n_954;
input n_627;
input n_440;
input n_793;
input n_478;
input n_476;
input n_534;
input n_884;
input n_345;
input n_944;
input n_91;
input n_182;
input n_143;
input n_647;
input n_237;
input n_407;
input n_1072;
input n_832;
input n_857;
input n_207;
input n_561;
input n_18;
input n_1027;
input n_971;
input n_1156;
input n_117;
input n_326;
input n_794;
input n_404;
input n_686;
input n_847;
input n_596;
input n_558;
input n_702;
input n_822;
input n_728;
input n_266;
input n_1162;
input n_272;
input n_1199;
input n_352;
input n_53;
input n_1038;
input n_520;
input n_409;
input n_887;
input n_154;
input n_71;
input n_300;
input n_809;
input n_870;
input n_931;
input n_599;
input n_434;
input n_868;
input n_639;
input n_914;
input n_411;
input n_414;
input n_965;
input n_935;
input n_121;
input n_1175;
input n_817;
input n_360;
input n_36;
input n_64;
input n_759;
input n_28;
input n_806;
input n_324;
input n_187;
input n_1189;
input n_103;
input n_97;
input n_11;
input n_7;
input n_706;
input n_746;
input n_747;
input n_52;
input n_784;
input n_110;
input n_1244;
input n_431;
input n_1194;
input n_615;
input n_851;
input n_843;
input n_523;
input n_913;
input n_705;
input n_865;
input n_61;
input n_678;
input n_697;
input n_127;
input n_1222;
input n_75;
input n_776;
input n_367;
input n_452;
input n_525;
input n_649;
input n_547;
input n_43;
input n_1191;
input n_116;
input n_284;
input n_1128;
input n_139;
input n_744;
input n_590;
input n_629;
input n_254;
input n_1233;
input n_23;
input n_526;
input n_293;
input n_372;
input n_677;
input n_244;
input n_47;
input n_1121;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_949;
input n_100;
input n_1008;
input n_946;
input n_1001;
input n_498;
input n_689;
input n_738;
input n_640;
input n_252;
input n_624;
input n_295;
input n_133;
input n_1010;
input n_1231;
input n_739;
input n_1195;
input n_610;
input n_936;
input n_568;
input n_39;
input n_1090;
input n_757;
input n_633;
input n_439;
input n_106;
input n_259;
input n_448;
input n_758;
input n_999;
input n_93;
input n_1158;
input n_563;
input n_1145;
input n_878;
input n_524;
input n_204;
input n_394;
input n_1049;
input n_1153;
input n_741;
input n_1068;
input n_122;
input n_331;
input n_10;
input n_906;
input n_1163;
input n_1207;
input n_919;
input n_908;
input n_90;
input n_724;
input n_658;
input n_456;
input n_959;
input n_535;
input n_152;
input n_940;
input n_9;
input n_592;
input n_1169;
input n_45;
input n_1017;
input n_123;
input n_978;
input n_1054;
input n_1095;
input n_267;
input n_514;
input n_457;
input n_1079;
input n_1045;
input n_1208;
input n_603;
input n_484;
input n_1033;
input n_442;
input n_131;
input n_636;
input n_660;
input n_1009;
input n_1148;
input n_109;
input n_742;
input n_750;
input n_995;
input n_454;
input n_374;
input n_185;
input n_396;
input n_1073;
input n_255;
input n_662;
input n_459;
input n_218;
input n_962;
input n_1215;
input n_1171;
input n_723;
input n_1065;
input n_473;
input n_1043;
input n_355;
input n_486;
input n_614;
input n_337;
input n_88;
input n_1177;
input n_168;
input n_974;
input n_727;
input n_1159;
input n_957;
input n_773;
input n_208;
input n_142;
input n_743;
input n_299;
input n_303;
input n_296;
input n_613;
input n_1119;
input n_1240;
input n_65;
input n_829;
input n_361;
input n_700;
input n_1237;
input n_573;
input n_69;
input n_1132;
input n_388;
input n_1127;
input n_761;
input n_1006;
input n_329;
input n_274;
input n_582;
input n_73;
input n_19;
input n_309;
input n_30;
input n_512;
input n_84;
input n_130;
input n_322;
input n_652;
input n_1111;
input n_25;
input n_1093;
input n_288;
input n_1031;
input n_263;
input n_609;
input n_1041;
input n_44;
input n_224;
input n_383;
input n_834;
input n_112;
input n_765;
input n_893;
input n_1015;
input n_1140;
input n_891;
input n_239;
input n_630;
input n_55;
input n_504;
input n_511;
input n_874;
input n_358;
input n_1101;
input n_77;
input n_102;
input n_1106;
input n_987;
input n_261;
input n_174;
input n_767;
input n_993;
input n_545;
input n_441;
input n_860;
input n_450;
input n_429;
input n_948;
input n_1217;
input n_628;
input n_365;
input n_729;
input n_1131;
input n_1084;
input n_970;
input n_911;
input n_83;
input n_513;
input n_1094;
input n_560;
input n_340;
input n_1044;
input n_1205;
input n_346;
input n_1209;
input n_495;
input n_602;
input n_574;
input n_879;
input n_16;
input n_58;
input n_623;
input n_405;
input n_824;
input n_359;
input n_490;
input n_996;
input n_921;
input n_233;
input n_572;
input n_366;
input n_815;
input n_128;
input n_120;
input n_327;
input n_135;
input n_1037;
input n_1080;
input n_426;
input n_1082;
input n_589;
input n_716;
input n_562;
input n_62;
input n_952;
input n_1229;
input n_391;
input n_701;
input n_1023;
input n_645;
input n_539;
input n_803;
input n_1092;
input n_238;
input n_531;
input n_890;
input n_764;
input n_1056;
input n_162;
input n_960;
input n_222;
input n_1123;
input n_1047;
input n_634;
input n_199;
input n_32;
input n_348;
input n_1029;
input n_925;
input n_1206;
input n_424;
input n_256;
input n_950;
input n_380;
input n_419;
input n_444;
input n_1060;
input n_1141;
input n_316;
input n_389;
input n_418;
input n_248;
input n_136;
input n_86;
input n_146;
input n_912;
input n_315;
input n_968;
input n_451;
input n_619;
input n_408;
input n_376;
input n_967;
input n_74;
input n_1139;
input n_515;
input n_57;
input n_351;
input n_885;
input n_397;
input n_483;
input n_683;
input n_1057;
input n_1051;
input n_1085;
input n_1066;
input n_721;
input n_1157;
input n_841;
input n_1050;
input n_22;
input n_802;
input n_46;
input n_983;
input n_38;
input n_280;
input n_873;
input n_378;
input n_1112;
input n_762;
input n_17;
input n_690;
input n_33;
input n_583;
input n_302;
input n_1203;
input n_821;
input n_321;
input n_1179;
input n_621;
input n_753;
input n_455;
input n_1048;
input n_212;
input n_385;
input n_507;
input n_330;
input n_1228;
input n_972;
input n_692;
input n_820;
input n_1200;
input n_1185;
input n_991;
input n_828;
input n_779;
input n_576;
input n_1143;
input n_804;
input n_537;
input n_945;
input n_492;
input n_153;
input n_943;
input n_341;
input n_250;
input n_992;
input n_543;
input n_260;
input n_842;
input n_650;
input n_984;
input n_694;
input n_286;
input n_883;
input n_470;
input n_325;
input n_449;
input n_132;
input n_1214;
input n_900;
input n_856;
input n_918;
input n_942;
input n_189;
input n_1147;
input n_13;
input n_1077;
input n_540;
input n_618;
input n_896;
input n_323;
input n_195;
input n_356;
input n_894;
input n_831;
input n_964;
input n_1096;
input n_234;
input n_833;
input n_5;
input n_225;
input n_988;
input n_814;
input n_192;
input n_1201;
input n_1114;
input n_655;
input n_669;
input n_472;
input n_1176;
input n_387;
input n_1149;
input n_398;
input n_635;
input n_763;
input n_1020;
input n_1062;
input n_211;
input n_1219;
input n_3;
input n_1204;
input n_178;
input n_1035;
input n_287;
input n_555;
input n_783;
input n_1188;
input n_661;
input n_41;
input n_849;
input n_15;
input n_336;
input n_584;
input n_681;
input n_50;
input n_430;
input n_510;
input n_216;
input n_311;
input n_830;
input n_801;
input n_241;
input n_875;
input n_357;
input n_1110;
input n_445;
input n_749;
input n_1134;
input n_717;
input n_165;
input n_939;
input n_482;
input n_1088;
input n_588;
input n_1173;
input n_789;
input n_1232;
input n_734;
input n_638;
input n_866;
input n_107;
input n_969;
input n_1019;
input n_1105;
input n_249;
input n_304;
input n_577;
input n_338;
input n_149;
input n_693;
input n_14;
input n_836;
input n_990;
input n_975;
input n_567;
input n_778;
input n_1122;
input n_151;
input n_306;
input n_458;
input n_770;
input n_1102;
input n_711;
input n_85;
input n_1187;
input n_1164;
input n_489;
input n_1174;
input n_617;
input n_876;
input n_1190;
input n_118;
input n_601;
input n_917;
input n_966;
input n_253;
input n_1116;
input n_1212;
input n_172;
input n_206;
input n_217;
input n_726;
input n_982;
input n_818;
input n_861;
input n_1183;
input n_899;
input n_210;
input n_774;
input n_1059;
input n_176;
input n_1133;
input n_557;
input n_1005;
input n_607;
input n_1003;
input n_679;
input n_710;
input n_527;
input n_1168;
input n_707;
input n_937;
input n_393;
input n_108;
input n_487;
input n_665;
input n_66;
input n_177;
input n_421;
input n_910;
input n_768;
input n_205;
input n_1136;
input n_754;
input n_179;
input n_1125;
input n_125;
input n_410;
input n_708;
input n_529;
input n_735;
input n_232;
input n_1109;
input n_126;
input n_895;
input n_202;
input n_427;
input n_791;
input n_732;
input n_193;
input n_808;
input n_797;
input n_1025;
input n_500;
input n_1067;
input n_148;
input n_435;
input n_159;
input n_766;
input n_541;
input n_538;
input n_1117;
input n_799;
input n_687;
input n_715;
input n_1213;
input n_536;
input n_872;
input n_594;
input n_200;
input n_1155;
input n_89;
input n_115;
input n_1011;
input n_1184;
input n_985;
input n_869;
input n_810;
input n_416;
input n_827;
input n_401;
input n_626;
input n_1144;
input n_1137;
input n_1170;
input n_305;
input n_137;
input n_676;
input n_294;
input n_318;
input n_653;
input n_642;
input n_194;
input n_855;
input n_1178;
input n_850;
input n_684;
input n_124;
input n_268;
input n_664;
input n_503;
input n_235;
input n_605;
input n_353;
input n_620;
input n_643;
input n_916;
input n_1081;
input n_493;
input n_1235;
input n_703;
input n_698;
input n_980;
input n_1115;
input n_780;
input n_998;
input n_467;
input n_1227;
input n_840;
input n_501;
input n_823;
input n_245;
input n_725;
input n_672;
input n_581;
input n_382;
input n_554;
input n_898;
input n_1013;
input n_718;
input n_265;
input n_1120;
input n_719;
input n_443;
input n_198;
input n_714;
input n_909;
input n_997;
input n_932;
input n_612;
input n_788;
input n_119;
input n_559;
input n_825;
input n_508;
input n_506;
input n_737;
input n_986;
input n_509;
input n_147;
input n_67;
input n_1192;
input n_1024;
input n_1063;
input n_209;
input n_733;
input n_941;
input n_981;
input n_68;
input n_867;
input n_186;
input n_134;
input n_587;
input n_63;
input n_792;
input n_756;
input n_399;
input n_1238;
input n_548;
input n_812;
input n_298;
input n_518;
input n_505;
input n_282;
input n_752;
input n_905;
input n_1108;
input n_782;
input n_1100;
input n_862;
input n_760;
input n_381;
input n_220;
input n_390;
input n_31;
input n_481;
input n_769;
input n_42;
input n_1046;
input n_271;
input n_934;
input n_826;
input n_886;
input n_1221;
input n_654;
input n_1172;
input n_167;
input n_379;
input n_428;
input n_570;
input n_853;
input n_377;
input n_751;
input n_786;
input n_1083;
input n_1142;
input n_1129;
input n_392;
input n_158;
input n_704;
input n_787;
input n_138;
input n_961;
input n_771;
input n_276;
input n_95;
input n_1225;
input n_169;
input n_522;
input n_400;
input n_930;
input n_181;
input n_221;
input n_622;
input n_1087;
input n_386;
input n_994;
input n_848;
input n_1223;
input n_104;
input n_682;
input n_56;
input n_141;
input n_1247;
input n_922;
input n_816;
input n_591;
input n_145;
input n_313;
input n_631;
input n_479;
input n_1246;
input n_432;
input n_839;
input n_1210;
input n_328;
input n_140;
input n_369;
input n_871;
input n_598;
input n_685;
input n_928;
input n_608;
input n_78;
input n_772;
input n_499;
input n_517;
input n_98;
input n_402;
input n_413;
input n_1086;
input n_796;
input n_236;
input n_1012;
input n_1;
input n_903;
input n_740;
input n_203;
input n_384;
input n_80;
input n_35;
input n_277;
input n_1061;
input n_92;
input n_333;
input n_462;
input n_1193;
input n_258;
input n_1113;
input n_29;
input n_79;
input n_1226;
input n_722;
input n_188;
input n_844;
input n_201;
input n_471;
input n_852;
input n_40;
input n_1028;
input n_781;
input n_474;
input n_542;
input n_463;
input n_595;
input n_502;
input n_466;
input n_420;
input n_632;
input n_699;
input n_979;
input n_1245;
input n_846;
input n_465;
input n_76;
input n_362;
input n_170;
input n_27;
input n_161;
input n_273;
input n_585;
input n_270;
input n_616;
input n_81;
input n_745;
input n_1103;
input n_648;
input n_312;
input n_1076;
input n_1091;
input n_494;
input n_641;
input n_730;
input n_354;
input n_575;
input n_480;
input n_425;
input n_795;
input n_695;
input n_180;
input n_656;
input n_1220;
input n_37;
input n_229;
input n_437;
input n_60;
input n_403;
input n_453;
input n_1130;
input n_720;
input n_0;
input n_863;
input n_805;
input n_113;
input n_712;
input n_246;
input n_1042;
input n_269;
input n_285;
input n_412;
input n_657;
input n_644;
input n_1160;
input n_491;
input n_1074;
input n_251;
input n_160;
input n_566;
input n_565;
input n_597;
input n_1181;
input n_1196;
input n_651;
input n_334;
input n_811;
input n_807;
input n_835;
input n_175;
input n_666;
input n_262;
input n_99;
input n_1026;
input n_1234;
input n_319;
input n_364;
input n_1138;
input n_927;
input n_20;
input n_1089;
input n_1004;
input n_1186;
input n_1032;
input n_242;
input n_1018;
input n_438;
input n_713;
input n_904;
input n_166;
input n_1180;
input n_533;
input n_278;

output n_5372;

wire n_2253;
wire n_2417;
wire n_2756;
wire n_4706;
wire n_2380;
wire n_3241;
wire n_3006;
wire n_5287;
wire n_2327;
wire n_1488;
wire n_2899;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_2395;
wire n_5161;
wire n_5207;
wire n_2347;
wire n_4963;
wire n_4240;
wire n_4508;
wire n_2021;
wire n_2391;
wire n_5035;
wire n_5282;
wire n_1960;
wire n_2843;
wire n_3615;
wire n_2059;
wire n_1466;
wire n_2487;
wire n_1695;
wire n_3202;
wire n_4977;
wire n_3813;
wire n_3341;
wire n_3587;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_4145;
wire n_3785;
wire n_5033;
wire n_1462;
wire n_4211;
wire n_3448;
wire n_3019;
wire n_2096;
wire n_3776;
wire n_2530;
wire n_4517;
wire n_2483;
wire n_1696;
wire n_4425;
wire n_4950;
wire n_4988;
wire n_1285;
wire n_1860;
wire n_4615;
wire n_1728;
wire n_2076;
wire n_2147;
wire n_3010;
wire n_2770;
wire n_4131;
wire n_2584;
wire n_3188;
wire n_3403;
wire n_3624;
wire n_3461;
wire n_3082;
wire n_2189;
wire n_3796;
wire n_5154;
wire n_3283;
wire n_2323;
wire n_2597;
wire n_3340;
wire n_3277;
wire n_2052;
wire n_4499;
wire n_4927;
wire n_5202;
wire n_1314;
wire n_1512;
wire n_1490;
wire n_3214;
wire n_2091;
wire n_1517;
wire n_4311;
wire n_3631;
wire n_3806;
wire n_4691;
wire n_1449;
wire n_4678;
wire n_2032;
wire n_1566;
wire n_2587;
wire n_3947;
wire n_3490;
wire n_3868;
wire n_1948;
wire n_3183;
wire n_3437;
wire n_3353;
wire n_4203;
wire n_3687;
wire n_5241;
wire n_2384;
wire n_3156;
wire n_3376;
wire n_5037;
wire n_4468;
wire n_3653;
wire n_3702;
wire n_4976;
wire n_2202;
wire n_2648;
wire n_5008;
wire n_2159;
wire n_2976;
wire n_3876;
wire n_2353;
wire n_2439;
wire n_4811;
wire n_2276;
wire n_2089;
wire n_3420;
wire n_1561;
wire n_5144;
wire n_3361;
wire n_4758;
wire n_1600;
wire n_4255;
wire n_1796;
wire n_4484;
wire n_3668;
wire n_4237;
wire n_2934;
wire n_1672;
wire n_1880;
wire n_3550;
wire n_1626;
wire n_2079;
wire n_2238;
wire n_1405;
wire n_1706;
wire n_3418;
wire n_4901;
wire n_2859;
wire n_3395;
wire n_4917;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_2968;
wire n_1585;
wire n_2684;
wire n_3593;
wire n_5343;
wire n_1599;
wire n_4421;
wire n_4836;
wire n_5062;
wire n_4020;
wire n_2730;
wire n_2251;
wire n_3915;
wire n_1377;
wire n_4469;
wire n_4414;
wire n_5184;
wire n_4532;
wire n_3339;
wire n_3349;
wire n_3735;
wire n_2248;
wire n_3007;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_2100;
wire n_5236;
wire n_3310;
wire n_3487;
wire n_2258;
wire n_1667;
wire n_3983;
wire n_4405;
wire n_1926;
wire n_1331;
wire n_4195;
wire n_4969;
wire n_4504;
wire n_1385;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_4531;
wire n_2987;
wire n_1527;
wire n_4567;
wire n_4164;
wire n_5315;
wire n_4234;
wire n_4130;
wire n_3611;
wire n_2862;
wire n_5348;
wire n_2175;
wire n_5055;
wire n_2324;
wire n_2606;
wire n_3187;
wire n_2828;
wire n_4471;
wire n_5031;
wire n_3392;
wire n_3975;
wire n_3430;
wire n_4444;
wire n_3208;
wire n_3331;
wire n_2379;
wire n_4983;
wire n_2911;
wire n_2154;
wire n_4916;
wire n_3649;
wire n_4302;
wire n_2514;
wire n_5189;
wire n_4786;
wire n_3257;
wire n_4160;
wire n_2293;
wire n_4051;
wire n_2028;
wire n_3009;
wire n_1276;
wire n_1412;
wire n_3981;
wire n_1841;
wire n_2581;
wire n_3224;
wire n_4647;
wire n_3752;
wire n_1711;
wire n_1891;
wire n_5254;
wire n_3526;
wire n_2546;
wire n_3790;
wire n_3491;
wire n_4613;
wire n_4649;
wire n_1888;
wire n_1963;
wire n_4795;
wire n_2226;
wire n_2891;
wire n_4028;
wire n_1690;
wire n_3819;
wire n_2449;
wire n_5083;
wire n_2297;
wire n_4186;
wire n_4731;
wire n_1759;
wire n_2177;
wire n_3747;
wire n_2227;
wire n_4618;
wire n_2190;
wire n_3346;
wire n_4742;
wire n_2876;
wire n_4099;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_2479;
wire n_1464;
wire n_4295;
wire n_5303;
wire n_1444;
wire n_4694;
wire n_4533;
wire n_3038;
wire n_5081;
wire n_5124;
wire n_3068;
wire n_2871;
wire n_4244;
wire n_4603;
wire n_2943;
wire n_4254;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_4697;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_4810;
wire n_3317;
wire n_4391;
wire n_3263;
wire n_2582;
wire n_4157;
wire n_4283;
wire n_4681;
wire n_1503;
wire n_4638;
wire n_1468;
wire n_3455;
wire n_5047;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_5346;
wire n_1994;
wire n_4707;
wire n_2577;
wire n_4527;
wire n_5109;
wire n_2796;
wire n_2342;
wire n_4156;
wire n_1851;
wire n_4848;
wire n_2937;
wire n_3095;
wire n_2805;
wire n_4918;
wire n_3856;
wire n_2914;
wire n_4898;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_5010;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_2925;
wire n_3773;
wire n_3918;
wire n_2398;
wire n_2857;
wire n_5358;
wire n_4528;
wire n_3932;
wire n_4619;
wire n_4673;
wire n_3516;
wire n_4822;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1596;
wire n_2947;
wire n_4299;
wire n_4801;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_3515;
wire n_2886;
wire n_2093;
wire n_2473;
wire n_3287;
wire n_3378;
wire n_1431;
wire n_4279;
wire n_4769;
wire n_4632;
wire n_4294;
wire n_1732;
wire n_5279;
wire n_4125;
wire n_4232;
wire n_4949;
wire n_2941;
wire n_2457;
wire n_4790;
wire n_2536;
wire n_1336;
wire n_1758;
wire n_2952;
wire n_4847;
wire n_5321;
wire n_3058;
wire n_5096;
wire n_4365;
wire n_1878;
wire n_3505;
wire n_4610;
wire n_3730;
wire n_4489;
wire n_5210;
wire n_4967;
wire n_4992;
wire n_3001;
wire n_3945;
wire n_4542;
wire n_2261;
wire n_2729;
wire n_3597;
wire n_1612;
wire n_2897;
wire n_2077;
wire n_4198;
wire n_2909;
wire n_4534;
wire n_4500;
wire n_5014;
wire n_3185;
wire n_1300;
wire n_3523;
wire n_1785;
wire n_2829;
wire n_4597;
wire n_4329;
wire n_4087;
wire n_3811;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_2231;
wire n_2017;
wire n_2604;
wire n_4257;
wire n_3453;
wire n_2390;
wire n_3213;
wire n_3077;
wire n_1562;
wire n_3474;
wire n_3984;
wire n_2151;
wire n_2106;
wire n_2716;
wire n_4665;
wire n_1913;
wire n_1823;
wire n_3679;
wire n_3422;
wire n_3888;
wire n_4189;
wire n_1875;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_3707;
wire n_1846;
wire n_3429;
wire n_1903;
wire n_3849;
wire n_3946;
wire n_3229;
wire n_4463;
wire n_1805;
wire n_4687;
wire n_4670;
wire n_4084;
wire n_4703;
wire n_4037;
wire n_2922;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2727;
wire n_3421;
wire n_2240;
wire n_2436;
wire n_1552;
wire n_3618;
wire n_2593;
wire n_5262;
wire n_3683;
wire n_3642;
wire n_3286;
wire n_3808;
wire n_1327;
wire n_4763;
wire n_1684;
wire n_3590;
wire n_5310;
wire n_4594;
wire n_3424;
wire n_1381;
wire n_2301;
wire n_3583;
wire n_3560;
wire n_4076;
wire n_4714;
wire n_2419;
wire n_3215;
wire n_5146;
wire n_4776;
wire n_2122;
wire n_2512;
wire n_4102;
wire n_2786;
wire n_3171;
wire n_1437;
wire n_5213;
wire n_3020;
wire n_3677;
wire n_3462;
wire n_3468;
wire n_2910;
wire n_1893;
wire n_1467;
wire n_2163;
wire n_2254;
wire n_1382;
wire n_3546;
wire n_2647;
wire n_1311;
wire n_1519;
wire n_4443;
wire n_4507;
wire n_2443;
wire n_1811;
wire n_2624;
wire n_3012;
wire n_4575;
wire n_3244;
wire n_3130;
wire n_3822;
wire n_3569;
wire n_4452;
wire n_4348;
wire n_5362;
wire n_4355;
wire n_3494;
wire n_5050;
wire n_5063;
wire n_5229;
wire n_2125;
wire n_3771;
wire n_5199;
wire n_3110;
wire n_3073;
wire n_4572;
wire n_4026;
wire n_2265;
wire n_4104;
wire n_1608;
wire n_4512;
wire n_3554;
wire n_4377;
wire n_1305;
wire n_5266;
wire n_3178;
wire n_5355;
wire n_2334;
wire n_4521;
wire n_4488;
wire n_2289;
wire n_3051;
wire n_1343;
wire n_2783;
wire n_2263;
wire n_3750;
wire n_2341;
wire n_3632;
wire n_4588;
wire n_2733;
wire n_1288;
wire n_2785;
wire n_2415;
wire n_3299;
wire n_4519;
wire n_3715;
wire n_3040;
wire n_1938;
wire n_2499;
wire n_3568;
wire n_3737;
wire n_1967;
wire n_1329;
wire n_3255;
wire n_4856;
wire n_2997;
wire n_4400;
wire n_5168;
wire n_3326;
wire n_3734;
wire n_4778;
wire n_2429;
wire n_5322;
wire n_1793;
wire n_4352;
wire n_4441;
wire n_4761;
wire n_1804;
wire n_4347;
wire n_4095;
wire n_3196;
wire n_4593;
wire n_2364;
wire n_2533;
wire n_3492;
wire n_2780;
wire n_4727;
wire n_4568;
wire n_5371;
wire n_2291;
wire n_4043;
wire n_1636;
wire n_3601;
wire n_1350;
wire n_1865;
wire n_2973;
wire n_2094;
wire n_1575;
wire n_2393;
wire n_1697;
wire n_5316;
wire n_3831;
wire n_3801;
wire n_2043;
wire n_2751;
wire n_4893;
wire n_5032;
wire n_1549;
wire n_1934;
wire n_4948;
wire n_4000;
wire n_3240;
wire n_2025;
wire n_1446;
wire n_4406;
wire n_2758;
wire n_1458;
wire n_1807;
wire n_2618;
wire n_5112;
wire n_2559;
wire n_4748;
wire n_2295;
wire n_3931;
wire n_4010;
wire n_2840;
wire n_5017;
wire n_1814;
wire n_2822;
wire n_4710;
wire n_4607;
wire n_5123;
wire n_4117;
wire n_3636;
wire n_1722;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_4487;
wire n_5001;
wire n_2795;
wire n_2981;
wire n_2282;
wire n_2800;
wire n_4817;
wire n_3380;
wire n_2098;
wire n_1296;
wire n_3460;
wire n_3409;
wire n_3538;
wire n_2068;
wire n_4849;
wire n_4867;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_4728;
wire n_4247;
wire n_4933;
wire n_4018;
wire n_3900;
wire n_4902;
wire n_4518;
wire n_4409;
wire n_4411;
wire n_3872;
wire n_4336;
wire n_2270;
wire n_4777;
wire n_2653;
wire n_2496;
wire n_1908;
wire n_2259;
wire n_3877;
wire n_2995;
wire n_2494;
wire n_3547;
wire n_3977;
wire n_4052;
wire n_3459;
wire n_1499;
wire n_4398;
wire n_3155;
wire n_2633;
wire n_4954;
wire n_2435;
wire n_1392;
wire n_2097;
wire n_4304;
wire n_3911;
wire n_5333;
wire n_1303;
wire n_4431;
wire n_4192;
wire n_3736;
wire n_4805;
wire n_4885;
wire n_1661;
wire n_3565;
wire n_4701;
wire n_2575;
wire n_5040;
wire n_1658;
wire n_1904;
wire n_1345;
wire n_1899;
wire n_2067;
wire n_2219;
wire n_3533;
wire n_2877;
wire n_2148;
wire n_1726;
wire n_4631;
wire n_3035;
wire n_5194;
wire n_1657;
wire n_1475;
wire n_1725;
wire n_1313;
wire n_1491;
wire n_3639;
wire n_2501;
wire n_3079;
wire n_4965;
wire n_1915;
wire n_5239;
wire n_1310;
wire n_2605;
wire n_4747;
wire n_5197;
wire n_1399;
wire n_1979;
wire n_2924;
wire n_4111;
wire n_2484;
wire n_4587;
wire n_3731;
wire n_2946;
wire n_5305;
wire n_4538;
wire n_2754;
wire n_1742;
wire n_2489;
wire n_5204;
wire n_2012;
wire n_1291;
wire n_4094;
wire n_3503;
wire n_2866;
wire n_3561;
wire n_1418;
wire n_2917;
wire n_2425;
wire n_3536;
wire n_3661;
wire n_4150;
wire n_4878;
wire n_1703;
wire n_1650;
wire n_3934;
wire n_4985;
wire n_3922;
wire n_3846;
wire n_2103;
wire n_2160;
wire n_2498;
wire n_2697;
wire n_3074;
wire n_1999;
wire n_2372;
wire n_3673;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_3943;
wire n_2430;
wire n_2433;
wire n_3293;
wire n_4022;
wire n_1531;
wire n_1334;
wire n_4852;
wire n_2528;
wire n_4869;
wire n_4700;
wire n_4035;
wire n_2316;
wire n_1898;
wire n_3294;
wire n_4426;
wire n_3415;
wire n_2284;
wire n_2817;
wire n_3139;
wire n_5292;
wire n_2598;
wire n_4601;
wire n_2687;
wire n_1890;
wire n_4220;
wire n_1944;
wire n_1497;
wire n_3431;
wire n_3169;
wire n_3151;
wire n_2078;
wire n_3284;
wire n_3070;
wire n_4066;
wire n_2884;
wire n_4515;
wire n_4351;
wire n_5264;
wire n_3126;
wire n_4403;
wire n_1981;
wire n_1663;
wire n_1718;
wire n_4509;
wire n_4858;
wire n_3700;
wire n_1518;
wire n_4223;
wire n_1281;
wire n_1889;
wire n_1489;
wire n_5025;
wire n_2966;
wire n_1376;
wire n_2326;
wire n_1569;
wire n_2188;
wire n_1429;
wire n_4644;
wire n_4456;
wire n_5060;
wire n_5334;
wire n_2448;
wire n_4346;
wire n_3170;
wire n_2748;
wire n_3311;
wire n_3272;
wire n_2898;
wire n_2717;
wire n_1861;
wire n_3628;
wire n_3691;
wire n_4235;
wire n_1867;
wire n_1945;
wire n_3018;
wire n_2573;
wire n_4435;
wire n_2939;
wire n_3807;
wire n_2447;
wire n_4764;
wire n_2774;
wire n_1707;
wire n_4655;
wire n_3161;
wire n_4581;
wire n_4827;
wire n_2488;
wire n_3477;
wire n_2476;
wire n_4399;
wire n_2781;
wire n_5309;
wire n_2778;
wire n_4782;
wire n_1520;
wire n_4363;
wire n_2887;
wire n_1287;
wire n_4864;
wire n_1262;
wire n_2691;
wire n_1411;
wire n_3054;
wire n_4335;
wire n_2526;
wire n_2703;
wire n_2167;
wire n_3391;
wire n_4259;
wire n_2709;
wire n_1536;
wire n_4865;
wire n_4056;
wire n_1344;
wire n_4564;
wire n_3840;
wire n_1339;
wire n_5085;
wire n_3518;
wire n_2956;
wire n_3733;
wire n_2173;
wire n_1842;
wire n_3738;
wire n_5116;
wire n_3464;
wire n_2018;
wire n_4526;
wire n_1555;
wire n_3245;
wire n_4417;
wire n_4899;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_2453;
wire n_4798;
wire n_1525;
wire n_3509;
wire n_3352;
wire n_3076;
wire n_3535;
wire n_2182;
wire n_3251;
wire n_2931;
wire n_5185;
wire n_3118;
wire n_3511;
wire n_3443;
wire n_2146;
wire n_1487;
wire n_3644;
wire n_5076;
wire n_3336;
wire n_3935;
wire n_3521;
wire n_3562;
wire n_3948;
wire n_4750;
wire n_1515;
wire n_2918;
wire n_3232;
wire n_1673;
wire n_2112;
wire n_1739;
wire n_2958;
wire n_4981;
wire n_3114;
wire n_3125;
wire n_2394;
wire n_3612;
wire n_2954;
wire n_4835;
wire n_4430;
wire n_4081;
wire n_3132;
wire n_4407;
wire n_3951;
wire n_4894;
wire n_3238;
wire n_3210;
wire n_2036;
wire n_3267;
wire n_4995;
wire n_3964;
wire n_3772;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_4446;
wire n_3884;
wire n_3726;
wire n_2525;
wire n_2892;
wire n_2907;
wire n_3577;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1741;
wire n_4057;
wire n_4332;
wire n_1258;
wire n_4314;
wire n_3347;
wire n_3216;
wire n_1621;
wire n_3809;
wire n_2113;
wire n_1448;
wire n_4288;
wire n_3567;
wire n_5066;
wire n_1634;
wire n_3939;
wire n_4241;
wire n_3321;
wire n_3212;
wire n_1433;
wire n_2256;
wire n_3152;
wire n_5106;
wire n_2920;
wire n_4265;
wire n_5319;
wire n_2247;
wire n_1622;
wire n_3705;
wire n_2802;
wire n_4705;
wire n_3159;
wire n_2268;
wire n_3778;
wire n_5337;
wire n_3304;
wire n_1378;
wire n_3912;
wire n_1729;
wire n_2739;
wire n_2771;
wire n_4604;
wire n_5223;
wire n_3795;
wire n_5020;
wire n_4419;
wire n_4477;
wire n_3179;
wire n_3256;
wire n_2386;
wire n_1501;
wire n_3086;
wire n_2369;
wire n_2927;
wire n_4217;
wire n_4395;
wire n_2821;
wire n_5074;
wire n_2568;
wire n_5364;
wire n_1738;
wire n_3728;
wire n_3064;
wire n_3088;
wire n_4639;
wire n_3713;
wire n_3663;
wire n_5046;
wire n_5166;
wire n_3246;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_5088;
wire n_2302;
wire n_1494;
wire n_2069;
wire n_3434;
wire n_1806;
wire n_1563;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_2024;
wire n_4780;
wire n_4243;
wire n_4982;
wire n_3695;
wire n_4330;
wire n_2482;
wire n_2677;
wire n_3832;
wire n_3987;
wire n_5352;
wire n_4991;
wire n_1698;
wire n_2329;
wire n_2142;
wire n_3332;
wire n_3048;
wire n_3937;
wire n_2203;
wire n_4525;
wire n_3782;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_3786;
wire n_2888;
wire n_3638;
wire n_1633;
wire n_4177;
wire n_3763;
wire n_2669;
wire n_1778;
wire n_2306;
wire n_3022;
wire n_4264;
wire n_3087;
wire n_3489;
wire n_2566;
wire n_5129;
wire n_2149;
wire n_3060;
wire n_4276;
wire n_5219;
wire n_3013;
wire n_1984;
wire n_5170;
wire n_2408;
wire n_5320;
wire n_1877;
wire n_3049;
wire n_1723;
wire n_5107;
wire n_4485;
wire n_4626;
wire n_2659;
wire n_1414;
wire n_4975;
wire n_1852;
wire n_3089;
wire n_2470;
wire n_3985;
wire n_5253;
wire n_1391;
wire n_4760;
wire n_4652;
wire n_4624;
wire n_2551;
wire n_1587;
wire n_2682;
wire n_1284;
wire n_3440;
wire n_1748;
wire n_4569;
wire n_2699;
wire n_4897;
wire n_2769;
wire n_3542;
wire n_3436;
wire n_2615;
wire n_3940;
wire n_2985;
wire n_5065;
wire n_2753;
wire n_1582;
wire n_3637;
wire n_2842;
wire n_4523;
wire n_1836;
wire n_2868;
wire n_3141;
wire n_5084;
wire n_3164;
wire n_3570;
wire n_5260;
wire n_4919;
wire n_4025;
wire n_2712;
wire n_5328;
wire n_3936;
wire n_4503;
wire n_3507;
wire n_3821;
wire n_2700;
wire n_3367;
wire n_4464;
wire n_3096;
wire n_3496;
wire n_4114;
wire n_2544;
wire n_2356;
wire n_4556;
wire n_2620;
wire n_1581;
wire n_4089;
wire n_2919;
wire n_4327;
wire n_4218;
wire n_2150;
wire n_3146;
wire n_5165;
wire n_2241;
wire n_2757;
wire n_4353;
wire n_2042;
wire n_1754;
wire n_1623;
wire n_2921;
wire n_2720;
wire n_1854;
wire n_4990;
wire n_1856;
wire n_4959;
wire n_4161;
wire n_1319;
wire n_3992;
wire n_2616;
wire n_1906;
wire n_4103;
wire n_1387;
wire n_4466;
wire n_2262;
wire n_2462;
wire n_1532;
wire n_3625;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_2837;
wire n_4844;
wire n_2979;
wire n_5257;
wire n_3655;
wire n_4688;
wire n_4765;
wire n_2548;
wire n_5180;
wire n_2108;
wire n_3640;
wire n_4388;
wire n_4206;
wire n_1538;
wire n_1779;
wire n_4738;
wire n_1369;
wire n_3909;
wire n_3207;
wire n_3944;
wire n_4434;
wire n_4837;
wire n_3042;
wire n_1942;
wire n_2510;
wire n_4219;
wire n_2804;
wire n_3659;
wire n_2120;
wire n_5012;
wire n_1293;
wire n_1876;
wire n_4620;
wire n_1810;
wire n_2813;
wire n_4438;
wire n_2009;
wire n_2222;
wire n_3510;
wire n_3218;
wire n_2667;
wire n_3150;
wire n_4325;
wire n_1733;
wire n_2413;
wire n_3775;
wire n_4133;
wire n_4184;
wire n_5203;
wire n_2518;
wire n_2629;
wire n_4481;
wire n_3416;
wire n_4379;
wire n_2181;
wire n_1829;
wire n_4030;
wire n_4490;
wire n_3138;
wire n_4397;
wire n_1710;
wire n_2928;
wire n_1734;
wire n_4820;
wire n_3770;
wire n_1308;
wire n_5094;
wire n_4938;
wire n_4179;
wire n_3469;
wire n_5336;
wire n_2723;
wire n_3220;
wire n_4641;
wire n_2539;
wire n_3855;
wire n_2054;
wire n_5339;
wire n_1559;
wire n_4931;
wire n_1765;
wire n_3158;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_3113;
wire n_2718;
wire n_3760;
wire n_4078;
wire n_1760;
wire n_2856;
wire n_1832;
wire n_4146;
wire n_4360;
wire n_3666;
wire n_3828;
wire n_3288;
wire n_4404;
wire n_5091;
wire n_1509;
wire n_1874;
wire n_4787;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_3667;
wire n_1306;
wire n_3703;
wire n_4903;
wire n_3558;
wire n_2545;
wire n_2787;
wire n_4356;
wire n_2061;
wire n_4432;
wire n_5251;
wire n_2378;
wire n_1740;
wire n_1586;
wire n_4291;
wire n_4386;
wire n_4149;
wire n_1492;
wire n_1692;
wire n_2982;
wire n_2481;
wire n_3545;
wire n_2507;
wire n_4019;
wire n_2900;
wire n_1614;
wire n_2339;
wire n_4637;
wire n_4935;
wire n_4785;
wire n_3426;
wire n_3454;
wire n_3820;
wire n_3741;
wire n_3410;
wire n_2029;
wire n_1609;
wire n_5298;
wire n_1887;
wire n_4413;
wire n_2346;
wire n_3990;
wire n_4493;
wire n_3475;
wire n_1592;
wire n_2882;
wire n_1721;
wire n_2338;
wire n_3672;
wire n_5290;
wire n_3197;
wire n_3109;
wire n_2721;
wire n_5095;
wire n_3002;
wire n_5324;
wire n_3897;
wire n_3845;
wire n_2081;
wire n_4570;
wire n_2156;
wire n_5101;
wire n_4296;
wire n_1820;
wire n_5019;
wire n_2418;
wire n_2179;
wire n_1416;
wire n_1724;
wire n_2521;
wire n_3458;
wire n_1420;
wire n_3330;
wire n_4606;
wire n_4774;
wire n_2477;
wire n_3887;
wire n_4093;
wire n_1486;
wire n_4672;
wire n_3519;
wire n_4174;
wire n_3374;
wire n_3045;
wire n_2367;
wire n_1870;
wire n_4766;
wire n_2896;
wire n_1365;
wire n_4074;
wire n_4600;
wire n_1927;
wire n_1349;
wire n_4460;
wire n_3645;
wire n_3223;
wire n_3929;
wire n_2255;
wire n_2272;
wire n_1965;
wire n_1902;
wire n_1941;
wire n_3938;
wire n_2878;
wire n_3498;
wire n_2015;
wire n_1982;
wire n_4110;
wire n_3189;
wire n_2066;
wire n_3154;
wire n_1551;
wire n_2905;
wire n_3965;
wire n_3566;
wire n_2220;
wire n_4349;
wire n_3788;
wire n_2410;
wire n_4313;
wire n_1935;
wire n_3366;
wire n_1534;
wire n_1351;
wire n_2696;
wire n_4863;
wire n_3242;
wire n_3525;
wire n_3486;
wire n_2405;
wire n_3995;
wire n_2088;
wire n_2953;
wire n_4036;
wire n_5100;
wire n_1795;
wire n_2578;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_3478;
wire n_4015;
wire n_3890;
wire n_2740;
wire n_5367;
wire n_2656;
wire n_1274;
wire n_3524;
wire n_5034;
wire n_1708;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_2092;
wire n_2075;
wire n_3658;
wire n_1776;
wire n_4807;
wire n_2281;
wire n_2131;
wire n_3026;
wire n_1757;
wire n_1919;
wire n_4230;
wire n_3419;
wire n_1290;
wire n_2053;
wire n_1958;
wire n_1252;
wire n_3784;
wire n_2969;
wire n_3941;
wire n_2864;
wire n_3195;
wire n_3190;
wire n_1553;
wire n_3678;
wire n_2664;
wire n_3456;
wire n_1808;
wire n_2266;
wire n_2650;
wire n_4428;
wire n_5003;
wire n_5252;
wire n_2731;
wire n_5134;
wire n_3953;
wire n_3166;
wire n_4122;
wire n_3976;
wire n_1357;
wire n_3979;
wire n_4582;
wire n_2998;
wire n_4684;
wire n_4840;
wire n_3162;
wire n_2760;
wire n_3377;
wire n_3749;
wire n_3962;
wire n_1826;
wire n_2304;
wire n_1283;
wire n_5325;
wire n_2637;
wire n_4384;
wire n_4423;
wire n_4096;
wire n_2881;
wire n_3282;
wire n_1763;
wire n_3231;
wire n_1966;
wire n_4996;
wire n_2475;
wire n_4598;
wire n_5064;
wire n_4478;
wire n_2646;
wire n_1605;
wire n_5173;
wire n_3920;
wire n_4890;
wire n_5027;
wire n_3203;
wire n_3866;
wire n_2903;
wire n_3921;
wire n_4106;
wire n_3717;
wire n_2743;
wire n_2675;
wire n_1439;
wire n_3052;
wire n_5215;
wire n_3743;
wire n_1932;
wire n_4721;
wire n_1983;
wire n_4029;
wire n_1594;
wire n_3870;
wire n_4496;
wire n_3529;
wire n_1977;
wire n_2153;
wire n_4338;
wire n_3094;
wire n_2310;
wire n_3952;
wire n_2287;
wire n_2860;
wire n_2056;
wire n_1470;
wire n_1735;
wire n_2318;
wire n_2502;
wire n_2504;
wire n_4495;
wire n_4762;
wire n_2974;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_3442;
wire n_3998;
wire n_2285;
wire n_3147;
wire n_4141;
wire n_5121;
wire n_1824;
wire n_1917;
wire n_3386;
wire n_4107;
wire n_4667;
wire n_2325;
wire n_2446;
wire n_3488;
wire n_4547;
wire n_2893;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_4668;
wire n_4953;
wire n_3898;
wire n_1786;
wire n_5284;
wire n_4997;
wire n_5308;
wire n_4274;
wire n_2627;
wire n_4759;
wire n_1413;
wire n_4467;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_3552;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_2361;
wire n_1603;
wire n_1401;
wire n_4113;
wire n_1998;
wire n_4686;
wire n_3759;
wire n_4321;
wire n_4342;
wire n_2034;
wire n_3933;
wire n_3206;
wire n_3966;
wire n_5243;
wire n_1702;
wire n_5221;
wire n_4183;
wire n_4068;
wire n_4872;
wire n_4233;
wire n_3192;
wire n_3764;
wire n_4709;
wire n_5038;
wire n_5311;
wire n_2649;
wire n_1929;
wire n_2807;
wire n_2542;
wire n_2313;
wire n_3324;
wire n_3914;
wire n_4625;
wire n_2558;
wire n_2063;
wire n_3803;
wire n_3742;
wire n_2252;
wire n_4819;
wire n_1685;
wire n_1714;
wire n_1541;
wire n_2576;
wire n_4900;
wire n_3390;
wire n_1573;
wire n_3746;
wire n_2373;
wire n_1713;
wire n_3817;
wire n_2745;
wire n_1253;
wire n_1737;
wire n_2493;
wire n_4930;
wire n_5276;
wire n_5078;
wire n_4537;
wire n_2885;
wire n_5011;
wire n_3318;
wire n_4070;
wire n_4282;
wire n_3485;
wire n_4180;
wire n_3839;
wire n_1440;
wire n_5205;
wire n_3333;
wire n_2845;
wire n_4143;
wire n_4659;
wire n_2602;
wire n_4579;
wire n_4616;
wire n_1496;
wire n_3014;
wire n_2547;
wire n_5023;
wire n_1812;
wire n_4105;
wire n_2532;
wire n_3791;
wire n_2665;
wire n_5351;
wire n_3905;
wire n_3368;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_3329;
wire n_2994;
wire n_2401;
wire n_3135;
wire n_2003;
wire n_1457;
wire n_4895;
wire n_3573;
wire n_3148;
wire n_2264;
wire n_3534;
wire n_1482;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_3438;
wire n_4098;
wire n_1297;
wire n_4789;
wire n_1972;
wire n_2806;
wire n_2184;
wire n_5312;
wire n_3217;
wire n_3404;
wire n_3425;
wire n_5111;
wire n_4055;
wire n_2926;
wire n_3540;
wire n_3670;
wire n_3973;
wire n_2023;
wire n_3249;
wire n_2351;
wire n_5113;
wire n_4442;
wire n_4698;
wire n_1602;
wire n_4779;
wire n_2286;
wire n_4966;
wire n_2065;
wire n_4017;
wire n_3397;
wire n_3740;
wire n_4418;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_1318;
wire n_2977;
wire n_1454;
wire n_3723;
wire n_3600;
wire n_4134;
wire n_1388;
wire n_2836;
wire n_1625;
wire n_2130;
wire n_5167;
wire n_3239;
wire n_5117;
wire n_2773;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_4913;
wire n_1452;
wire n_1791;
wire n_2850;
wire n_1747;
wire n_4251;
wire n_1817;
wire n_3982;
wire n_2654;
wire n_4621;
wire n_1326;
wire n_3176;
wire n_4559;
wire n_2186;
wire n_4368;
wire n_4740;
wire n_5301;
wire n_5007;
wire n_3581;
wire n_2562;
wire n_4077;
wire n_4642;
wire n_2221;
wire n_3576;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_4049;
wire n_3862;
wire n_5214;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_4724;
wire n_1772;
wire n_1476;
wire n_2818;
wire n_3646;
wire n_2129;
wire n_3345;
wire n_1395;
wire n_4546;
wire n_3584;
wire n_3756;
wire n_2889;
wire n_5021;
wire n_2772;
wire n_1675;
wire n_1924;
wire n_4382;
wire n_1554;
wire n_3999;
wire n_2844;
wire n_2138;
wire n_5211;
wire n_5230;
wire n_2260;
wire n_1813;
wire n_4833;
wire n_3056;
wire n_2345;
wire n_5110;
wire n_1341;
wire n_3295;
wire n_2382;
wire n_4719;
wire n_4178;
wire n_3062;
wire n_2317;
wire n_3289;
wire n_1973;
wire n_2579;
wire n_1770;
wire n_4228;
wire n_4401;
wire n_1756;
wire n_1716;
wire n_2788;
wire n_2984;
wire n_3364;
wire n_1873;
wire n_3201;
wire n_3472;
wire n_2874;
wire n_5179;
wire n_4605;
wire n_4877;
wire n_3235;
wire n_4968;
wire n_1272;
wire n_5030;
wire n_3949;
wire n_3543;
wire n_3050;
wire n_1478;
wire n_3903;
wire n_4834;
wire n_1364;
wire n_5272;
wire n_2183;
wire n_2742;
wire n_3314;
wire n_4158;
wire n_2360;
wire n_3254;
wire n_5361;
wire n_4171;
wire n_4045;
wire n_1367;
wire n_4562;
wire n_5068;
wire n_3634;
wire n_1460;
wire n_2834;
wire n_2531;
wire n_5015;
wire n_2702;
wire n_2030;
wire n_3115;
wire n_4749;
wire n_4390;
wire n_5302;
wire n_4979;
wire n_1404;
wire n_1794;
wire n_2234;
wire n_4804;
wire n_2209;
wire n_4270;
wire n_2797;
wire n_1255;
wire n_5152;
wire n_2321;
wire n_3680;
wire n_3497;
wire n_1601;
wire n_2940;
wire n_2612;
wire n_1495;
wire n_5128;
wire n_4566;
wire n_2841;
wire n_3322;
wire n_4576;
wire n_2427;
wire n_2505;
wire n_4061;
wire n_2070;
wire n_3250;
wire n_2594;
wire n_1914;
wire n_2335;
wire n_2904;
wire n_5307;
wire n_4767;
wire n_4328;
wire n_3004;
wire n_3112;
wire n_2349;
wire n_1379;
wire n_3874;
wire n_4676;
wire n_4544;
wire n_2170;
wire n_3175;
wire n_3522;
wire n_4429;
wire n_4591;
wire n_3266;
wire n_4646;
wire n_4563;
wire n_4725;
wire n_2210;
wire n_4169;
wire n_5331;
wire n_3247;
wire n_3091;
wire n_3066;
wire n_2426;
wire n_4320;
wire n_5341;
wire n_4881;
wire n_5271;
wire n_5089;
wire n_5263;
wire n_3613;
wire n_3444;
wire n_1505;
wire n_4012;
wire n_4636;
wire n_4584;
wire n_3910;
wire n_4711;
wire n_3319;
wire n_5240;
wire n_3335;
wire n_3413;
wire n_1969;
wire n_4680;
wire n_2044;
wire n_2689;
wire n_3259;
wire n_4191;
wire n_5224;
wire n_4293;
wire n_2010;
wire n_3688;
wire n_3016;
wire n_1693;
wire n_2599;
wire n_3338;
wire n_3414;
wire n_1827;
wire n_4671;
wire n_4209;
wire n_1271;
wire n_1542;
wire n_5041;
wire n_1423;
wire n_1751;
wire n_1508;
wire n_2200;
wire n_3261;
wire n_5026;
wire n_3863;
wire n_3027;
wire n_2746;
wire n_5059;
wire n_3127;
wire n_1780;
wire n_3732;
wire n_4250;
wire n_5329;
wire n_3596;
wire n_4699;
wire n_3906;
wire n_4127;
wire n_3297;
wire n_2683;
wire n_1370;
wire n_1360;
wire n_2388;
wire n_4292;
wire n_3641;
wire n_4577;
wire n_4854;
wire n_4202;
wire n_5212;
wire n_5000;
wire n_2853;
wire n_1323;
wire n_3766;
wire n_1353;
wire n_2880;
wire n_3350;
wire n_1666;
wire n_2389;
wire n_4165;
wire n_4866;
wire n_4038;
wire n_4109;
wire n_5297;
wire n_1264;
wire n_4412;
wire n_3407;
wire n_3599;
wire n_3621;
wire n_1580;
wire n_5234;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_1607;
wire n_2538;
wire n_2105;
wire n_5259;
wire n_3163;
wire n_1686;
wire n_3710;
wire n_4155;
wire n_1359;
wire n_2031;
wire n_3891;
wire n_4144;
wire n_2165;
wire n_3379;
wire n_4374;
wire n_3532;
wire n_5131;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_1294;
wire n_1257;
wire n_3531;
wire n_2963;
wire n_3834;
wire n_4548;
wire n_3258;
wire n_4989;
wire n_4622;
wire n_4315;
wire n_2959;
wire n_2047;
wire n_1845;
wire n_2193;
wire n_2478;
wire n_5140;
wire n_4816;
wire n_1483;
wire n_2983;
wire n_3810;
wire n_1289;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_5306;
wire n_4483;
wire n_5342;
wire n_2782;
wire n_2672;
wire n_1670;
wire n_2651;
wire n_4358;
wire n_5147;
wire n_3656;
wire n_2071;
wire n_2561;
wire n_2643;
wire n_1374;
wire n_4793;
wire n_4168;
wire n_3446;
wire n_3028;
wire n_4806;
wire n_4350;
wire n_5280;
wire n_1428;
wire n_5235;
wire n_3836;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1931;
wire n_4187;
wire n_4166;
wire n_5206;
wire n_3222;
wire n_1267;
wire n_1801;
wire n_1513;
wire n_2970;
wire n_2235;
wire n_4937;
wire n_3980;
wire n_2791;
wire n_5103;
wire n_1473;
wire n_3755;
wire n_4258;
wire n_4498;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_5285;
wire n_3563;
wire n_2506;
wire n_4064;
wire n_4936;
wire n_1556;
wire n_1863;
wire n_3841;
wire n_2118;
wire n_4770;
wire n_2944;
wire n_2407;
wire n_4907;
wire n_5058;
wire n_3262;
wire n_1450;
wire n_5018;
wire n_4006;
wire n_4861;
wire n_1322;
wire n_3690;
wire n_2358;
wire n_5192;
wire n_5141;
wire n_3716;
wire n_5133;
wire n_1700;
wire n_2833;
wire n_4712;
wire n_3191;
wire n_3837;
wire n_3193;
wire n_1971;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3273;
wire n_3544;
wire n_4310;
wire n_1523;
wire n_1950;
wire n_1447;
wire n_2370;
wire n_5159;
wire n_3954;
wire n_3025;
wire n_4674;
wire n_4908;
wire n_5097;
wire n_2750;
wire n_3899;
wire n_1278;
wire n_4159;
wire n_3714;
wire n_3071;
wire n_3739;
wire n_4069;
wire n_2784;
wire n_3718;
wire n_3092;
wire n_3470;
wire n_4862;
wire n_2557;
wire n_5300;
wire n_4850;
wire n_3781;
wire n_4813;
wire n_4912;
wire n_2590;
wire n_2330;
wire n_2942;
wire n_3106;
wire n_1882;
wire n_3328;
wire n_3889;
wire n_4256;
wire n_4224;
wire n_3508;
wire n_4024;
wire n_2218;
wire n_2267;
wire n_2636;
wire n_1951;
wire n_1825;
wire n_1883;
wire n_2759;
wire n_4415;
wire n_4702;
wire n_4252;
wire n_4457;
wire n_5139;
wire n_1393;
wire n_2319;
wire n_3481;
wire n_2808;
wire n_2679;
wire n_2676;
wire n_1709;
wire n_4491;
wire n_2930;
wire n_1838;
wire n_3514;
wire n_2777;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_2611;
wire n_4261;
wire n_1660;
wire n_4886;
wire n_4090;
wire n_2529;
wire n_2698;
wire n_5043;
wire n_1662;
wire n_1481;
wire n_4001;
wire n_3047;
wire n_2454;
wire n_4371;
wire n_5281;
wire n_4473;
wire n_3120;
wire n_4007;
wire n_1743;
wire n_4268;
wire n_5048;
wire n_5028;
wire n_1479;
wire n_4480;
wire n_2350;
wire n_3895;
wire n_4194;
wire n_4824;
wire n_1892;
wire n_4120;
wire n_4427;
wire n_3745;
wire n_2990;
wire n_1766;
wire n_1571;
wire n_3119;
wire n_4142;
wire n_4082;
wire n_3479;
wire n_4085;
wire n_4073;
wire n_4260;
wire n_1649;
wire n_4163;
wire n_4439;
wire n_2064;
wire n_3867;
wire n_4372;
wire n_3500;
wire n_3279;
wire n_2621;
wire n_5073;
wire n_5024;
wire n_1537;
wire n_4262;
wire n_2671;
wire n_1798;
wire n_1790;
wire n_4720;
wire n_1647;
wire n_4685;
wire n_2563;
wire n_2387;
wire n_4334;
wire n_1674;
wire n_1830;
wire n_2073;
wire n_4511;
wire n_4014;
wire n_5250;
wire n_3144;
wire n_4757;
wire n_2913;
wire n_2336;
wire n_1615;
wire n_4175;
wire n_2005;
wire n_1916;
wire n_4648;
wire n_1333;
wire n_5006;
wire n_1443;
wire n_1539;
wire n_4892;
wire n_3823;
wire n_1866;
wire n_4173;
wire n_1624;
wire n_4970;
wire n_3816;
wire n_1279;
wire n_4108;
wire n_4486;
wire n_2960;
wire n_4627;
wire n_2290;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_2040;
wire n_3199;
wire n_3843;
wire n_2145;
wire n_1639;
wire n_3030;
wire n_2580;
wire n_3685;
wire n_4249;
wire n_5163;
wire n_2039;
wire n_4961;
wire n_3753;
wire n_2035;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_5190;
wire n_2509;
wire n_3236;
wire n_4317;
wire n_1362;
wire n_4855;
wire n_3969;
wire n_2459;
wire n_4154;
wire n_3396;
wire n_1445;
wire n_4023;
wire n_4420;
wire n_1923;
wire n_5138;
wire n_2116;
wire n_1434;
wire n_1828;
wire n_2320;
wire n_5349;
wire n_2038;
wire n_2137;
wire n_4973;
wire n_4640;
wire n_2583;
wire n_4396;
wire n_5127;
wire n_4367;
wire n_2087;
wire n_5216;
wire n_1989;
wire n_3818;
wire n_2523;
wire n_4387;
wire n_4951;
wire n_4453;
wire n_4170;
wire n_1578;
wire n_3719;
wire n_1959;
wire n_3681;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_4308;
wire n_2812;
wire n_2355;
wire n_2133;
wire n_1426;
wire n_3830;
wire n_2585;
wire n_2725;
wire n_5175;
wire n_3883;
wire n_1355;
wire n_2565;
wire n_4152;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_3268;
wire n_4281;
wire n_4661;
wire n_4200;
wire n_3614;
wire n_2111;
wire n_3301;
wire n_3466;
wire n_4962;
wire n_2595;
wire n_3411;
wire n_4958;
wire n_4271;
wire n_5171;
wire n_3586;
wire n_1390;
wire n_4071;
wire n_4921;
wire n_1980;
wire n_3065;
wire n_4361;
wire n_4614;
wire n_1265;
wire n_2681;
wire n_3103;
wire n_4945;
wire n_2424;
wire n_4922;
wire n_4732;
wire n_1651;
wire n_2775;
wire n_4693;
wire n_4326;
wire n_3557;
wire n_2230;
wire n_4744;
wire n_2851;
wire n_4305;
wire n_1455;
wire n_2490;
wire n_1407;
wire n_4213;
wire n_2849;
wire n_3692;
wire n_2204;
wire n_4929;
wire n_1961;
wire n_4964;
wire n_1430;
wire n_4802;
wire n_1354;
wire n_4139;
wire n_3029;
wire n_2508;
wire n_4031;
wire n_2416;
wire n_3881;
wire n_2461;
wire n_2243;
wire n_4583;
wire n_4210;
wire n_5245;
wire n_4666;
wire n_2929;
wire n_3751;
wire n_2555;
wire n_2662;
wire n_1611;
wire n_2368;
wire n_2890;
wire n_2554;
wire n_3698;
wire n_3927;
wire n_1840;
wire n_4540;
wire n_3961;
wire n_1630;
wire n_4891;
wire n_3559;
wire n_2661;
wire n_2572;
wire n_3993;
wire n_4940;
wire n_5208;
wire n_3588;
wire n_2308;
wire n_4590;
wire n_4830;
wire n_5231;
wire n_5237;
wire n_4664;
wire n_3860;
wire n_3160;
wire n_2191;
wire n_5093;
wire n_2428;
wire n_3847;
wire n_4946;
wire n_1346;
wire n_4906;
wire n_2158;
wire n_3290;
wire n_4663;
wire n_5347;
wire n_2824;
wire n_3033;
wire n_3298;
wire n_2440;
wire n_4883;
wire n_1386;
wire n_2923;
wire n_1442;
wire n_4162;
wire n_3665;
wire n_5115;
wire n_3264;
wire n_2333;
wire n_2916;
wire n_4297;
wire n_1632;
wire n_3800;
wire n_2403;
wire n_4608;
wire n_5232;
wire n_2792;
wire n_2870;
wire n_3991;
wire n_3134;
wire n_4172;
wire n_4791;
wire n_4536;
wire n_5149;
wire n_2463;
wire n_5151;
wire n_4773;
wire n_5345;
wire n_5357;
wire n_4497;
wire n_2472;
wire n_4611;
wire n_4755;
wire n_1768;
wire n_2294;
wire n_4960;
wire n_2993;
wire n_1719;
wire n_3864;
wire n_4658;
wire n_5135;
wire n_2732;
wire n_2309;
wire n_2948;
wire n_1560;
wire n_4362;
wire n_4306;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2685;
wire n_2037;
wire n_1953;
wire n_4422;
wire n_2589;
wire n_1363;
wire n_1301;
wire n_3482;
wire n_2233;
wire n_1312;
wire n_4555;
wire n_2827;
wire n_5136;
wire n_5228;
wire n_1504;
wire n_3956;
wire n_5323;
wire n_3572;
wire n_4215;
wire n_4280;
wire n_3375;
wire n_4047;
wire n_2082;
wire n_1643;
wire n_3167;
wire n_5350;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_5338;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3854;
wire n_2468;
wire n_1610;
wire n_1422;
wire n_3078;
wire n_3253;
wire n_4027;
wire n_2280;
wire n_4599;
wire n_3363;
wire n_4812;
wire n_1511;
wire n_3689;
wire n_2020;
wire n_4628;
wire n_1881;
wire n_2749;
wire n_3451;
wire n_4873;
wire n_4657;
wire n_2971;
wire n_2311;
wire n_3950;
wire n_4458;
wire n_4121;
wire n_1616;
wire n_5090;
wire n_4476;
wire n_2298;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_5104;
wire n_5042;
wire n_4860;
wire n_4359;
wire n_2303;
wire n_2810;
wire n_2747;
wire n_1848;
wire n_2126;
wire n_4573;
wire n_5289;
wire n_4118;
wire n_4803;
wire n_4079;
wire n_4091;
wire n_1638;
wire n_2002;
wire n_5145;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_5132;
wire n_5191;
wire n_3085;
wire n_1655;
wire n_5359;
wire n_2574;
wire n_5293;
wire n_1358;
wire n_4316;
wire n_3697;
wire n_2638;
wire n_4044;
wire n_4062;
wire n_4524;
wire n_4843;
wire n_3971;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_2711;
wire n_5363;
wire n_5200;
wire n_1653;
wire n_1506;
wire n_2867;
wire n_1894;
wire n_2794;
wire n_3145;
wire n_3124;
wire n_4253;
wire n_5356;
wire n_5369;
wire n_2608;
wire n_5258;
wire n_2657;
wire n_5255;
wire n_2852;
wire n_2392;
wire n_3517;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_1834;
wire n_3758;
wire n_3356;
wire n_2835;
wire n_1572;
wire n_1968;
wire n_3269;
wire n_5080;
wire n_1516;
wire n_3506;
wire n_1736;
wire n_3605;
wire n_2409;
wire n_3402;
wire n_5295;
wire n_4679;
wire n_4115;
wire n_4998;
wire n_2988;
wire n_1731;
wire n_1970;
wire n_2766;
wire n_2201;
wire n_2117;
wire n_4167;
wire n_1993;
wire n_5155;
wire n_3835;
wire n_2205;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_3967;
wire n_5016;
wire n_1912;
wire n_3401;
wire n_3226;
wire n_1410;
wire n_3902;
wire n_4730;
wire n_2779;
wire n_1584;
wire n_3654;
wire n_2164;
wire n_2115;
wire n_2232;
wire n_5327;
wire n_1302;
wire n_1774;
wire n_4713;
wire n_5137;
wire n_2811;
wire n_3348;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_4204;
wire n_5098;
wire n_1991;
wire n_2224;
wire n_1543;
wire n_4743;
wire n_3805;
wire n_3825;
wire n_3657;
wire n_4924;
wire n_3928;
wire n_4859;
wire n_2692;
wire n_2008;
wire n_4654;
wire n_4733;
wire n_3792;
wire n_4272;
wire n_3974;
wire n_3871;
wire n_1753;
wire n_2283;
wire n_3278;
wire n_1689;
wire n_4269;
wire n_4695;
wire n_1855;
wire n_3312;
wire n_1352;
wire n_2197;
wire n_2199;
wire n_5069;
wire n_3285;
wire n_3968;
wire n_5099;
wire n_2228;
wire n_4704;
wire n_4551;
wire n_5052;
wire n_2421;
wire n_2902;
wire n_4957;
wire n_2480;
wire n_2363;
wire n_4072;
wire n_4781;
wire n_3606;
wire n_5004;
wire n_2550;
wire n_4424;
wire n_3055;
wire n_3711;
wire n_3315;
wire n_3172;
wire n_3292;
wire n_4436;
wire n_3878;
wire n_4450;
wire n_3553;
wire n_4746;
wire n_1683;
wire n_1530;
wire n_3131;
wire n_5118;
wire n_5105;
wire n_1409;
wire n_3850;
wire n_4459;
wire n_1268;
wire n_2996;
wire n_1320;
wire n_4050;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_2102;
wire n_4853;
wire n_2422;
wire n_2239;
wire n_5256;
wire n_2950;
wire n_5220;
wire n_3852;
wire n_5178;
wire n_4520;
wire n_2057;
wire n_4008;
wire n_5077;
wire n_3858;
wire n_1901;
wire n_4502;
wire n_3032;
wire n_4851;
wire n_1330;
wire n_3072;
wire n_3081;
wire n_3313;
wire n_2710;
wire n_1745;
wire n_3924;
wire n_4571;
wire n_2006;
wire n_5314;
wire n_1618;
wire n_2343;
wire n_3439;
wire n_5049;
wire n_2535;
wire n_4205;
wire n_2726;
wire n_5277;
wire n_4723;
wire n_5176;
wire n_2799;
wire n_4454;
wire n_4229;
wire n_4739;
wire n_2376;
wire n_3017;
wire n_2456;
wire n_3904;
wire n_5150;
wire n_2678;
wire n_4838;
wire n_2872;
wire n_2451;
wire n_5075;
wire n_4879;
wire n_5051;
wire n_3926;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2854;
wire n_1701;
wire n_4181;
wire n_1550;
wire n_2764;
wire n_1498;
wire n_4225;
wire n_2567;
wire n_5142;
wire n_3102;
wire n_1648;
wire n_4153;
wire n_5156;
wire n_3627;
wire n_4300;
wire n_3551;
wire n_1769;
wire n_4783;
wire n_2964;
wire n_3769;
wire n_2673;
wire n_4530;
wire n_4267;
wire n_2292;
wire n_3865;
wire n_3859;
wire n_3722;
wire n_2442;
wire n_1943;
wire n_3117;
wire n_3428;
wire n_2961;
wire n_3351;
wire n_3527;
wire n_1396;
wire n_1348;
wire n_2883;
wire n_1752;
wire n_4182;
wire n_2912;
wire n_1315;
wire n_4825;
wire n_4440;
wire n_4549;
wire n_1910;
wire n_3955;
wire n_5120;
wire n_4565;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_4574;
wire n_4839;
wire n_5222;
wire n_4016;
wire n_3435;
wire n_3575;
wire n_1546;
wire n_4231;
wire n_3165;
wire n_4923;
wire n_3652;
wire n_4097;
wire n_4083;
wire n_1937;
wire n_4461;
wire n_3234;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_3916;
wire n_2569;
wire n_3556;
wire n_4101;
wire n_2196;
wire n_3591;
wire n_4273;
wire n_3024;
wire n_3512;
wire n_4939;
wire n_5169;
wire n_4389;
wire n_3930;
wire n_4448;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_2404;
wire n_2083;
wire n_2503;
wire n_1540;
wire n_1936;
wire n_2027;
wire n_2642;
wire n_2500;
wire n_1918;
wire n_4831;
wire n_2513;
wire n_2695;
wire n_3480;
wire n_3057;
wire n_3194;
wire n_2414;
wire n_1402;
wire n_3662;
wire n_4319;
wire n_2229;
wire n_1397;
wire n_4596;
wire n_2004;
wire n_3694;
wire n_2586;
wire n_4726;
wire n_1398;
wire n_1879;
wire n_4751;
wire n_4222;
wire n_2274;
wire n_2972;
wire n_3225;
wire n_4119;
wire n_3799;
wire n_4298;
wire n_5201;
wire n_4474;
wire n_5217;
wire n_2511;
wire n_1681;
wire n_3383;
wire n_3585;
wire n_2975;
wire n_5029;
wire n_2704;
wire n_4214;
wire n_5158;
wire n_4884;
wire n_4366;
wire n_1251;
wire n_4009;
wire n_4580;
wire n_1263;
wire n_4129;
wire n_4871;
wire n_2617;
wire n_4999;
wire n_1859;
wire n_1677;
wire n_2955;
wire n_4112;
wire n_4337;
wire n_4138;
wire n_1528;
wire n_5335;
wire n_1292;
wire n_2520;
wire n_2134;
wire n_4236;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_5002;
wire n_3595;
wire n_1347;
wire n_5143;
wire n_4238;
wire n_1451;
wire n_2374;
wire n_1545;
wire n_1947;
wire n_2114;
wire n_3571;
wire n_2396;
wire n_1799;
wire n_4734;
wire n_1939;
wire n_2486;
wire n_4635;
wire n_3501;
wire n_1869;
wire n_4013;
wire n_3039;
wire n_2011;
wire n_4242;
wire n_4984;
wire n_3851;
wire n_2543;
wire n_3036;
wire n_1896;
wire n_3180;
wire n_5283;
wire n_5268;
wire n_1705;
wire n_4561;
wire n_2639;
wire n_3325;
wire n_3107;
wire n_4021;
wire n_3880;
wire n_5122;
wire n_1261;
wire n_3186;
wire n_4955;
wire n_4501;
wire n_3696;
wire n_1280;
wire n_3650;
wire n_2761;
wire n_3157;
wire n_2537;
wire n_2144;
wire n_2515;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_5330;
wire n_4197;
wire n_4829;
wire n_1949;
wire n_1946;
wire n_2936;
wire n_1484;
wire n_1328;
wire n_4715;
wire n_5039;
wire n_2141;
wire n_4369;
wire n_4543;
wire n_2099;
wire n_4941;
wire n_1831;
wire n_1598;
wire n_4394;
wire n_1850;
wire n_1749;
wire n_3101;
wire n_3669;
wire n_5278;
wire n_2663;
wire n_1394;
wire n_2693;
wire n_3798;
wire n_4065;
wire n_5187;
wire n_4944;
wire n_2180;
wire n_2249;
wire n_4135;
wire n_2632;
wire n_1547;
wire n_1755;
wire n_2908;
wire n_3744;
wire n_4263;
wire n_1862;
wire n_2915;
wire n_2300;
wire n_3291;
wire n_4716;
wire n_4942;
wire n_2432;
wire n_1521;
wire n_3405;
wire n_4745;
wire n_2337;
wire n_1384;
wire n_3907;
wire n_5344;
wire n_4629;
wire n_2932;
wire n_2980;
wire n_5225;
wire n_3306;
wire n_1784;
wire n_4857;
wire n_3136;
wire n_4080;
wire n_4226;
wire n_4741;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_4752;
wire n_5265;
wire n_1750;
wire n_1459;
wire n_3986;
wire n_4376;
wire n_4753;
wire n_4552;
wire n_3885;
wire n_2713;
wire n_5196;
wire n_5181;
wire n_2644;
wire n_2951;
wire n_3008;
wire n_3709;
wire n_5126;
wire n_2214;
wire n_3427;
wire n_2055;
wire n_4067;
wire n_1403;
wire n_4042;
wire n_4176;
wire n_4385;
wire n_3320;
wire n_5009;
wire n_2688;
wire n_5368;
wire n_1463;
wire n_3651;
wire n_4333;
wire n_3359;
wire n_2865;
wire n_2706;
wire n_3676;
wire n_4375;
wire n_4788;
wire n_4717;
wire n_4986;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_4815;
wire n_4246;
wire n_3580;
wire n_2139;
wire n_4609;
wire n_5291;
wire n_5114;
wire n_2674;
wire n_1565;
wire n_4088;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_4462;
wire n_4472;
wire n_3433;
wire n_5288;
wire n_2305;
wire n_2450;
wire n_3447;
wire n_3305;
wire n_4151;
wire n_4148;
wire n_1712;
wire n_3528;
wire n_4373;
wire n_4934;
wire n_5218;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_4630;
wire n_4643;
wire n_4331;
wire n_3989;
wire n_4475;
wire n_4846;
wire n_3804;
wire n_4344;
wire n_3296;
wire n_1775;
wire n_1368;
wire n_2762;
wire n_4683;
wire n_5366;
wire n_1847;
wire n_2767;
wire n_2603;
wire n_3116;
wire n_1884;
wire n_3602;
wire n_2967;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_2195;
wire n_3923;
wire n_4696;
wire n_2626;
wire n_3441;
wire n_1978;
wire n_1544;
wire n_5086;
wire n_1629;
wire n_2801;
wire n_4011;
wire n_4905;
wire n_2763;
wire n_2825;
wire n_3643;
wire n_4876;
wire n_1997;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_4278;
wire n_1635;
wire n_4623;
wire n_4910;
wire n_2690;
wire n_4410;
wire n_3370;
wire n_2215;
wire n_5053;
wire n_1259;
wire n_4553;
wire n_3978;
wire n_4809;
wire n_5226;
wire n_1925;
wire n_3660;
wire n_1815;
wire n_2491;
wire n_1788;
wire n_5079;
wire n_3833;
wire n_1679;
wire n_4841;
wire n_2022;
wire n_3814;
wire n_1415;
wire n_2592;
wire n_2838;
wire n_4842;
wire n_4911;
wire n_4340;
wire n_3513;
wire n_3133;
wire n_4645;
wire n_2992;
wire n_3725;
wire n_1833;
wire n_4920;
wire n_4972;
wire n_2517;
wire n_3128;
wire n_2631;
wire n_2178;
wire n_1767;
wire n_1529;
wire n_2469;
wire n_3355;
wire n_2007;
wire n_3917;
wire n_3942;
wire n_2736;
wire n_3765;
wire n_3000;
wire n_1406;
wire n_3108;
wire n_3111;
wire n_1837;
wire n_1839;
wire n_4557;
wire n_5248;
wire n_4451;
wire n_2875;
wire n_1500;
wire n_3844;
wire n_3280;
wire n_4054;
wire n_3471;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_5160;
wire n_2741;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_1656;
wire n_3564;
wire n_3988;
wire n_3457;
wire n_1678;
wire n_4324;
wire n_4821;
wire n_1871;
wire n_3630;
wire n_3271;
wire n_4771;
wire n_4086;
wire n_2412;
wire n_4814;
wire n_2084;
wire n_1781;
wire n_3648;
wire n_3075;
wire n_3173;
wire n_5332;
wire n_5108;
wire n_4692;
wire n_3031;
wire n_3701;
wire n_1773;
wire n_3243;
wire n_2666;
wire n_3385;
wire n_2171;
wire n_4708;
wire n_2768;
wire n_2314;
wire n_4826;
wire n_2420;
wire n_3343;
wire n_1593;
wire n_3767;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_4589;
wire n_5057;
wire n_4578;
wire n_1640;
wire n_2162;
wire n_2847;
wire n_2051;
wire n_3221;
wire n_2168;
wire n_2790;
wire n_5072;
wire n_3629;
wire n_3021;
wire n_2359;
wire n_3674;
wire n_5286;
wire n_3502;
wire n_3098;
wire n_1383;
wire n_5013;
wire n_2312;
wire n_3015;
wire n_1920;
wire n_4147;
wire n_2048;
wire n_3607;
wire n_4925;
wire n_1921;
wire n_1309;
wire n_4974;
wire n_1800;
wire n_1548;
wire n_4932;
wire n_1421;
wire n_4510;
wire n_2571;
wire n_1286;
wire n_3276;
wire n_3787;
wire n_5119;
wire n_2124;
wire n_3827;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_4447;
wire n_4285;
wire n_4651;
wire n_4818;
wire n_4514;
wire n_1366;
wire n_4800;
wire n_3960;
wire n_3248;
wire n_2277;
wire n_1568;
wire n_2110;
wire n_1332;
wire n_4433;
wire n_2879;
wire n_2474;
wire n_2090;
wire n_3153;
wire n_1591;
wire n_2033;
wire n_4341;
wire n_1682;
wire n_4312;
wire n_2628;
wire n_3399;
wire n_1249;
wire n_2132;
wire n_2400;
wire n_4633;
wire n_3838;
wire n_1909;
wire n_4277;
wire n_4140;
wire n_3675;
wire n_5092;
wire n_3387;
wire n_5186;
wire n_4662;
wire n_3779;
wire n_2464;
wire n_2831;
wire n_1456;
wire n_4882;
wire n_4993;
wire n_2365;
wire n_4832;
wire n_4207;
wire n_4545;
wire n_3037;
wire n_4868;
wire n_1885;
wire n_2452;
wire n_3925;
wire n_2176;
wire n_1816;
wire n_5238;
wire n_4059;
wire n_2455;
wire n_4595;
wire n_1849;
wire n_5054;
wire n_2467;
wire n_2288;
wire n_4063;
wire n_3592;
wire n_4650;
wire n_4888;
wire n_5326;
wire n_1435;
wire n_3394;
wire n_4874;
wire n_3793;
wire n_4669;
wire n_4339;
wire n_1645;
wire n_4041;
wire n_2858;
wire n_4060;
wire n_2658;
wire n_1717;
wire n_2895;
wire n_2128;
wire n_3097;
wire n_4541;
wire n_3824;
wire n_3388;
wire n_5267;
wire n_4494;
wire n_3059;
wire n_3465;
wire n_1316;
wire n_4796;
wire n_1438;
wire n_3589;
wire n_2534;
wire n_4799;
wire n_5153;
wire n_3449;
wire n_2694;
wire n_2198;
wire n_2610;
wire n_2989;
wire n_2789;
wire n_4775;
wire n_2216;
wire n_5044;
wire n_1897;
wire n_1424;
wire n_5365;
wire n_2933;
wire n_5045;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_5354;
wire n_4455;
wire n_2328;
wire n_4248;
wire n_4754;
wire n_4554;
wire n_4845;
wire n_3053;
wire n_1299;
wire n_3893;
wire n_2465;
wire n_3548;
wire n_4585;
wire n_1699;
wire n_3334;
wire n_2541;
wire n_4383;
wire n_1432;
wire n_3875;
wire n_5370;
wire n_4003;
wire n_5299;
wire n_2402;
wire n_4301;
wire n_4586;
wire n_1954;
wire n_4048;
wire n_1844;
wire n_3777;
wire n_4784;
wire n_2999;
wire n_1644;
wire n_5082;
wire n_4046;
wire n_1974;
wire n_2086;
wire n_3537;
wire n_5209;
wire n_3080;
wire n_4199;
wire n_2701;
wire n_3362;
wire n_1631;
wire n_3105;
wire n_4286;
wire n_5102;
wire n_2556;
wire n_2269;
wire n_3274;
wire n_3041;
wire n_4470;
wire n_2236;
wire n_2816;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3664;
wire n_4188;
wire n_1668;
wire n_3913;
wire n_3417;
wire n_1579;
wire n_4034;
wire n_1688;
wire n_3327;
wire n_5275;
wire n_4689;
wire n_5071;
wire n_3067;
wire n_2755;
wire n_3237;
wire n_1992;
wire n_4402;
wire n_4239;
wire n_3400;
wire n_4550;
wire n_1342;
wire n_1400;
wire n_3382;
wire n_3574;
wire n_5227;
wire n_2169;
wire n_1557;
wire n_4201;
wire n_3316;
wire n_5242;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_1730;
wire n_3603;
wire n_4123;
wire n_2192;
wire n_3633;
wire n_4479;
wire n_1373;
wire n_2670;
wire n_1646;
wire n_1307;
wire n_4416;
wire n_3372;
wire n_4539;
wire n_2707;
wire n_2471;
wire n_1472;
wire n_1671;
wire n_3230;
wire n_3342;
wire n_4682;
wire n_5353;
wire n_3708;
wire n_5294;
wire n_3729;
wire n_4978;
wire n_4690;
wire n_4437;
wire n_3861;
wire n_4736;
wire n_3780;
wire n_1928;
wire n_5244;
wire n_3957;
wire n_5274;
wire n_3848;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_3608;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_3177;
wire n_4053;
wire n_2352;
wire n_5125;
wire n_4040;
wire n_2207;
wire n_2619;
wire n_2444;
wire n_3123;
wire n_5056;
wire n_5249;
wire n_3393;
wire n_5198;
wire n_5360;
wire n_5233;
wire n_4887;
wire n_4617;
wire n_5269;
wire n_3520;
wire n_2492;
wire n_4005;
wire n_1687;
wire n_1637;
wire n_4904;
wire n_1419;
wire n_4792;
wire n_3578;
wire n_3812;
wire n_1886;
wire n_1389;
wire n_1256;
wire n_4980;
wire n_1465;
wire n_4290;
wire n_5247;
wire n_1375;
wire n_3727;
wire n_5317;
wire n_3774;
wire n_3093;
wire n_1843;
wire n_3061;
wire n_1597;
wire n_1659;
wire n_2431;
wire n_1371;
wire n_4956;
wire n_2206;
wire n_3182;
wire n_2564;
wire n_4947;
wire n_4656;
wire n_3896;
wire n_3958;
wire n_3450;
wire n_4729;
wire n_4987;
wire n_5182;
wire n_4971;
wire n_2000;
wire n_2074;
wire n_3174;
wire n_2217;
wire n_1453;
wire n_3398;
wire n_2307;
wire n_3408;
wire n_2722;
wire n_2640;
wire n_4823;
wire n_4875;
wire n_3432;
wire n_1628;
wire n_1514;
wire n_1771;
wire n_3090;
wire n_2437;
wire n_3762;
wire n_2445;
wire n_1427;
wire n_1835;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_4137;
wire n_2634;
wire n_4529;
wire n_4323;
wire n_3034;
wire n_2212;
wire n_3972;
wire n_3308;
wire n_1533;
wire n_5036;
wire n_4772;
wire n_3467;
wire n_4322;
wire n_1720;
wire n_2830;
wire n_4354;
wire n_4653;
wire n_2354;
wire n_2246;
wire n_5273;
wire n_4677;
wire n_3901;
wire n_1480;
wire n_5261;
wire n_3757;
wire n_3381;
wire n_5193;
wire n_2245;
wire n_1782;
wire n_4909;
wire n_1524;
wire n_1485;
wire n_2965;
wire n_3635;
wire n_5022;
wire n_5005;
wire n_2814;
wire n_1570;
wire n_3882;
wire n_3046;
wire n_2213;
wire n_3826;
wire n_3211;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_4634;
wire n_3337;
wire n_2527;
wire n_1461;
wire n_3204;
wire n_2136;
wire n_5174;
wire n_1273;
wire n_1822;
wire n_4952;
wire n_5157;
wire n_3005;
wire n_4380;
wire n_3129;
wire n_4126;
wire n_1282;
wire n_1783;
wire n_2601;
wire n_5087;
wire n_3043;
wire n_3802;
wire n_2375;
wire n_4506;
wire n_4880;
wire n_1907;
wire n_2686;
wire n_2344;
wire n_3892;
wire n_4896;
wire n_1417;
wire n_1295;
wire n_5061;
wire n_1985;
wire n_2107;
wire n_3219;
wire n_2906;
wire n_4943;
wire n_2187;
wire n_1762;
wire n_3023;
wire n_4193;
wire n_4075;
wire n_3104;
wire n_4737;
wire n_3647;
wire n_2819;
wire n_5195;
wire n_3609;
wire n_4136;
wire n_1715;
wire n_1952;
wire n_4393;
wire n_3720;
wire n_4535;
wire n_1922;
wire n_2560;
wire n_4522;
wire n_4794;
wire n_3959;
wire n_3140;
wire n_5246;
wire n_3724;
wire n_2104;
wire n_3011;
wire n_5164;
wire n_4196;
wire n_1425;
wire n_4592;
wire n_4675;
wire n_5340;
wire n_3069;
wire n_4370;
wire n_1900;
wire n_1620;
wire n_5183;
wire n_3084;
wire n_1727;
wire n_2735;
wire n_2497;
wire n_3412;
wire n_1995;
wire n_2411;
wire n_3761;
wire n_4889;
wire n_2014;
wire n_2986;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_4828;
wire n_4558;
wire n_2172;
wire n_4722;
wire n_3626;
wire n_4768;
wire n_4100;
wire n_2250;
wire n_4092;
wire n_3908;
wire n_2423;
wire n_3671;
wire n_3344;
wire n_2194;
wire n_4465;
wire n_3302;
wire n_5304;
wire n_2680;
wire n_5130;
wire n_1567;
wire n_3122;
wire n_5162;
wire n_4808;
wire n_3842;
wire n_3265;
wire n_1857;
wire n_4482;
wire n_2041;
wire n_1797;
wire n_2957;
wire n_2357;
wire n_1250;
wire n_3309;
wire n_3260;
wire n_4926;
wire n_3357;
wire n_1589;
wire n_4116;
wire n_2570;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_3754;
wire n_4612;
wire n_1469;
wire n_2744;
wire n_4287;
wire n_2397;
wire n_2208;
wire n_3063;
wire n_5177;
wire n_3617;
wire n_1298;
wire n_1652;
wire n_4516;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_4505;
wire n_1676;
wire n_1277;
wire n_2591;
wire n_3384;
wire n_4602;
wire n_5172;
wire n_4449;
wire n_1864;
wire n_5070;
wire n_1337;
wire n_4445;
wire n_1627;
wire n_4870;
wire n_2438;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_3181;
wire n_2278;
wire n_4915;
wire n_5296;
wire n_2135;
wire n_3493;
wire n_5313;
wire n_3323;
wire n_2734;
wire n_4914;
wire n_2823;
wire n_1408;
wire n_1761;
wire n_5270;
wire n_4345;
wire n_5188;
wire n_3281;
wire n_3307;
wire n_1606;
wire n_1694;
wire n_4318;
wire n_2485;
wire n_2655;
wire n_4185;
wire n_4797;
wire n_2366;
wire n_1526;
wire n_3997;
wire n_1604;
wire n_1275;
wire n_4032;
wire n_1764;
wire n_3582;
wire n_1583;
wire n_2826;
wire n_3539;
wire n_4343;
wire n_1493;
wire n_4212;
wire n_4124;
wire n_4492;
wire n_2708;
wire n_5148;
wire n_4994;
wire n_4245;
wire n_4364;
wire n_4928;
wire n_2225;
wire n_1507;
wire n_4378;
wire n_2383;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_3853;
wire n_4216;
wire n_2019;
wire n_1340;
wire n_1558;
wire n_2166;
wire n_2938;
wire n_4309;
wire n_3594;
wire n_1704;
wire n_3721;
wire n_1254;
wire n_2026;
wire n_2109;
wire n_2013;
wire n_1990;
wire n_2614;
wire n_2991;
wire n_2242;
wire n_2752;
wire n_2894;
wire n_3473;
wire n_4560;
wire n_5318;
wire n_2839;
wire n_1588;
wire n_2237;
wire n_3463;
wire n_3699;
wire n_5067;
wire n_3360;
wire n_2524;
wire n_3873;
wire n_3693;
wire n_2728;
wire n_3857;

INVx1_ASAP7_75t_L g1249 ( 
.A(n_220),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_613),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_1110),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1194),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_1182),
.Y(n_1253)
);

INVx2_ASAP7_75t_SL g1254 ( 
.A(n_188),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1005),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_374),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1205),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_949),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1096),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_757),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_76),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_480),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_246),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_480),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_349),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_554),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_763),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_452),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_216),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_807),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_260),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1075),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_1216),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_1044),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_27),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_160),
.Y(n_1276)
);

BUFx5_ASAP7_75t_L g1277 ( 
.A(n_583),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_575),
.Y(n_1278)
);

INVx2_ASAP7_75t_SL g1279 ( 
.A(n_481),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1015),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_335),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_702),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_955),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_1125),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1242),
.Y(n_1285)
);

CKINVDCx16_ASAP7_75t_R g1286 ( 
.A(n_287),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1074),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_809),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_1025),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_718),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1046),
.Y(n_1291)
);

BUFx10_ASAP7_75t_L g1292 ( 
.A(n_677),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_72),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_266),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1137),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1163),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1080),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_1141),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_984),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_505),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_554),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1162),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1231),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1128),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_168),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_354),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_132),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1209),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_1212),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_957),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_188),
.Y(n_1311)
);

CKINVDCx14_ASAP7_75t_R g1312 ( 
.A(n_935),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_916),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_44),
.Y(n_1314)
);

CKINVDCx14_ASAP7_75t_R g1315 ( 
.A(n_264),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_161),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_672),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_474),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_580),
.Y(n_1319)
);

BUFx5_ASAP7_75t_L g1320 ( 
.A(n_1201),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_1109),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1052),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1090),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_1179),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1244),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_498),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1225),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1183),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_937),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_1121),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_1131),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_1136),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_579),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1007),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_911),
.Y(n_1335)
);

BUFx5_ASAP7_75t_L g1336 ( 
.A(n_1053),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_922),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1146),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_934),
.Y(n_1339)
);

INVx1_ASAP7_75t_SL g1340 ( 
.A(n_661),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_920),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1189),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_760),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_616),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1185),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_1239),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_238),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_828),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1026),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_1145),
.Y(n_1350)
);

CKINVDCx16_ASAP7_75t_R g1351 ( 
.A(n_1199),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1060),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_943),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1172),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_556),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_742),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_544),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_632),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1035),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_942),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1228),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_123),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_35),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_946),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_39),
.Y(n_1365)
);

BUFx8_ASAP7_75t_SL g1366 ( 
.A(n_1048),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1222),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1023),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_252),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_380),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1036),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_167),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_54),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_331),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_147),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_526),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_24),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_121),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_737),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_891),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_1029),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1012),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_427),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_833),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_695),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_220),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1119),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1157),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_265),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1215),
.Y(n_1390)
);

CKINVDCx20_ASAP7_75t_R g1391 ( 
.A(n_615),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_451),
.Y(n_1392)
);

CKINVDCx14_ASAP7_75t_R g1393 ( 
.A(n_1021),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_816),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_294),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_719),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_366),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_260),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_219),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_954),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_952),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_440),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_914),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_671),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1106),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_1057),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_567),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1129),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_832),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_679),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_498),
.Y(n_1411)
);

CKINVDCx12_ASAP7_75t_R g1412 ( 
.A(n_1120),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1169),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_444),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_33),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1031),
.Y(n_1416)
);

BUFx5_ASAP7_75t_L g1417 ( 
.A(n_5),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1115),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_538),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_488),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_943),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1186),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_1217),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_678),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1000),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1101),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_869),
.Y(n_1427)
);

BUFx6f_ASAP7_75t_L g1428 ( 
.A(n_1175),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1087),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1093),
.Y(n_1430)
);

BUFx6f_ASAP7_75t_L g1431 ( 
.A(n_1122),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_978),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1078),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_457),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_598),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1065),
.Y(n_1436)
);

INVx1_ASAP7_75t_SL g1437 ( 
.A(n_1192),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_1108),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1001),
.Y(n_1439)
);

CKINVDCx20_ASAP7_75t_R g1440 ( 
.A(n_1223),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1143),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1195),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_703),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1016),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1160),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_715),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_274),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1210),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_394),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1142),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_577),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_898),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1177),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_1170),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1140),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_682),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_496),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_314),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_103),
.Y(n_1459)
);

CKINVDCx20_ASAP7_75t_R g1460 ( 
.A(n_47),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_163),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_372),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_956),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_895),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_662),
.Y(n_1465)
);

CKINVDCx16_ASAP7_75t_R g1466 ( 
.A(n_523),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1155),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1095),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1245),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1117),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_913),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_44),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_618),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1059),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_571),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_790),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_744),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_750),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_242),
.Y(n_1479)
);

INVx2_ASAP7_75t_SL g1480 ( 
.A(n_2),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_1167),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_1126),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1113),
.Y(n_1483)
);

INVx2_ASAP7_75t_SL g1484 ( 
.A(n_941),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1127),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_124),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_578),
.Y(n_1487)
);

BUFx6f_ASAP7_75t_L g1488 ( 
.A(n_1105),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_98),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_458),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_538),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_467),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_388),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_393),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1236),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_342),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_1100),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_527),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_380),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_1041),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1220),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_529),
.Y(n_1502)
);

CKINVDCx20_ASAP7_75t_R g1503 ( 
.A(n_172),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1134),
.Y(n_1504)
);

CKINVDCx20_ASAP7_75t_R g1505 ( 
.A(n_859),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_167),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_987),
.Y(n_1507)
);

CKINVDCx20_ASAP7_75t_R g1508 ( 
.A(n_1247),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_252),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_189),
.Y(n_1510)
);

INVx1_ASAP7_75t_SL g1511 ( 
.A(n_562),
.Y(n_1511)
);

CKINVDCx16_ASAP7_75t_R g1512 ( 
.A(n_330),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_288),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_503),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_468),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_568),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_1040),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_908),
.Y(n_1518)
);

BUFx3_ASAP7_75t_L g1519 ( 
.A(n_192),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_514),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_942),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_899),
.Y(n_1522)
);

CKINVDCx20_ASAP7_75t_R g1523 ( 
.A(n_1181),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_457),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_202),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_135),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_985),
.Y(n_1527)
);

CKINVDCx16_ASAP7_75t_R g1528 ( 
.A(n_74),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_615),
.Y(n_1529)
);

INVx1_ASAP7_75t_SL g1530 ( 
.A(n_939),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_583),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_930),
.Y(n_1532)
);

INVx1_ASAP7_75t_SL g1533 ( 
.A(n_169),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_156),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_528),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1237),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_761),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_369),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_107),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1161),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_586),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_L g1542 ( 
.A(n_190),
.Y(n_1542)
);

CKINVDCx20_ASAP7_75t_R g1543 ( 
.A(n_816),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1028),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_193),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_712),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1148),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_729),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_105),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_300),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_917),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1203),
.Y(n_1552)
);

BUFx6f_ASAP7_75t_L g1553 ( 
.A(n_419),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_698),
.Y(n_1554)
);

INVx1_ASAP7_75t_SL g1555 ( 
.A(n_53),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_1056),
.Y(n_1556)
);

BUFx3_ASAP7_75t_L g1557 ( 
.A(n_931),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_321),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_628),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_131),
.Y(n_1560)
);

BUFx10_ASAP7_75t_L g1561 ( 
.A(n_938),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_19),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_977),
.Y(n_1563)
);

CKINVDCx20_ASAP7_75t_R g1564 ( 
.A(n_845),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_801),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_763),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_744),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_360),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_862),
.Y(n_1569)
);

INVxp67_ASAP7_75t_L g1570 ( 
.A(n_1099),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_L g1571 ( 
.A(n_1063),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_112),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1198),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_718),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1178),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_726),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1073),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_607),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_940),
.Y(n_1579)
);

CKINVDCx20_ASAP7_75t_R g1580 ( 
.A(n_1184),
.Y(n_1580)
);

CKINVDCx20_ASAP7_75t_R g1581 ( 
.A(n_548),
.Y(n_1581)
);

CKINVDCx16_ASAP7_75t_R g1582 ( 
.A(n_340),
.Y(n_1582)
);

INVxp67_ASAP7_75t_L g1583 ( 
.A(n_1039),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_504),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_850),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_134),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_493),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_524),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1214),
.Y(n_1589)
);

BUFx10_ASAP7_75t_L g1590 ( 
.A(n_1094),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_567),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_397),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1116),
.Y(n_1593)
);

CKINVDCx20_ASAP7_75t_R g1594 ( 
.A(n_1033),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_933),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1118),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_144),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_894),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_224),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_605),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_927),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_884),
.Y(n_1602)
);

CKINVDCx20_ASAP7_75t_R g1603 ( 
.A(n_1164),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_1227),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_671),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_596),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_1010),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1069),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1097),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_755),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_124),
.Y(n_1611)
);

CKINVDCx20_ASAP7_75t_R g1612 ( 
.A(n_1152),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_384),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_389),
.Y(n_1614)
);

CKINVDCx20_ASAP7_75t_R g1615 ( 
.A(n_155),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_555),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_289),
.Y(n_1617)
);

CKINVDCx16_ASAP7_75t_R g1618 ( 
.A(n_588),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_1149),
.Y(n_1619)
);

CKINVDCx20_ASAP7_75t_R g1620 ( 
.A(n_285),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_959),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_624),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_118),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_392),
.Y(n_1624)
);

BUFx10_ASAP7_75t_L g1625 ( 
.A(n_314),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_591),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_626),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_929),
.Y(n_1628)
);

CKINVDCx20_ASAP7_75t_R g1629 ( 
.A(n_205),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_963),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_975),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1076),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1081),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_449),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1079),
.Y(n_1635)
);

CKINVDCx20_ASAP7_75t_R g1636 ( 
.A(n_921),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_361),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_473),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_971),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1176),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_347),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_12),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1112),
.Y(n_1643)
);

BUFx3_ASAP7_75t_L g1644 ( 
.A(n_308),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_873),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_639),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_51),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_611),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1207),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_1138),
.Y(n_1650)
);

BUFx6f_ASAP7_75t_L g1651 ( 
.A(n_945),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_932),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_261),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_419),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_909),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_1018),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_105),
.Y(n_1657)
);

BUFx10_ASAP7_75t_L g1658 ( 
.A(n_1219),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_1088),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_1102),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_1173),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_33),
.Y(n_1662)
);

CKINVDCx20_ASAP7_75t_R g1663 ( 
.A(n_214),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1206),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1208),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_947),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_94),
.Y(n_1667)
);

BUFx6f_ASAP7_75t_L g1668 ( 
.A(n_398),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_817),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_9),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_919),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_791),
.Y(n_1672)
);

BUFx6f_ASAP7_75t_L g1673 ( 
.A(n_327),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_600),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_799),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_469),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1054),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_1022),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1133),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_73),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1229),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_269),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1055),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_1171),
.Y(n_1684)
);

INVxp67_ASAP7_75t_SL g1685 ( 
.A(n_134),
.Y(n_1685)
);

BUFx3_ASAP7_75t_L g1686 ( 
.A(n_910),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_557),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_1221),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_118),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_1006),
.Y(n_1690)
);

BUFx3_ASAP7_75t_L g1691 ( 
.A(n_910),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_1091),
.Y(n_1692)
);

INVx1_ASAP7_75t_SL g1693 ( 
.A(n_283),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_983),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_1211),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1240),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_965),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_948),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_354),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_805),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_879),
.Y(n_1701)
);

BUFx10_ASAP7_75t_L g1702 ( 
.A(n_1234),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1083),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_344),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_170),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_8),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_890),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_928),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_973),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_911),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_681),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_958),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_1034),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_918),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_1200),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_422),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_344),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_806),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_964),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_309),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_316),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_991),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_1049),
.Y(n_1723)
);

BUFx5_ASAP7_75t_L g1724 ( 
.A(n_365),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_470),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_334),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_993),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_82),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_862),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_836),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_559),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_590),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_1188),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_878),
.Y(n_1734)
);

BUFx3_ASAP7_75t_L g1735 ( 
.A(n_1191),
.Y(n_1735)
);

INVx1_ASAP7_75t_SL g1736 ( 
.A(n_1037),
.Y(n_1736)
);

INVx3_ASAP7_75t_L g1737 ( 
.A(n_164),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_646),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_1197),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_276),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_192),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_892),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_1248),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_604),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1086),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_445),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_946),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_1062),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_874),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_800),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_1224),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_648),
.Y(n_1752)
);

INVx2_ASAP7_75t_SL g1753 ( 
.A(n_904),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_514),
.Y(n_1754)
);

CKINVDCx20_ASAP7_75t_R g1755 ( 
.A(n_662),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_84),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_1061),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_914),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_1092),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_144),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_485),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_1003),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_937),
.Y(n_1763)
);

INVx1_ASAP7_75t_SL g1764 ( 
.A(n_76),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_399),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_403),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_834),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1165),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_944),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_893),
.Y(n_1770)
);

CKINVDCx20_ASAP7_75t_R g1771 ( 
.A(n_695),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_1156),
.Y(n_1772)
);

CKINVDCx20_ASAP7_75t_R g1773 ( 
.A(n_672),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_888),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_371),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_83),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_839),
.Y(n_1777)
);

CKINVDCx5p33_ASAP7_75t_R g1778 ( 
.A(n_846),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1089),
.Y(n_1779)
);

CKINVDCx20_ASAP7_75t_R g1780 ( 
.A(n_115),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_901),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_996),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_319),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_818),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_277),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_833),
.Y(n_1786)
);

CKINVDCx5p33_ASAP7_75t_R g1787 ( 
.A(n_1166),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_30),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_856),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_1002),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_876),
.Y(n_1791)
);

BUFx3_ASAP7_75t_L g1792 ( 
.A(n_84),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1174),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_524),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_229),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_281),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_1202),
.Y(n_1797)
);

CKINVDCx20_ASAP7_75t_R g1798 ( 
.A(n_1233),
.Y(n_1798)
);

CKINVDCx5p33_ASAP7_75t_R g1799 ( 
.A(n_902),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1180),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_3),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_1246),
.Y(n_1802)
);

CKINVDCx5p33_ASAP7_75t_R g1803 ( 
.A(n_540),
.Y(n_1803)
);

BUFx10_ASAP7_75t_L g1804 ( 
.A(n_373),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_1004),
.Y(n_1805)
);

BUFx5_ASAP7_75t_L g1806 ( 
.A(n_8),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_348),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_297),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_72),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_497),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1135),
.Y(n_1811)
);

CKINVDCx5p33_ASAP7_75t_R g1812 ( 
.A(n_635),
.Y(n_1812)
);

CKINVDCx5p33_ASAP7_75t_R g1813 ( 
.A(n_37),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_208),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_934),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_254),
.Y(n_1816)
);

CKINVDCx20_ASAP7_75t_R g1817 ( 
.A(n_728),
.Y(n_1817)
);

CKINVDCx16_ASAP7_75t_R g1818 ( 
.A(n_147),
.Y(n_1818)
);

BUFx3_ASAP7_75t_L g1819 ( 
.A(n_1124),
.Y(n_1819)
);

CKINVDCx20_ASAP7_75t_R g1820 ( 
.A(n_115),
.Y(n_1820)
);

CKINVDCx20_ASAP7_75t_R g1821 ( 
.A(n_267),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1027),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_309),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1123),
.Y(n_1824)
);

CKINVDCx5p33_ASAP7_75t_R g1825 ( 
.A(n_7),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_622),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_1038),
.Y(n_1827)
);

CKINVDCx20_ASAP7_75t_R g1828 ( 
.A(n_476),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_557),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_408),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_814),
.Y(n_1831)
);

INVx2_ASAP7_75t_SL g1832 ( 
.A(n_55),
.Y(n_1832)
);

CKINVDCx5p33_ASAP7_75t_R g1833 ( 
.A(n_1067),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_182),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_604),
.Y(n_1835)
);

CKINVDCx20_ASAP7_75t_R g1836 ( 
.A(n_660),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_723),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_951),
.Y(n_1838)
);

CKINVDCx5p33_ASAP7_75t_R g1839 ( 
.A(n_460),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_102),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_441),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_198),
.Y(n_1842)
);

BUFx3_ASAP7_75t_L g1843 ( 
.A(n_713),
.Y(n_1843)
);

CKINVDCx20_ASAP7_75t_R g1844 ( 
.A(n_1071),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_1235),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_801),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_925),
.Y(n_1847)
);

CKINVDCx5p33_ASAP7_75t_R g1848 ( 
.A(n_789),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_25),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_888),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_944),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_504),
.Y(n_1852)
);

INVx1_ASAP7_75t_SL g1853 ( 
.A(n_926),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1104),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_722),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1050),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_529),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_1098),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_585),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_1072),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_872),
.Y(n_1861)
);

CKINVDCx16_ASAP7_75t_R g1862 ( 
.A(n_1158),
.Y(n_1862)
);

BUFx6f_ASAP7_75t_L g1863 ( 
.A(n_454),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1153),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_212),
.Y(n_1865)
);

CKINVDCx5p33_ASAP7_75t_R g1866 ( 
.A(n_927),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_915),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1204),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1085),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_683),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_357),
.Y(n_1871)
);

BUFx3_ASAP7_75t_L g1872 ( 
.A(n_473),
.Y(n_1872)
);

CKINVDCx5p33_ASAP7_75t_R g1873 ( 
.A(n_1132),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_858),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_1238),
.Y(n_1875)
);

INVxp67_ASAP7_75t_L g1876 ( 
.A(n_1150),
.Y(n_1876)
);

CKINVDCx5p33_ASAP7_75t_R g1877 ( 
.A(n_1),
.Y(n_1877)
);

BUFx3_ASAP7_75t_L g1878 ( 
.A(n_999),
.Y(n_1878)
);

CKINVDCx16_ASAP7_75t_R g1879 ( 
.A(n_53),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_803),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_408),
.Y(n_1881)
);

BUFx6f_ASAP7_75t_L g1882 ( 
.A(n_364),
.Y(n_1882)
);

CKINVDCx20_ASAP7_75t_R g1883 ( 
.A(n_722),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_527),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_997),
.Y(n_1885)
);

CKINVDCx5p33_ASAP7_75t_R g1886 ( 
.A(n_1019),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_74),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_706),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1009),
.Y(n_1889)
);

CKINVDCx5p33_ASAP7_75t_R g1890 ( 
.A(n_614),
.Y(n_1890)
);

BUFx3_ASAP7_75t_L g1891 ( 
.A(n_1196),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_923),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_34),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_808),
.Y(n_1894)
);

BUFx10_ASAP7_75t_L g1895 ( 
.A(n_840),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_262),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_613),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_326),
.Y(n_1898)
);

INVx1_ASAP7_75t_SL g1899 ( 
.A(n_729),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_477),
.Y(n_1900)
);

BUFx6f_ASAP7_75t_L g1901 ( 
.A(n_1020),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_912),
.Y(n_1902)
);

CKINVDCx5p33_ASAP7_75t_R g1903 ( 
.A(n_820),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_343),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_533),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_273),
.Y(n_1906)
);

INVx2_ASAP7_75t_SL g1907 ( 
.A(n_692),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_123),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_924),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_979),
.Y(n_1910)
);

CKINVDCx5p33_ASAP7_75t_R g1911 ( 
.A(n_627),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_1230),
.Y(n_1912)
);

CKINVDCx5p33_ASAP7_75t_R g1913 ( 
.A(n_222),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_687),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_1064),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_302),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1213),
.Y(n_1917)
);

INVxp67_ASAP7_75t_L g1918 ( 
.A(n_1241),
.Y(n_1918)
);

CKINVDCx16_ASAP7_75t_R g1919 ( 
.A(n_630),
.Y(n_1919)
);

BUFx10_ASAP7_75t_L g1920 ( 
.A(n_741),
.Y(n_1920)
);

BUFx3_ASAP7_75t_L g1921 ( 
.A(n_552),
.Y(n_1921)
);

CKINVDCx5p33_ASAP7_75t_R g1922 ( 
.A(n_1043),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_658),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_304),
.Y(n_1924)
);

INVx1_ASAP7_75t_SL g1925 ( 
.A(n_612),
.Y(n_1925)
);

CKINVDCx5p33_ASAP7_75t_R g1926 ( 
.A(n_1114),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_223),
.Y(n_1927)
);

INVx2_ASAP7_75t_SL g1928 ( 
.A(n_905),
.Y(n_1928)
);

CKINVDCx5p33_ASAP7_75t_R g1929 ( 
.A(n_104),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_187),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_92),
.Y(n_1931)
);

CKINVDCx5p33_ASAP7_75t_R g1932 ( 
.A(n_654),
.Y(n_1932)
);

CKINVDCx16_ASAP7_75t_R g1933 ( 
.A(n_1193),
.Y(n_1933)
);

CKINVDCx16_ASAP7_75t_R g1934 ( 
.A(n_907),
.Y(n_1934)
);

CKINVDCx20_ASAP7_75t_R g1935 ( 
.A(n_1187),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_803),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_358),
.Y(n_1937)
);

CKINVDCx5p33_ASAP7_75t_R g1938 ( 
.A(n_93),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_565),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_82),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1008),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_106),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_228),
.Y(n_1943)
);

CKINVDCx5p33_ASAP7_75t_R g1944 ( 
.A(n_698),
.Y(n_1944)
);

CKINVDCx5p33_ASAP7_75t_R g1945 ( 
.A(n_994),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1107),
.Y(n_1946)
);

CKINVDCx16_ASAP7_75t_R g1947 ( 
.A(n_704),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_1139),
.Y(n_1948)
);

CKINVDCx20_ASAP7_75t_R g1949 ( 
.A(n_1042),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1218),
.Y(n_1950)
);

BUFx6f_ASAP7_75t_L g1951 ( 
.A(n_737),
.Y(n_1951)
);

BUFx10_ASAP7_75t_L g1952 ( 
.A(n_1232),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_936),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1084),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1014),
.Y(n_1955)
);

BUFx10_ASAP7_75t_L g1956 ( 
.A(n_441),
.Y(n_1956)
);

CKINVDCx20_ASAP7_75t_R g1957 ( 
.A(n_1030),
.Y(n_1957)
);

CKINVDCx5p33_ASAP7_75t_R g1958 ( 
.A(n_276),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_701),
.Y(n_1959)
);

BUFx2_ASAP7_75t_SL g1960 ( 
.A(n_762),
.Y(n_1960)
);

INVx2_ASAP7_75t_SL g1961 ( 
.A(n_1103),
.Y(n_1961)
);

CKINVDCx5p33_ASAP7_75t_R g1962 ( 
.A(n_669),
.Y(n_1962)
);

BUFx3_ASAP7_75t_L g1963 ( 
.A(n_995),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_159),
.Y(n_1964)
);

CKINVDCx5p33_ASAP7_75t_R g1965 ( 
.A(n_896),
.Y(n_1965)
);

CKINVDCx5p33_ASAP7_75t_R g1966 ( 
.A(n_187),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_368),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1047),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_813),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_97),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1243),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_332),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1147),
.Y(n_1973)
);

INVx2_ASAP7_75t_SL g1974 ( 
.A(n_399),
.Y(n_1974)
);

CKINVDCx5p33_ASAP7_75t_R g1975 ( 
.A(n_924),
.Y(n_1975)
);

CKINVDCx5p33_ASAP7_75t_R g1976 ( 
.A(n_443),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_203),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_562),
.Y(n_1978)
);

CKINVDCx5p33_ASAP7_75t_R g1979 ( 
.A(n_992),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_720),
.Y(n_1980)
);

CKINVDCx5p33_ASAP7_75t_R g1981 ( 
.A(n_332),
.Y(n_1981)
);

CKINVDCx5p33_ASAP7_75t_R g1982 ( 
.A(n_1154),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_953),
.Y(n_1983)
);

CKINVDCx5p33_ASAP7_75t_R g1984 ( 
.A(n_1070),
.Y(n_1984)
);

CKINVDCx5p33_ASAP7_75t_R g1985 ( 
.A(n_976),
.Y(n_1985)
);

CKINVDCx5p33_ASAP7_75t_R g1986 ( 
.A(n_1077),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1159),
.Y(n_1987)
);

CKINVDCx5p33_ASAP7_75t_R g1988 ( 
.A(n_156),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_900),
.Y(n_1989)
);

CKINVDCx5p33_ASAP7_75t_R g1990 ( 
.A(n_355),
.Y(n_1990)
);

CKINVDCx20_ASAP7_75t_R g1991 ( 
.A(n_1024),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_535),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_974),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_906),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_237),
.Y(n_1995)
);

BUFx6f_ASAP7_75t_L g1996 ( 
.A(n_769),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_392),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_405),
.Y(n_1998)
);

CKINVDCx5p33_ASAP7_75t_R g1999 ( 
.A(n_298),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_547),
.Y(n_2000)
);

CKINVDCx5p33_ASAP7_75t_R g2001 ( 
.A(n_101),
.Y(n_2001)
);

CKINVDCx5p33_ASAP7_75t_R g2002 ( 
.A(n_1066),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_972),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_1013),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_318),
.Y(n_2005)
);

CKINVDCx5p33_ASAP7_75t_R g2006 ( 
.A(n_960),
.Y(n_2006)
);

CKINVDCx20_ASAP7_75t_R g2007 ( 
.A(n_382),
.Y(n_2007)
);

CKINVDCx5p33_ASAP7_75t_R g2008 ( 
.A(n_201),
.Y(n_2008)
);

BUFx3_ASAP7_75t_L g2009 ( 
.A(n_1130),
.Y(n_2009)
);

BUFx6f_ASAP7_75t_L g2010 ( 
.A(n_466),
.Y(n_2010)
);

CKINVDCx5p33_ASAP7_75t_R g2011 ( 
.A(n_858),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_734),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_470),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_182),
.Y(n_2014)
);

CKINVDCx20_ASAP7_75t_R g2015 ( 
.A(n_403),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1082),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_94),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_119),
.Y(n_2018)
);

CKINVDCx20_ASAP7_75t_R g2019 ( 
.A(n_79),
.Y(n_2019)
);

CKINVDCx20_ASAP7_75t_R g2020 ( 
.A(n_952),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_834),
.Y(n_2021)
);

CKINVDCx5p33_ASAP7_75t_R g2022 ( 
.A(n_897),
.Y(n_2022)
);

INVx2_ASAP7_75t_SL g2023 ( 
.A(n_1226),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1017),
.Y(n_2024)
);

CKINVDCx5p33_ASAP7_75t_R g2025 ( 
.A(n_1168),
.Y(n_2025)
);

CKINVDCx16_ASAP7_75t_R g2026 ( 
.A(n_1051),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_1068),
.Y(n_2027)
);

BUFx2_ASAP7_75t_L g2028 ( 
.A(n_596),
.Y(n_2028)
);

CKINVDCx5p33_ASAP7_75t_R g2029 ( 
.A(n_646),
.Y(n_2029)
);

CKINVDCx5p33_ASAP7_75t_R g2030 ( 
.A(n_1144),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_7),
.Y(n_2031)
);

BUFx3_ASAP7_75t_L g2032 ( 
.A(n_307),
.Y(n_2032)
);

CKINVDCx5p33_ASAP7_75t_R g2033 ( 
.A(n_331),
.Y(n_2033)
);

BUFx5_ASAP7_75t_L g2034 ( 
.A(n_520),
.Y(n_2034)
);

CKINVDCx5p33_ASAP7_75t_R g2035 ( 
.A(n_1111),
.Y(n_2035)
);

CKINVDCx5p33_ASAP7_75t_R g2036 ( 
.A(n_285),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_217),
.Y(n_2037)
);

CKINVDCx5p33_ASAP7_75t_R g2038 ( 
.A(n_600),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_889),
.Y(n_2039)
);

CKINVDCx5p33_ASAP7_75t_R g2040 ( 
.A(n_1045),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1151),
.Y(n_2041)
);

CKINVDCx5p33_ASAP7_75t_R g2042 ( 
.A(n_925),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_949),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1190),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_517),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_637),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1058),
.Y(n_2047)
);

CKINVDCx5p33_ASAP7_75t_R g2048 ( 
.A(n_903),
.Y(n_2048)
);

CKINVDCx5p33_ASAP7_75t_R g2049 ( 
.A(n_476),
.Y(n_2049)
);

CKINVDCx20_ASAP7_75t_R g2050 ( 
.A(n_628),
.Y(n_2050)
);

CKINVDCx5p33_ASAP7_75t_R g2051 ( 
.A(n_786),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1011),
.Y(n_2052)
);

CKINVDCx5p33_ASAP7_75t_R g2053 ( 
.A(n_372),
.Y(n_2053)
);

CKINVDCx5p33_ASAP7_75t_R g2054 ( 
.A(n_998),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_298),
.Y(n_2055)
);

CKINVDCx5p33_ASAP7_75t_R g2056 ( 
.A(n_691),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_922),
.Y(n_2057)
);

INVxp67_ASAP7_75t_L g2058 ( 
.A(n_612),
.Y(n_2058)
);

CKINVDCx20_ASAP7_75t_R g2059 ( 
.A(n_306),
.Y(n_2059)
);

CKINVDCx5p33_ASAP7_75t_R g2060 ( 
.A(n_50),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_46),
.Y(n_2061)
);

CKINVDCx5p33_ASAP7_75t_R g2062 ( 
.A(n_887),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_568),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_143),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_902),
.Y(n_2065)
);

CKINVDCx5p33_ASAP7_75t_R g2066 ( 
.A(n_950),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1032),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_664),
.Y(n_2068)
);

CKINVDCx5p33_ASAP7_75t_R g2069 ( 
.A(n_656),
.Y(n_2069)
);

INVx2_ASAP7_75t_SL g2070 ( 
.A(n_1292),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1277),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1277),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1277),
.Y(n_2073)
);

CKINVDCx5p33_ASAP7_75t_R g2074 ( 
.A(n_1366),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1277),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1277),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1417),
.Y(n_2077)
);

CKINVDCx20_ASAP7_75t_R g2078 ( 
.A(n_1284),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1417),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1417),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1417),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1417),
.Y(n_2082)
);

CKINVDCx20_ASAP7_75t_R g2083 ( 
.A(n_1298),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1724),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1724),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1724),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1724),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1724),
.Y(n_2088)
);

CKINVDCx5p33_ASAP7_75t_R g2089 ( 
.A(n_1251),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1806),
.Y(n_2090)
);

CKINVDCx5p33_ASAP7_75t_R g2091 ( 
.A(n_1252),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1806),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1806),
.Y(n_2093)
);

INVxp33_ASAP7_75t_L g2094 ( 
.A(n_1290),
.Y(n_2094)
);

CKINVDCx5p33_ASAP7_75t_R g2095 ( 
.A(n_1253),
.Y(n_2095)
);

INVx1_ASAP7_75t_SL g2096 ( 
.A(n_1353),
.Y(n_2096)
);

INVxp67_ASAP7_75t_L g2097 ( 
.A(n_2028),
.Y(n_2097)
);

BUFx3_ASAP7_75t_L g2098 ( 
.A(n_1590),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1806),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1806),
.Y(n_2100)
);

INVxp33_ASAP7_75t_SL g2101 ( 
.A(n_1487),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2034),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2034),
.Y(n_2103)
);

INVxp67_ASAP7_75t_SL g2104 ( 
.A(n_1504),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2034),
.Y(n_2105)
);

BUFx3_ASAP7_75t_L g2106 ( 
.A(n_1590),
.Y(n_2106)
);

CKINVDCx5p33_ASAP7_75t_R g2107 ( 
.A(n_1255),
.Y(n_2107)
);

CKINVDCx5p33_ASAP7_75t_R g2108 ( 
.A(n_1257),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2034),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2034),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1737),
.Y(n_2111)
);

CKINVDCx16_ASAP7_75t_R g2112 ( 
.A(n_1286),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1737),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1363),
.Y(n_2114)
);

CKINVDCx20_ASAP7_75t_R g2115 ( 
.A(n_1330),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1363),
.Y(n_2116)
);

CKINVDCx14_ASAP7_75t_R g2117 ( 
.A(n_1312),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1363),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1509),
.Y(n_2119)
);

CKINVDCx5p33_ASAP7_75t_R g2120 ( 
.A(n_1272),
.Y(n_2120)
);

INVx1_ASAP7_75t_SL g2121 ( 
.A(n_1434),
.Y(n_2121)
);

CKINVDCx5p33_ASAP7_75t_R g2122 ( 
.A(n_1273),
.Y(n_2122)
);

CKINVDCx5p33_ASAP7_75t_R g2123 ( 
.A(n_1274),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1509),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1509),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1542),
.Y(n_2126)
);

CKINVDCx20_ASAP7_75t_R g2127 ( 
.A(n_1332),
.Y(n_2127)
);

INVx1_ASAP7_75t_SL g2128 ( 
.A(n_1503),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1542),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1542),
.Y(n_2130)
);

INVxp67_ASAP7_75t_SL g2131 ( 
.A(n_1633),
.Y(n_2131)
);

INVxp67_ASAP7_75t_SL g2132 ( 
.A(n_1352),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1553),
.Y(n_2133)
);

INVxp67_ASAP7_75t_L g2134 ( 
.A(n_1652),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1553),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1553),
.Y(n_2136)
);

INVxp67_ASAP7_75t_SL g2137 ( 
.A(n_1735),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1651),
.Y(n_2138)
);

INVxp33_ASAP7_75t_SL g2139 ( 
.A(n_1250),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1651),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1651),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1668),
.Y(n_2142)
);

CKINVDCx5p33_ASAP7_75t_R g2143 ( 
.A(n_1280),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1668),
.Y(n_2144)
);

CKINVDCx5p33_ASAP7_75t_R g2145 ( 
.A(n_1287),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1668),
.Y(n_2146)
);

CKINVDCx16_ASAP7_75t_R g2147 ( 
.A(n_1466),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1673),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1673),
.Y(n_2149)
);

INVxp33_ASAP7_75t_SL g2150 ( 
.A(n_1258),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1673),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1863),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1863),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1863),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1882),
.Y(n_2155)
);

INVxp67_ASAP7_75t_SL g2156 ( 
.A(n_1819),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_1882),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1882),
.Y(n_2158)
);

CKINVDCx14_ASAP7_75t_R g2159 ( 
.A(n_1315),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1951),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_1951),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1951),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1996),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1996),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1996),
.Y(n_2165)
);

CKINVDCx20_ASAP7_75t_R g2166 ( 
.A(n_1423),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2010),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2010),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2010),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_1320),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1313),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1377),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_1320),
.Y(n_2173)
);

CKINVDCx20_ASAP7_75t_R g2174 ( 
.A(n_1440),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1458),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1519),
.Y(n_2176)
);

INVxp33_ASAP7_75t_L g2177 ( 
.A(n_1249),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_1320),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1557),
.Y(n_2179)
);

CKINVDCx5p33_ASAP7_75t_R g2180 ( 
.A(n_1289),
.Y(n_2180)
);

INVxp67_ASAP7_75t_L g2181 ( 
.A(n_1292),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_1320),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1637),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1644),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1686),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1691),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1792),
.Y(n_2187)
);

CKINVDCx5p33_ASAP7_75t_R g2188 ( 
.A(n_1295),
.Y(n_2188)
);

BUFx2_ASAP7_75t_L g2189 ( 
.A(n_1843),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1872),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1921),
.Y(n_2191)
);

INVx1_ASAP7_75t_SL g2192 ( 
.A(n_1505),
.Y(n_2192)
);

HB1xp67_ASAP7_75t_L g2193 ( 
.A(n_1512),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2032),
.Y(n_2194)
);

CKINVDCx14_ASAP7_75t_R g2195 ( 
.A(n_1393),
.Y(n_2195)
);

CKINVDCx5p33_ASAP7_75t_R g2196 ( 
.A(n_1296),
.Y(n_2196)
);

HB1xp67_ASAP7_75t_L g2197 ( 
.A(n_1528),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2063),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2064),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2065),
.Y(n_2200)
);

HB1xp67_ASAP7_75t_L g2201 ( 
.A(n_1582),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_1320),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2068),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1256),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1262),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1263),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2057),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2061),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1265),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1270),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1271),
.Y(n_2211)
);

CKINVDCx5p33_ASAP7_75t_R g2212 ( 
.A(n_1297),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1275),
.Y(n_2213)
);

BUFx10_ASAP7_75t_L g2214 ( 
.A(n_1264),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1278),
.Y(n_2215)
);

INVx1_ASAP7_75t_SL g2216 ( 
.A(n_1780),
.Y(n_2216)
);

BUFx3_ASAP7_75t_L g2217 ( 
.A(n_1658),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1283),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1293),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1307),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1311),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1314),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1317),
.Y(n_2223)
);

BUFx3_ASAP7_75t_L g2224 ( 
.A(n_1658),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1326),
.Y(n_2225)
);

INVxp67_ASAP7_75t_SL g2226 ( 
.A(n_1878),
.Y(n_2226)
);

BUFx3_ASAP7_75t_L g2227 ( 
.A(n_1702),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1335),
.Y(n_2228)
);

INVxp33_ASAP7_75t_SL g2229 ( 
.A(n_1267),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1337),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1341),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1343),
.Y(n_2232)
);

OR2x2_ASAP7_75t_L g2233 ( 
.A(n_1254),
.B(n_0),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1362),
.Y(n_2234)
);

NOR2xp33_ASAP7_75t_L g2235 ( 
.A(n_1570),
.B(n_1583),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1365),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1373),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1380),
.Y(n_2238)
);

INVxp33_ASAP7_75t_L g2239 ( 
.A(n_1385),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1386),
.Y(n_2240)
);

BUFx6f_ASAP7_75t_L g2241 ( 
.A(n_2133),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_2142),
.Y(n_2242)
);

BUFx6f_ASAP7_75t_L g2243 ( 
.A(n_2157),
.Y(n_2243)
);

AND2x6_ASAP7_75t_L g2244 ( 
.A(n_2098),
.B(n_1260),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2161),
.Y(n_2245)
);

BUFx12f_ASAP7_75t_L g2246 ( 
.A(n_2074),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2089),
.B(n_1323),
.Y(n_2247)
);

AOI22xp5_ASAP7_75t_L g2248 ( 
.A1(n_2101),
.A2(n_1862),
.B1(n_1933),
.B2(n_1351),
.Y(n_2248)
);

BUFx2_ASAP7_75t_L g2249 ( 
.A(n_2117),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2114),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2116),
.Y(n_2251)
);

CKINVDCx5p33_ASAP7_75t_R g2252 ( 
.A(n_2091),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2118),
.Y(n_2253)
);

CKINVDCx5p33_ASAP7_75t_R g2254 ( 
.A(n_2095),
.Y(n_2254)
);

INVx3_ASAP7_75t_L g2255 ( 
.A(n_2119),
.Y(n_2255)
);

OA21x2_ASAP7_75t_L g2256 ( 
.A1(n_2071),
.A2(n_1918),
.B(n_1876),
.Y(n_2256)
);

NOR2x1_ASAP7_75t_L g2257 ( 
.A(n_2106),
.B(n_1891),
.Y(n_2257)
);

BUFx6f_ASAP7_75t_L g2258 ( 
.A(n_2124),
.Y(n_2258)
);

BUFx6f_ASAP7_75t_L g2259 ( 
.A(n_2125),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2107),
.B(n_1547),
.Y(n_2260)
);

BUFx6f_ASAP7_75t_L g2261 ( 
.A(n_2126),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_2129),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_2130),
.Y(n_2263)
);

INVx3_ASAP7_75t_L g2264 ( 
.A(n_2135),
.Y(n_2264)
);

AND2x4_ASAP7_75t_L g2265 ( 
.A(n_2217),
.B(n_1963),
.Y(n_2265)
);

AND2x4_ASAP7_75t_L g2266 ( 
.A(n_2224),
.B(n_2009),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2136),
.Y(n_2267)
);

NOR2x1_ASAP7_75t_L g2268 ( 
.A(n_2227),
.B(n_1259),
.Y(n_2268)
);

BUFx6f_ASAP7_75t_L g2269 ( 
.A(n_2138),
.Y(n_2269)
);

INVx2_ASAP7_75t_SL g2270 ( 
.A(n_2214),
.Y(n_2270)
);

BUFx2_ASAP7_75t_L g2271 ( 
.A(n_2159),
.Y(n_2271)
);

INVx3_ASAP7_75t_L g2272 ( 
.A(n_2140),
.Y(n_2272)
);

AND2x4_ASAP7_75t_L g2273 ( 
.A(n_2132),
.B(n_1437),
.Y(n_2273)
);

CKINVDCx6p67_ASAP7_75t_R g2274 ( 
.A(n_2112),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_2141),
.Y(n_2275)
);

AND2x2_ASAP7_75t_L g2276 ( 
.A(n_2195),
.B(n_1618),
.Y(n_2276)
);

BUFx6f_ASAP7_75t_L g2277 ( 
.A(n_2144),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2108),
.B(n_1961),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2146),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_2148),
.Y(n_2280)
);

BUFx2_ASAP7_75t_L g2281 ( 
.A(n_2193),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_2137),
.B(n_1818),
.Y(n_2282)
);

INVx5_ASAP7_75t_L g2283 ( 
.A(n_2214),
.Y(n_2283)
);

INVx5_ASAP7_75t_L g2284 ( 
.A(n_2070),
.Y(n_2284)
);

BUFx12f_ASAP7_75t_L g2285 ( 
.A(n_2120),
.Y(n_2285)
);

BUFx12f_ASAP7_75t_L g2286 ( 
.A(n_2122),
.Y(n_2286)
);

BUFx3_ASAP7_75t_L g2287 ( 
.A(n_2189),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_2149),
.Y(n_2288)
);

BUFx6f_ASAP7_75t_L g2289 ( 
.A(n_2151),
.Y(n_2289)
);

HB1xp67_ASAP7_75t_L g2290 ( 
.A(n_2197),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2152),
.Y(n_2291)
);

BUFx2_ASAP7_75t_L g2292 ( 
.A(n_2201),
.Y(n_2292)
);

HB1xp67_ASAP7_75t_L g2293 ( 
.A(n_2147),
.Y(n_2293)
);

INVx3_ASAP7_75t_L g2294 ( 
.A(n_2153),
.Y(n_2294)
);

BUFx2_ASAP7_75t_L g2295 ( 
.A(n_2123),
.Y(n_2295)
);

OA21x2_ASAP7_75t_L g2296 ( 
.A1(n_2072),
.A2(n_2076),
.B(n_2073),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2154),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_2155),
.Y(n_2298)
);

BUFx12f_ASAP7_75t_L g2299 ( 
.A(n_2143),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2158),
.Y(n_2300)
);

OA21x2_ASAP7_75t_L g2301 ( 
.A1(n_2077),
.A2(n_2080),
.B(n_2079),
.Y(n_2301)
);

AND2x4_ASAP7_75t_L g2302 ( 
.A(n_2156),
.B(n_2226),
.Y(n_2302)
);

BUFx12f_ASAP7_75t_L g2303 ( 
.A(n_2145),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_2160),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2162),
.Y(n_2305)
);

HB1xp67_ASAP7_75t_L g2306 ( 
.A(n_2121),
.Y(n_2306)
);

CKINVDCx5p33_ASAP7_75t_R g2307 ( 
.A(n_2180),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2163),
.Y(n_2308)
);

OA21x2_ASAP7_75t_L g2309 ( 
.A1(n_2081),
.A2(n_1291),
.B(n_1285),
.Y(n_2309)
);

INVx4_ASAP7_75t_L g2310 ( 
.A(n_2188),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2196),
.B(n_2023),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2164),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2165),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2167),
.Y(n_2314)
);

OAI21x1_ASAP7_75t_L g2315 ( 
.A1(n_2075),
.A2(n_1322),
.B(n_1299),
.Y(n_2315)
);

BUFx12f_ASAP7_75t_L g2316 ( 
.A(n_2212),
.Y(n_2316)
);

INVx5_ASAP7_75t_L g2317 ( 
.A(n_2170),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2168),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2235),
.B(n_1388),
.Y(n_2319)
);

INVx5_ASAP7_75t_L g2320 ( 
.A(n_2173),
.Y(n_2320)
);

AND2x4_ASAP7_75t_L g2321 ( 
.A(n_2104),
.B(n_1736),
.Y(n_2321)
);

INVxp33_ASAP7_75t_SL g2322 ( 
.A(n_2128),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2169),
.Y(n_2323)
);

BUFx12f_ASAP7_75t_L g2324 ( 
.A(n_2233),
.Y(n_2324)
);

INVx5_ASAP7_75t_L g2325 ( 
.A(n_2178),
.Y(n_2325)
);

BUFx6f_ASAP7_75t_L g2326 ( 
.A(n_2198),
.Y(n_2326)
);

INVx3_ASAP7_75t_L g2327 ( 
.A(n_2171),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2082),
.Y(n_2328)
);

OAI22xp5_ASAP7_75t_L g2329 ( 
.A1(n_2096),
.A2(n_2097),
.B1(n_2131),
.B2(n_2094),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2084),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2085),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_2086),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2087),
.Y(n_2333)
);

HB1xp67_ASAP7_75t_L g2334 ( 
.A(n_2192),
.Y(n_2334)
);

BUFx12f_ASAP7_75t_L g2335 ( 
.A(n_2139),
.Y(n_2335)
);

INVx4_ASAP7_75t_L g2336 ( 
.A(n_2182),
.Y(n_2336)
);

BUFx6f_ASAP7_75t_L g2337 ( 
.A(n_2199),
.Y(n_2337)
);

BUFx2_ASAP7_75t_L g2338 ( 
.A(n_2181),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2088),
.Y(n_2339)
);

INVx5_ASAP7_75t_L g2340 ( 
.A(n_2202),
.Y(n_2340)
);

BUFx12f_ASAP7_75t_L g2341 ( 
.A(n_2150),
.Y(n_2341)
);

NOR2x1_ASAP7_75t_L g2342 ( 
.A(n_2090),
.B(n_1302),
.Y(n_2342)
);

AND2x4_ASAP7_75t_L g2343 ( 
.A(n_2134),
.B(n_1303),
.Y(n_2343)
);

NOR2xp33_ASAP7_75t_L g2344 ( 
.A(n_2229),
.B(n_2026),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2092),
.Y(n_2345)
);

BUFx6f_ASAP7_75t_L g2346 ( 
.A(n_2200),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_2093),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2177),
.B(n_1879),
.Y(n_2348)
);

BUFx6f_ASAP7_75t_L g2349 ( 
.A(n_2203),
.Y(n_2349)
);

INVx6_ASAP7_75t_L g2350 ( 
.A(n_2239),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2099),
.Y(n_2351)
);

OAI22xp5_ASAP7_75t_L g2352 ( 
.A1(n_2216),
.A2(n_1934),
.B1(n_1947),
.B2(n_1919),
.Y(n_2352)
);

AND2x4_ASAP7_75t_L g2353 ( 
.A(n_2172),
.B(n_1308),
.Y(n_2353)
);

AOI22x1_ASAP7_75t_SL g2354 ( 
.A1(n_2078),
.A2(n_1269),
.B1(n_1360),
.B2(n_1261),
.Y(n_2354)
);

BUFx6f_ASAP7_75t_L g2355 ( 
.A(n_2204),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2100),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2102),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2103),
.Y(n_2358)
);

AND2x4_ASAP7_75t_L g2359 ( 
.A(n_2175),
.B(n_1325),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2176),
.B(n_1430),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2105),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2109),
.Y(n_2362)
);

INVx2_ASAP7_75t_SL g2363 ( 
.A(n_2179),
.Y(n_2363)
);

BUFx3_ASAP7_75t_L g2364 ( 
.A(n_2183),
.Y(n_2364)
);

AND2x4_ASAP7_75t_L g2365 ( 
.A(n_2184),
.B(n_1327),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2110),
.Y(n_2366)
);

BUFx12f_ASAP7_75t_L g2367 ( 
.A(n_2083),
.Y(n_2367)
);

BUFx6f_ASAP7_75t_L g2368 ( 
.A(n_2205),
.Y(n_2368)
);

CKINVDCx6p67_ASAP7_75t_R g2369 ( 
.A(n_2115),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2185),
.B(n_1608),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_2186),
.B(n_1702),
.Y(n_2371)
);

BUFx6f_ASAP7_75t_L g2372 ( 
.A(n_2206),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2111),
.Y(n_2373)
);

BUFx8_ASAP7_75t_L g2374 ( 
.A(n_2187),
.Y(n_2374)
);

INVx4_ASAP7_75t_L g2375 ( 
.A(n_2190),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2113),
.Y(n_2376)
);

HB1xp67_ASAP7_75t_L g2377 ( 
.A(n_2191),
.Y(n_2377)
);

BUFx2_ASAP7_75t_L g2378 ( 
.A(n_2194),
.Y(n_2378)
);

BUFx12f_ASAP7_75t_L g2379 ( 
.A(n_2127),
.Y(n_2379)
);

BUFx6f_ASAP7_75t_L g2380 ( 
.A(n_2207),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2208),
.Y(n_2381)
);

INVx5_ASAP7_75t_L g2382 ( 
.A(n_2209),
.Y(n_2382)
);

NAND2x1p5_ASAP7_75t_L g2383 ( 
.A(n_2210),
.B(n_1387),
.Y(n_2383)
);

BUFx6f_ASAP7_75t_L g2384 ( 
.A(n_2211),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_2213),
.Y(n_2385)
);

AND2x2_ASAP7_75t_L g2386 ( 
.A(n_2215),
.B(n_1952),
.Y(n_2386)
);

CKINVDCx5p33_ASAP7_75t_R g2387 ( 
.A(n_2166),
.Y(n_2387)
);

INVx3_ASAP7_75t_L g2388 ( 
.A(n_2218),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_2219),
.B(n_1952),
.Y(n_2389)
);

AND2x6_ASAP7_75t_L g2390 ( 
.A(n_2220),
.B(n_1340),
.Y(n_2390)
);

BUFx8_ASAP7_75t_L g2391 ( 
.A(n_2221),
.Y(n_2391)
);

BUFx6f_ASAP7_75t_L g2392 ( 
.A(n_2222),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2223),
.Y(n_2393)
);

AND2x2_ASAP7_75t_L g2394 ( 
.A(n_2225),
.B(n_1685),
.Y(n_2394)
);

CKINVDCx11_ASAP7_75t_R g2395 ( 
.A(n_2174),
.Y(n_2395)
);

BUFx2_ASAP7_75t_L g2396 ( 
.A(n_2228),
.Y(n_2396)
);

BUFx6f_ASAP7_75t_L g2397 ( 
.A(n_2230),
.Y(n_2397)
);

AND2x4_ASAP7_75t_L g2398 ( 
.A(n_2231),
.B(n_1328),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2232),
.Y(n_2399)
);

INVx4_ASAP7_75t_L g2400 ( 
.A(n_2234),
.Y(n_2400)
);

OA21x2_ASAP7_75t_L g2401 ( 
.A1(n_2236),
.A2(n_1359),
.B(n_1349),
.Y(n_2401)
);

INVxp33_ASAP7_75t_SL g2402 ( 
.A(n_2237),
.Y(n_2402)
);

AND2x2_ASAP7_75t_L g2403 ( 
.A(n_2238),
.B(n_1279),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2240),
.B(n_1664),
.Y(n_2404)
);

BUFx12f_ASAP7_75t_L g2405 ( 
.A(n_2074),
.Y(n_2405)
);

BUFx3_ASAP7_75t_L g2406 ( 
.A(n_2189),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2133),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_2133),
.Y(n_2408)
);

AOI22xp5_ASAP7_75t_L g2409 ( 
.A1(n_2101),
.A2(n_1523),
.B1(n_1580),
.B2(n_1508),
.Y(n_2409)
);

INVx3_ASAP7_75t_L g2410 ( 
.A(n_2133),
.Y(n_2410)
);

AND2x4_ASAP7_75t_L g2411 ( 
.A(n_2098),
.B(n_1367),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2133),
.Y(n_2412)
);

AOI22xp5_ASAP7_75t_L g2413 ( 
.A1(n_2101),
.A2(n_1603),
.B1(n_1612),
.B2(n_1594),
.Y(n_2413)
);

BUFx8_ASAP7_75t_SL g2414 ( 
.A(n_2074),
.Y(n_2414)
);

OAI21x1_ASAP7_75t_L g2415 ( 
.A1(n_2075),
.A2(n_1703),
.B(n_1679),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_2133),
.Y(n_2416)
);

INVx2_ASAP7_75t_SL g2417 ( 
.A(n_2214),
.Y(n_2417)
);

HB1xp67_ASAP7_75t_L g2418 ( 
.A(n_2193),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2133),
.Y(n_2419)
);

BUFx8_ASAP7_75t_SL g2420 ( 
.A(n_2074),
.Y(n_2420)
);

INVx5_ASAP7_75t_L g2421 ( 
.A(n_2214),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2117),
.B(n_1465),
.Y(n_2422)
);

INVx3_ASAP7_75t_L g2423 ( 
.A(n_2133),
.Y(n_2423)
);

INVx4_ASAP7_75t_L g2424 ( 
.A(n_2089),
.Y(n_2424)
);

BUFx3_ASAP7_75t_L g2425 ( 
.A(n_2189),
.Y(n_2425)
);

HB1xp67_ASAP7_75t_L g2426 ( 
.A(n_2193),
.Y(n_2426)
);

INVxp67_ASAP7_75t_L g2427 ( 
.A(n_2193),
.Y(n_2427)
);

AOI22xp5_ASAP7_75t_L g2428 ( 
.A1(n_2101),
.A2(n_1844),
.B1(n_1935),
.B2(n_1798),
.Y(n_2428)
);

BUFx12f_ASAP7_75t_L g2429 ( 
.A(n_2074),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2133),
.Y(n_2430)
);

OA21x2_ASAP7_75t_L g2431 ( 
.A1(n_2071),
.A2(n_1371),
.B(n_1368),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2133),
.Y(n_2432)
);

INVx4_ASAP7_75t_L g2433 ( 
.A(n_2089),
.Y(n_2433)
);

BUFx6f_ASAP7_75t_L g2434 ( 
.A(n_2133),
.Y(n_2434)
);

INVx3_ASAP7_75t_L g2435 ( 
.A(n_2133),
.Y(n_2435)
);

BUFx12f_ASAP7_75t_L g2436 ( 
.A(n_2074),
.Y(n_2436)
);

OAI21x1_ASAP7_75t_L g2437 ( 
.A1(n_2075),
.A2(n_1824),
.B(n_1719),
.Y(n_2437)
);

BUFx3_ASAP7_75t_L g2438 ( 
.A(n_2189),
.Y(n_2438)
);

BUFx2_ASAP7_75t_L g2439 ( 
.A(n_2117),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2133),
.Y(n_2440)
);

INVx3_ASAP7_75t_L g2441 ( 
.A(n_2133),
.Y(n_2441)
);

BUFx12f_ASAP7_75t_L g2442 ( 
.A(n_2074),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2133),
.Y(n_2443)
);

BUFx12f_ASAP7_75t_L g2444 ( 
.A(n_2074),
.Y(n_2444)
);

AOI22x1_ASAP7_75t_SL g2445 ( 
.A1(n_2078),
.A2(n_1460),
.B1(n_1506),
.B2(n_1391),
.Y(n_2445)
);

HB1xp67_ASAP7_75t_L g2446 ( 
.A(n_2193),
.Y(n_2446)
);

INVx5_ASAP7_75t_L g2447 ( 
.A(n_2214),
.Y(n_2447)
);

INVx4_ASAP7_75t_L g2448 ( 
.A(n_2089),
.Y(n_2448)
);

BUFx12f_ASAP7_75t_L g2449 ( 
.A(n_2074),
.Y(n_2449)
);

AND2x6_ASAP7_75t_L g2450 ( 
.A(n_2098),
.B(n_1511),
.Y(n_2450)
);

CKINVDCx5p33_ASAP7_75t_R g2451 ( 
.A(n_2089),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2133),
.Y(n_2452)
);

BUFx8_ASAP7_75t_SL g2453 ( 
.A(n_2074),
.Y(n_2453)
);

BUFx6f_ASAP7_75t_L g2454 ( 
.A(n_2133),
.Y(n_2454)
);

OAI21x1_ASAP7_75t_L g2455 ( 
.A1(n_2075),
.A2(n_1955),
.B(n_1946),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2133),
.Y(n_2456)
);

INVx3_ASAP7_75t_L g2457 ( 
.A(n_2133),
.Y(n_2457)
);

BUFx8_ASAP7_75t_SL g2458 ( 
.A(n_2074),
.Y(n_2458)
);

BUFx3_ASAP7_75t_L g2459 ( 
.A(n_2189),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2133),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2133),
.Y(n_2461)
);

BUFx6f_ASAP7_75t_L g2462 ( 
.A(n_2133),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2133),
.Y(n_2463)
);

BUFx6f_ASAP7_75t_L g2464 ( 
.A(n_2133),
.Y(n_2464)
);

NOR2xp33_ASAP7_75t_L g2465 ( 
.A(n_2235),
.B(n_1390),
.Y(n_2465)
);

BUFx3_ASAP7_75t_L g2466 ( 
.A(n_2189),
.Y(n_2466)
);

AOI22xp5_ASAP7_75t_L g2467 ( 
.A1(n_2101),
.A2(n_1957),
.B1(n_1991),
.B2(n_1949),
.Y(n_2467)
);

INVx2_ASAP7_75t_SL g2468 ( 
.A(n_2214),
.Y(n_2468)
);

INVx5_ASAP7_75t_L g2469 ( 
.A(n_2214),
.Y(n_2469)
);

INVx6_ASAP7_75t_L g2470 ( 
.A(n_2214),
.Y(n_2470)
);

AND2x2_ASAP7_75t_L g2471 ( 
.A(n_2117),
.B(n_1480),
.Y(n_2471)
);

BUFx6f_ASAP7_75t_L g2472 ( 
.A(n_2133),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2133),
.Y(n_2473)
);

HB1xp67_ASAP7_75t_L g2474 ( 
.A(n_2193),
.Y(n_2474)
);

INVx3_ASAP7_75t_L g2475 ( 
.A(n_2133),
.Y(n_2475)
);

INVx5_ASAP7_75t_L g2476 ( 
.A(n_2214),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2133),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2133),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2133),
.Y(n_2479)
);

CKINVDCx5p33_ASAP7_75t_R g2480 ( 
.A(n_2089),
.Y(n_2480)
);

AND2x4_ASAP7_75t_L g2481 ( 
.A(n_2098),
.B(n_1408),
.Y(n_2481)
);

BUFx6f_ASAP7_75t_L g2482 ( 
.A(n_2133),
.Y(n_2482)
);

BUFx6f_ASAP7_75t_L g2483 ( 
.A(n_2133),
.Y(n_2483)
);

BUFx12f_ASAP7_75t_L g2484 ( 
.A(n_2074),
.Y(n_2484)
);

BUFx6f_ASAP7_75t_L g2485 ( 
.A(n_2133),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_2133),
.Y(n_2486)
);

INVx5_ASAP7_75t_L g2487 ( 
.A(n_2214),
.Y(n_2487)
);

BUFx3_ASAP7_75t_L g2488 ( 
.A(n_2189),
.Y(n_2488)
);

BUFx6f_ASAP7_75t_L g2489 ( 
.A(n_2133),
.Y(n_2489)
);

BUFx6f_ASAP7_75t_L g2490 ( 
.A(n_2133),
.Y(n_2490)
);

OAI21x1_ASAP7_75t_L g2491 ( 
.A1(n_2075),
.A2(n_2041),
.B(n_2016),
.Y(n_2491)
);

AND2x2_ASAP7_75t_L g2492 ( 
.A(n_2117),
.B(n_1484),
.Y(n_2492)
);

AND2x4_ASAP7_75t_L g2493 ( 
.A(n_2098),
.B(n_1413),
.Y(n_2493)
);

HB1xp67_ASAP7_75t_L g2494 ( 
.A(n_2193),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2133),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2133),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2133),
.Y(n_2497)
);

BUFx6f_ASAP7_75t_L g2498 ( 
.A(n_2133),
.Y(n_2498)
);

BUFx12f_ASAP7_75t_L g2499 ( 
.A(n_2074),
.Y(n_2499)
);

INVx2_ASAP7_75t_L g2500 ( 
.A(n_2133),
.Y(n_2500)
);

INVx3_ASAP7_75t_L g2501 ( 
.A(n_2133),
.Y(n_2501)
);

BUFx6f_ASAP7_75t_L g2502 ( 
.A(n_2133),
.Y(n_2502)
);

BUFx12f_ASAP7_75t_L g2503 ( 
.A(n_2074),
.Y(n_2503)
);

BUFx2_ASAP7_75t_L g2504 ( 
.A(n_2117),
.Y(n_2504)
);

AND2x4_ASAP7_75t_L g2505 ( 
.A(n_2098),
.B(n_1418),
.Y(n_2505)
);

BUFx6f_ASAP7_75t_L g2506 ( 
.A(n_2133),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2133),
.Y(n_2507)
);

NOR2xp33_ASAP7_75t_L g2508 ( 
.A(n_2235),
.B(n_1425),
.Y(n_2508)
);

AND2x2_ASAP7_75t_L g2509 ( 
.A(n_2117),
.B(n_1753),
.Y(n_2509)
);

BUFx3_ASAP7_75t_L g2510 ( 
.A(n_2189),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2133),
.Y(n_2511)
);

AND2x4_ASAP7_75t_L g2512 ( 
.A(n_2098),
.B(n_1444),
.Y(n_2512)
);

OAI22x1_ASAP7_75t_SL g2513 ( 
.A1(n_2101),
.A2(n_1564),
.B1(n_1581),
.B2(n_1543),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2133),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_2089),
.B(n_2052),
.Y(n_2515)
);

CKINVDCx5p33_ASAP7_75t_R g2516 ( 
.A(n_2089),
.Y(n_2516)
);

NOR2x1_ASAP7_75t_L g2517 ( 
.A(n_2098),
.B(n_1450),
.Y(n_2517)
);

BUFx8_ASAP7_75t_L g2518 ( 
.A(n_2070),
.Y(n_2518)
);

INVx2_ASAP7_75t_L g2519 ( 
.A(n_2133),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2133),
.Y(n_2520)
);

BUFx12f_ASAP7_75t_L g2521 ( 
.A(n_2074),
.Y(n_2521)
);

BUFx6f_ASAP7_75t_L g2522 ( 
.A(n_2133),
.Y(n_2522)
);

AND2x6_ASAP7_75t_L g2523 ( 
.A(n_2098),
.B(n_1530),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2089),
.B(n_1453),
.Y(n_2524)
);

BUFx3_ASAP7_75t_L g2525 ( 
.A(n_2189),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2089),
.B(n_1467),
.Y(n_2526)
);

BUFx6f_ASAP7_75t_L g2527 ( 
.A(n_2133),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2133),
.Y(n_2528)
);

BUFx12f_ASAP7_75t_L g2529 ( 
.A(n_2074),
.Y(n_2529)
);

AND2x2_ASAP7_75t_L g2530 ( 
.A(n_2117),
.B(n_1832),
.Y(n_2530)
);

BUFx6f_ASAP7_75t_L g2531 ( 
.A(n_2133),
.Y(n_2531)
);

BUFx6f_ASAP7_75t_L g2532 ( 
.A(n_2133),
.Y(n_2532)
);

CKINVDCx5p33_ASAP7_75t_R g2533 ( 
.A(n_2089),
.Y(n_2533)
);

BUFx6f_ASAP7_75t_L g2534 ( 
.A(n_2133),
.Y(n_2534)
);

AND2x4_ASAP7_75t_L g2535 ( 
.A(n_2098),
.B(n_1469),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_2133),
.Y(n_2536)
);

BUFx12f_ASAP7_75t_L g2537 ( 
.A(n_2074),
.Y(n_2537)
);

INVx5_ASAP7_75t_L g2538 ( 
.A(n_2214),
.Y(n_2538)
);

OAI22xp33_ASAP7_75t_R g2539 ( 
.A1(n_2121),
.A2(n_1555),
.B1(n_1693),
.B2(n_1533),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2089),
.B(n_1470),
.Y(n_2540)
);

BUFx2_ASAP7_75t_L g2541 ( 
.A(n_2117),
.Y(n_2541)
);

AND2x4_ASAP7_75t_L g2542 ( 
.A(n_2098),
.B(n_1485),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2133),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2133),
.Y(n_2544)
);

BUFx6f_ASAP7_75t_L g2545 ( 
.A(n_2133),
.Y(n_2545)
);

BUFx6f_ASAP7_75t_L g2546 ( 
.A(n_2133),
.Y(n_2546)
);

INVx3_ASAP7_75t_L g2547 ( 
.A(n_2133),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2133),
.Y(n_2548)
);

INVx3_ASAP7_75t_L g2549 ( 
.A(n_2133),
.Y(n_2549)
);

BUFx6f_ASAP7_75t_L g2550 ( 
.A(n_2133),
.Y(n_2550)
);

HB1xp67_ASAP7_75t_L g2551 ( 
.A(n_2193),
.Y(n_2551)
);

CKINVDCx5p33_ASAP7_75t_R g2552 ( 
.A(n_2089),
.Y(n_2552)
);

OA21x2_ASAP7_75t_L g2553 ( 
.A1(n_2071),
.A2(n_1552),
.B(n_1544),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2133),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2117),
.B(n_1907),
.Y(n_2555)
);

INVx5_ASAP7_75t_L g2556 ( 
.A(n_2214),
.Y(n_2556)
);

AND2x2_ASAP7_75t_L g2557 ( 
.A(n_2117),
.B(n_1928),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2133),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2133),
.Y(n_2559)
);

BUFx3_ASAP7_75t_L g2560 ( 
.A(n_2189),
.Y(n_2560)
);

INVx2_ASAP7_75t_L g2561 ( 
.A(n_2133),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2133),
.Y(n_2562)
);

AND2x2_ASAP7_75t_L g2563 ( 
.A(n_2117),
.B(n_1974),
.Y(n_2563)
);

BUFx6f_ASAP7_75t_L g2564 ( 
.A(n_2133),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_SL g2565 ( 
.A(n_2112),
.B(n_1561),
.Y(n_2565)
);

AND2x4_ASAP7_75t_L g2566 ( 
.A(n_2098),
.B(n_1593),
.Y(n_2566)
);

AND2x4_ASAP7_75t_L g2567 ( 
.A(n_2098),
.B(n_1609),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2133),
.Y(n_2568)
);

AOI22x1_ASAP7_75t_SL g2569 ( 
.A1(n_2078),
.A2(n_1620),
.B1(n_1629),
.B2(n_1615),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2133),
.Y(n_2570)
);

BUFx6f_ASAP7_75t_L g2571 ( 
.A(n_2133),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2381),
.Y(n_2572)
);

BUFx6f_ASAP7_75t_L g2573 ( 
.A(n_2241),
.Y(n_2573)
);

BUFx6f_ASAP7_75t_L g2574 ( 
.A(n_2243),
.Y(n_2574)
);

HB1xp67_ASAP7_75t_L g2575 ( 
.A(n_2350),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2393),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2399),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2326),
.Y(n_2578)
);

INVx3_ASAP7_75t_L g2579 ( 
.A(n_2434),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2454),
.Y(n_2580)
);

AND2x4_ASAP7_75t_L g2581 ( 
.A(n_2287),
.B(n_2058),
.Y(n_2581)
);

BUFx6f_ASAP7_75t_L g2582 ( 
.A(n_2462),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2464),
.Y(n_2583)
);

INVx2_ASAP7_75t_L g2584 ( 
.A(n_2472),
.Y(n_2584)
);

NOR2xp33_ASAP7_75t_L g2585 ( 
.A(n_2515),
.B(n_1268),
.Y(n_2585)
);

AND2x6_ASAP7_75t_L g2586 ( 
.A(n_2276),
.B(n_1764),
.Y(n_2586)
);

BUFx6f_ASAP7_75t_L g2587 ( 
.A(n_2482),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2483),
.Y(n_2588)
);

BUFx6f_ASAP7_75t_L g2589 ( 
.A(n_2485),
.Y(n_2589)
);

NOR2xp33_ASAP7_75t_L g2590 ( 
.A(n_2524),
.B(n_1276),
.Y(n_2590)
);

AND2x2_ASAP7_75t_L g2591 ( 
.A(n_2348),
.B(n_1561),
.Y(n_2591)
);

NOR2xp33_ASAP7_75t_L g2592 ( 
.A(n_2526),
.B(n_1281),
.Y(n_2592)
);

CKINVDCx16_ASAP7_75t_R g2593 ( 
.A(n_2306),
.Y(n_2593)
);

AND2x2_ASAP7_75t_L g2594 ( 
.A(n_2282),
.B(n_1625),
.Y(n_2594)
);

AND2x4_ASAP7_75t_L g2595 ( 
.A(n_2406),
.B(n_1394),
.Y(n_2595)
);

INVx2_ASAP7_75t_L g2596 ( 
.A(n_2489),
.Y(n_2596)
);

NOR2x1_ASAP7_75t_L g2597 ( 
.A(n_2344),
.B(n_1631),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_SL g2598 ( 
.A(n_2556),
.B(n_1304),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2337),
.Y(n_2599)
);

BUFx6f_ASAP7_75t_L g2600 ( 
.A(n_2490),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2346),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2498),
.Y(n_2602)
);

HB1xp67_ASAP7_75t_L g2603 ( 
.A(n_2334),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_L g2604 ( 
.A(n_2302),
.B(n_1309),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_2540),
.B(n_1321),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2502),
.Y(n_2606)
);

AND2x4_ASAP7_75t_L g2607 ( 
.A(n_2425),
.B(n_1398),
.Y(n_2607)
);

CKINVDCx16_ASAP7_75t_R g2608 ( 
.A(n_2293),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2349),
.Y(n_2609)
);

INVxp67_ASAP7_75t_L g2610 ( 
.A(n_2338),
.Y(n_2610)
);

HB1xp67_ASAP7_75t_L g2611 ( 
.A(n_2438),
.Y(n_2611)
);

INVx4_ASAP7_75t_L g2612 ( 
.A(n_2285),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2355),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2368),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2336),
.B(n_1324),
.Y(n_2615)
);

HB1xp67_ASAP7_75t_L g2616 ( 
.A(n_2459),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2506),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2372),
.Y(n_2618)
);

INVx3_ASAP7_75t_L g2619 ( 
.A(n_2522),
.Y(n_2619)
);

NOR2xp33_ASAP7_75t_L g2620 ( 
.A(n_2247),
.B(n_1282),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_2527),
.Y(n_2621)
);

NOR2xp33_ASAP7_75t_L g2622 ( 
.A(n_2260),
.B(n_1288),
.Y(n_2622)
);

OR2x2_ASAP7_75t_L g2623 ( 
.A(n_2281),
.B(n_1853),
.Y(n_2623)
);

AND2x4_ASAP7_75t_L g2624 ( 
.A(n_2466),
.B(n_1399),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2380),
.Y(n_2625)
);

BUFx6f_ASAP7_75t_L g2626 ( 
.A(n_2531),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2384),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2392),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2397),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_SL g2630 ( 
.A(n_2556),
.B(n_1331),
.Y(n_2630)
);

INVx3_ASAP7_75t_L g2631 ( 
.A(n_2532),
.Y(n_2631)
);

OA21x2_ASAP7_75t_L g2632 ( 
.A1(n_2315),
.A2(n_1635),
.B(n_1632),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_2465),
.B(n_1334),
.Y(n_2633)
);

AND2x2_ASAP7_75t_L g2634 ( 
.A(n_2321),
.B(n_2273),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2534),
.Y(n_2635)
);

BUFx6f_ASAP7_75t_L g2636 ( 
.A(n_2545),
.Y(n_2636)
);

BUFx6f_ASAP7_75t_L g2637 ( 
.A(n_2546),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2328),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2331),
.Y(n_2639)
);

INVx3_ASAP7_75t_L g2640 ( 
.A(n_2550),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2564),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_L g2642 ( 
.A(n_2508),
.B(n_1338),
.Y(n_2642)
);

OAI22xp5_ASAP7_75t_L g2643 ( 
.A1(n_2248),
.A2(n_2319),
.B1(n_2311),
.B2(n_2278),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2333),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2345),
.Y(n_2645)
);

INVx3_ASAP7_75t_L g2646 ( 
.A(n_2571),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2256),
.B(n_2351),
.Y(n_2647)
);

CKINVDCx20_ASAP7_75t_R g2648 ( 
.A(n_2395),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2357),
.B(n_1342),
.Y(n_2649)
);

HB1xp67_ASAP7_75t_L g2650 ( 
.A(n_2488),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_2358),
.B(n_1345),
.Y(n_2651)
);

AND2x2_ASAP7_75t_L g2652 ( 
.A(n_2386),
.B(n_1625),
.Y(n_2652)
);

INVxp67_ASAP7_75t_L g2653 ( 
.A(n_2292),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2361),
.B(n_1346),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2362),
.Y(n_2655)
);

AOI22xp5_ASAP7_75t_L g2656 ( 
.A1(n_2427),
.A2(n_1412),
.B1(n_1925),
.B2(n_1899),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_SL g2657 ( 
.A(n_2283),
.B(n_2421),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2366),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2242),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2330),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2408),
.Y(n_2661)
);

BUFx6f_ASAP7_75t_L g2662 ( 
.A(n_2258),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2416),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2432),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2332),
.Y(n_2665)
);

AND2x4_ASAP7_75t_L g2666 ( 
.A(n_2510),
.B(n_1401),
.Y(n_2666)
);

AND2x2_ASAP7_75t_L g2667 ( 
.A(n_2389),
.B(n_1804),
.Y(n_2667)
);

HB1xp67_ASAP7_75t_L g2668 ( 
.A(n_2525),
.Y(n_2668)
);

BUFx6f_ASAP7_75t_L g2669 ( 
.A(n_2259),
.Y(n_2669)
);

BUFx6f_ASAP7_75t_L g2670 ( 
.A(n_2261),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2339),
.Y(n_2671)
);

OR2x2_ASAP7_75t_L g2672 ( 
.A(n_2329),
.B(n_1960),
.Y(n_2672)
);

AND2x2_ASAP7_75t_L g2673 ( 
.A(n_2371),
.B(n_1804),
.Y(n_2673)
);

HB1xp67_ASAP7_75t_L g2674 ( 
.A(n_2560),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2347),
.B(n_1350),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2356),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2364),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2443),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2373),
.Y(n_2679)
);

OA21x2_ASAP7_75t_L g2680 ( 
.A1(n_2415),
.A2(n_1643),
.B(n_1640),
.Y(n_2680)
);

AND2x2_ASAP7_75t_L g2681 ( 
.A(n_2422),
.B(n_1895),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2376),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2452),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2385),
.Y(n_2684)
);

BUFx6f_ASAP7_75t_L g2685 ( 
.A(n_2263),
.Y(n_2685)
);

BUFx2_ASAP7_75t_L g2686 ( 
.A(n_2324),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2377),
.Y(n_2687)
);

CKINVDCx5p33_ASAP7_75t_R g2688 ( 
.A(n_2252),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2460),
.Y(n_2689)
);

AND2x4_ASAP7_75t_L g2690 ( 
.A(n_2265),
.B(n_1403),
.Y(n_2690)
);

OA21x2_ASAP7_75t_L g2691 ( 
.A1(n_2437),
.A2(n_1677),
.B(n_1649),
.Y(n_2691)
);

OAI22xp5_ASAP7_75t_L g2692 ( 
.A1(n_2310),
.A2(n_1294),
.B1(n_1301),
.B2(n_1300),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2388),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2250),
.Y(n_2694)
);

BUFx6f_ASAP7_75t_L g2695 ( 
.A(n_2269),
.Y(n_2695)
);

AND2x4_ASAP7_75t_L g2696 ( 
.A(n_2266),
.B(n_1409),
.Y(n_2696)
);

HB1xp67_ASAP7_75t_L g2697 ( 
.A(n_2290),
.Y(n_2697)
);

AND2x4_ASAP7_75t_L g2698 ( 
.A(n_2394),
.B(n_1411),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2461),
.Y(n_2699)
);

INVx2_ASAP7_75t_L g2700 ( 
.A(n_2478),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2251),
.Y(n_2701)
);

AND2x2_ASAP7_75t_L g2702 ( 
.A(n_2471),
.B(n_1895),
.Y(n_2702)
);

AND2x4_ASAP7_75t_L g2703 ( 
.A(n_2411),
.B(n_1414),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2253),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2479),
.Y(n_2705)
);

INVx3_ASAP7_75t_L g2706 ( 
.A(n_2277),
.Y(n_2706)
);

INVx3_ASAP7_75t_L g2707 ( 
.A(n_2289),
.Y(n_2707)
);

AND2x2_ASAP7_75t_L g2708 ( 
.A(n_2492),
.B(n_1920),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2486),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2267),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2296),
.B(n_1354),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2301),
.B(n_1361),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2297),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2305),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2317),
.B(n_1381),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_L g2716 ( 
.A(n_2317),
.B(n_1382),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2308),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2313),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2496),
.Y(n_2719)
);

AOI22xp5_ASAP7_75t_L g2720 ( 
.A1(n_2352),
.A2(n_1406),
.B1(n_1416),
.B2(n_1405),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2318),
.Y(n_2721)
);

INVxp67_ASAP7_75t_L g2722 ( 
.A(n_2418),
.Y(n_2722)
);

BUFx6f_ASAP7_75t_L g2723 ( 
.A(n_2398),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2323),
.Y(n_2724)
);

HB1xp67_ASAP7_75t_L g2725 ( 
.A(n_2426),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2497),
.Y(n_2726)
);

HB1xp67_ASAP7_75t_L g2727 ( 
.A(n_2446),
.Y(n_2727)
);

BUFx6f_ASAP7_75t_L g2728 ( 
.A(n_2353),
.Y(n_2728)
);

INVx6_ASAP7_75t_L g2729 ( 
.A(n_2374),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2500),
.Y(n_2730)
);

BUFx3_ASAP7_75t_L g2731 ( 
.A(n_2286),
.Y(n_2731)
);

AND2x2_ASAP7_75t_L g2732 ( 
.A(n_2509),
.B(n_1920),
.Y(n_2732)
);

AND2x2_ASAP7_75t_L g2733 ( 
.A(n_2530),
.B(n_1956),
.Y(n_2733)
);

BUFx6f_ASAP7_75t_L g2734 ( 
.A(n_2359),
.Y(n_2734)
);

BUFx6f_ASAP7_75t_L g2735 ( 
.A(n_2365),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2507),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2342),
.B(n_1422),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2519),
.Y(n_2738)
);

AND2x2_ASAP7_75t_L g2739 ( 
.A(n_2555),
.B(n_2557),
.Y(n_2739)
);

INVx2_ASAP7_75t_L g2740 ( 
.A(n_2520),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2563),
.B(n_1426),
.Y(n_2741)
);

INVx1_ASAP7_75t_SL g2742 ( 
.A(n_2322),
.Y(n_2742)
);

OAI22xp5_ASAP7_75t_L g2743 ( 
.A1(n_2424),
.A2(n_1305),
.B1(n_1316),
.B2(n_1310),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2536),
.Y(n_2744)
);

BUFx3_ASAP7_75t_L g2745 ( 
.A(n_2299),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2548),
.Y(n_2746)
);

INVxp67_ASAP7_75t_L g2747 ( 
.A(n_2474),
.Y(n_2747)
);

HB1xp67_ASAP7_75t_L g2748 ( 
.A(n_2494),
.Y(n_2748)
);

BUFx6f_ASAP7_75t_L g2749 ( 
.A(n_2401),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2558),
.Y(n_2750)
);

AND2x6_ASAP7_75t_L g2751 ( 
.A(n_2257),
.B(n_1420),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2561),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2562),
.Y(n_2753)
);

HB1xp67_ASAP7_75t_L g2754 ( 
.A(n_2551),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2568),
.Y(n_2755)
);

BUFx8_ASAP7_75t_L g2756 ( 
.A(n_2246),
.Y(n_2756)
);

BUFx6f_ASAP7_75t_L g2757 ( 
.A(n_2455),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2570),
.Y(n_2758)
);

NOR2xp33_ASAP7_75t_L g2759 ( 
.A(n_2402),
.B(n_1318),
.Y(n_2759)
);

INVx2_ASAP7_75t_L g2760 ( 
.A(n_2262),
.Y(n_2760)
);

CKINVDCx5p33_ASAP7_75t_R g2761 ( 
.A(n_2254),
.Y(n_2761)
);

BUFx2_ASAP7_75t_L g2762 ( 
.A(n_2244),
.Y(n_2762)
);

AOI22xp5_ASAP7_75t_L g2763 ( 
.A1(n_2307),
.A2(n_2451),
.B1(n_2516),
.B2(n_2480),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2363),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2275),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2279),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2327),
.Y(n_2767)
);

BUFx6f_ASAP7_75t_L g2768 ( 
.A(n_2491),
.Y(n_2768)
);

HB1xp67_ASAP7_75t_L g2769 ( 
.A(n_2378),
.Y(n_2769)
);

HB1xp67_ASAP7_75t_L g2770 ( 
.A(n_2396),
.Y(n_2770)
);

OAI22xp5_ASAP7_75t_SL g2771 ( 
.A1(n_2409),
.A2(n_1663),
.B1(n_1755),
.B2(n_1636),
.Y(n_2771)
);

AND2x2_ASAP7_75t_L g2772 ( 
.A(n_2284),
.B(n_1956),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2320),
.B(n_1429),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2255),
.Y(n_2774)
);

AND2x2_ASAP7_75t_L g2775 ( 
.A(n_2447),
.B(n_1319),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2264),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2325),
.B(n_1432),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2280),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2272),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2294),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2288),
.Y(n_2781)
);

INVx6_ASAP7_75t_L g2782 ( 
.A(n_2391),
.Y(n_2782)
);

AND2x2_ASAP7_75t_L g2783 ( 
.A(n_2469),
.B(n_1329),
.Y(n_2783)
);

BUFx2_ASAP7_75t_L g2784 ( 
.A(n_2244),
.Y(n_2784)
);

BUFx6f_ASAP7_75t_L g2785 ( 
.A(n_2410),
.Y(n_2785)
);

AOI22xp5_ASAP7_75t_L g2786 ( 
.A1(n_2533),
.A2(n_1436),
.B1(n_1438),
.B2(n_1433),
.Y(n_2786)
);

BUFx6f_ASAP7_75t_L g2787 ( 
.A(n_2423),
.Y(n_2787)
);

INVx2_ASAP7_75t_L g2788 ( 
.A(n_2291),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2298),
.Y(n_2789)
);

AND2x4_ASAP7_75t_L g2790 ( 
.A(n_2481),
.B(n_1427),
.Y(n_2790)
);

OA21x2_ASAP7_75t_L g2791 ( 
.A1(n_2404),
.A2(n_1696),
.B(n_1683),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2300),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2304),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2312),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2314),
.Y(n_2795)
);

AND2x2_ASAP7_75t_L g2796 ( 
.A(n_2476),
.B(n_2487),
.Y(n_2796)
);

BUFx6f_ASAP7_75t_L g2797 ( 
.A(n_2435),
.Y(n_2797)
);

AND2x2_ASAP7_75t_L g2798 ( 
.A(n_2538),
.B(n_1333),
.Y(n_2798)
);

AND2x4_ASAP7_75t_L g2799 ( 
.A(n_2493),
.B(n_1435),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2441),
.Y(n_2800)
);

INVx2_ASAP7_75t_L g2801 ( 
.A(n_2457),
.Y(n_2801)
);

AND2x6_ASAP7_75t_L g2802 ( 
.A(n_2268),
.B(n_1443),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2475),
.Y(n_2803)
);

NAND2xp33_ASAP7_75t_L g2804 ( 
.A(n_2517),
.B(n_1387),
.Y(n_2804)
);

INVx3_ASAP7_75t_L g2805 ( 
.A(n_2501),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2547),
.Y(n_2806)
);

OAI22xp5_ASAP7_75t_SL g2807 ( 
.A1(n_2413),
.A2(n_1773),
.B1(n_1817),
.B2(n_1771),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2340),
.B(n_1439),
.Y(n_2808)
);

OA21x2_ASAP7_75t_L g2809 ( 
.A1(n_2360),
.A2(n_1768),
.B(n_1722),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2549),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2400),
.Y(n_2811)
);

BUFx6f_ASAP7_75t_L g2812 ( 
.A(n_2505),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2245),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2407),
.Y(n_2814)
);

NOR2xp33_ASAP7_75t_SL g2815 ( 
.A(n_2270),
.B(n_1820),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2370),
.B(n_1442),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2412),
.Y(n_2817)
);

INVx2_ASAP7_75t_L g2818 ( 
.A(n_2419),
.Y(n_2818)
);

NOR2xp33_ASAP7_75t_L g2819 ( 
.A(n_2433),
.B(n_1339),
.Y(n_2819)
);

BUFx8_ASAP7_75t_L g2820 ( 
.A(n_2405),
.Y(n_2820)
);

AND2x2_ASAP7_75t_L g2821 ( 
.A(n_2295),
.B(n_1347),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2430),
.Y(n_2822)
);

INVx3_ASAP7_75t_L g2823 ( 
.A(n_2375),
.Y(n_2823)
);

INVx2_ASAP7_75t_L g2824 ( 
.A(n_2440),
.Y(n_2824)
);

AND2x2_ASAP7_75t_L g2825 ( 
.A(n_2249),
.B(n_1348),
.Y(n_2825)
);

BUFx2_ASAP7_75t_L g2826 ( 
.A(n_2450),
.Y(n_2826)
);

OAI21x1_ASAP7_75t_L g2827 ( 
.A1(n_2309),
.A2(n_1793),
.B(n_1779),
.Y(n_2827)
);

BUFx6f_ASAP7_75t_L g2828 ( 
.A(n_2512),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2456),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2463),
.Y(n_2830)
);

BUFx3_ASAP7_75t_L g2831 ( 
.A(n_2303),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_2473),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2477),
.Y(n_2833)
);

BUFx6f_ASAP7_75t_L g2834 ( 
.A(n_2535),
.Y(n_2834)
);

INVx3_ASAP7_75t_L g2835 ( 
.A(n_2542),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2495),
.Y(n_2836)
);

AND2x2_ASAP7_75t_L g2837 ( 
.A(n_2271),
.B(n_1355),
.Y(n_2837)
);

INVx1_ASAP7_75t_SL g2838 ( 
.A(n_2470),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2431),
.B(n_2553),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2511),
.Y(n_2840)
);

AND3x2_ASAP7_75t_L g2841 ( 
.A(n_2439),
.B(n_1306),
.C(n_1266),
.Y(n_2841)
);

INVx5_ASAP7_75t_L g2842 ( 
.A(n_2450),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2448),
.B(n_1445),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2514),
.Y(n_2844)
);

BUFx6f_ASAP7_75t_L g2845 ( 
.A(n_2566),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2403),
.B(n_1448),
.Y(n_2846)
);

INVx3_ASAP7_75t_L g2847 ( 
.A(n_2567),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2528),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2543),
.Y(n_2849)
);

AND2x2_ASAP7_75t_L g2850 ( 
.A(n_2504),
.B(n_1356),
.Y(n_2850)
);

HB1xp67_ASAP7_75t_L g2851 ( 
.A(n_2383),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2544),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2554),
.B(n_1454),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2559),
.Y(n_2854)
);

AND2x2_ASAP7_75t_L g2855 ( 
.A(n_2541),
.B(n_1357),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2382),
.Y(n_2856)
);

INVx3_ASAP7_75t_L g2857 ( 
.A(n_2343),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2390),
.Y(n_2858)
);

BUFx2_ASAP7_75t_L g2859 ( 
.A(n_2523),
.Y(n_2859)
);

AND2x4_ASAP7_75t_L g2860 ( 
.A(n_2565),
.B(n_1451),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_2552),
.B(n_1455),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2390),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2523),
.Y(n_2863)
);

AND2x2_ASAP7_75t_L g2864 ( 
.A(n_2417),
.B(n_1358),
.Y(n_2864)
);

BUFx6f_ASAP7_75t_L g2865 ( 
.A(n_2468),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2428),
.B(n_1468),
.Y(n_2866)
);

CKINVDCx5p33_ASAP7_75t_R g2867 ( 
.A(n_2414),
.Y(n_2867)
);

AOI22xp5_ASAP7_75t_L g2868 ( 
.A1(n_2467),
.A2(n_1481),
.B1(n_1482),
.B2(n_1474),
.Y(n_2868)
);

INVx2_ASAP7_75t_L g2869 ( 
.A(n_2316),
.Y(n_2869)
);

BUFx8_ASAP7_75t_L g2870 ( 
.A(n_2429),
.Y(n_2870)
);

INVx3_ASAP7_75t_L g2871 ( 
.A(n_2274),
.Y(n_2871)
);

INVx3_ASAP7_75t_L g2872 ( 
.A(n_2335),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2518),
.Y(n_2873)
);

BUFx6f_ASAP7_75t_L g2874 ( 
.A(n_2341),
.Y(n_2874)
);

AND3x2_ASAP7_75t_L g2875 ( 
.A(n_2539),
.B(n_1370),
.C(n_1344),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2436),
.Y(n_2876)
);

OAI21x1_ASAP7_75t_L g2877 ( 
.A1(n_2369),
.A2(n_1822),
.B(n_1811),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2442),
.Y(n_2878)
);

NAND2xp33_ASAP7_75t_L g2879 ( 
.A(n_2387),
.B(n_1387),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2444),
.B(n_1483),
.Y(n_2880)
);

BUFx3_ASAP7_75t_L g2881 ( 
.A(n_2367),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2449),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2484),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2499),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2503),
.Y(n_2885)
);

BUFx6f_ASAP7_75t_L g2886 ( 
.A(n_2573),
.Y(n_2886)
);

AND2x2_ASAP7_75t_L g2887 ( 
.A(n_2634),
.B(n_2379),
.Y(n_2887)
);

NOR2xp33_ASAP7_75t_L g2888 ( 
.A(n_2759),
.B(n_2521),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_SL g2889 ( 
.A(n_2842),
.B(n_1495),
.Y(n_2889)
);

NOR2xp33_ASAP7_75t_L g2890 ( 
.A(n_2633),
.B(n_2529),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_SL g2891 ( 
.A(n_2842),
.B(n_1497),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2572),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2576),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2577),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_2659),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2642),
.B(n_1854),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2661),
.Y(n_2897)
);

INVx3_ASAP7_75t_L g2898 ( 
.A(n_2573),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2590),
.B(n_1856),
.Y(n_2899)
);

NOR2xp33_ASAP7_75t_L g2900 ( 
.A(n_2592),
.B(n_2537),
.Y(n_2900)
);

INVx3_ASAP7_75t_L g2901 ( 
.A(n_2574),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2663),
.Y(n_2902)
);

AOI22xp5_ASAP7_75t_L g2903 ( 
.A1(n_2643),
.A2(n_1500),
.B1(n_1507),
.B2(n_1501),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2585),
.B(n_1864),
.Y(n_2904)
);

INVx1_ASAP7_75t_SL g2905 ( 
.A(n_2742),
.Y(n_2905)
);

INVxp33_ASAP7_75t_L g2906 ( 
.A(n_2603),
.Y(n_2906)
);

CKINVDCx6p67_ASAP7_75t_R g2907 ( 
.A(n_2593),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2679),
.Y(n_2908)
);

INVx2_ASAP7_75t_L g2909 ( 
.A(n_2664),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2682),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2678),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2683),
.Y(n_2912)
);

AND2x2_ASAP7_75t_L g2913 ( 
.A(n_2594),
.B(n_2652),
.Y(n_2913)
);

INVxp67_ASAP7_75t_SL g2914 ( 
.A(n_2749),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2694),
.Y(n_2915)
);

BUFx2_ASAP7_75t_L g2916 ( 
.A(n_2575),
.Y(n_2916)
);

AND3x2_ASAP7_75t_L g2917 ( 
.A(n_2762),
.B(n_1424),
.C(n_1389),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_2620),
.B(n_1868),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2701),
.Y(n_2919)
);

INVx3_ASAP7_75t_L g2920 ( 
.A(n_2574),
.Y(n_2920)
);

INVx2_ASAP7_75t_L g2921 ( 
.A(n_2689),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2699),
.Y(n_2922)
);

AND3x2_ASAP7_75t_L g2923 ( 
.A(n_2784),
.B(n_1566),
.C(n_1546),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2704),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2710),
.Y(n_2925)
);

AND2x2_ASAP7_75t_SL g2926 ( 
.A(n_2815),
.B(n_2354),
.Y(n_2926)
);

INVx2_ASAP7_75t_L g2927 ( 
.A(n_2700),
.Y(n_2927)
);

INVx2_ASAP7_75t_L g2928 ( 
.A(n_2705),
.Y(n_2928)
);

INVxp67_ASAP7_75t_SL g2929 ( 
.A(n_2749),
.Y(n_2929)
);

NOR2xp33_ASAP7_75t_L g2930 ( 
.A(n_2622),
.B(n_2420),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2709),
.Y(n_2931)
);

NAND2xp5_ASAP7_75t_L g2932 ( 
.A(n_2739),
.B(n_1885),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_SL g2933 ( 
.A(n_2597),
.B(n_2667),
.Y(n_2933)
);

BUFx10_ASAP7_75t_L g2934 ( 
.A(n_2867),
.Y(n_2934)
);

INVx2_ASAP7_75t_L g2935 ( 
.A(n_2719),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_2726),
.Y(n_2936)
);

AND2x6_ASAP7_75t_L g2937 ( 
.A(n_2673),
.B(n_2647),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2713),
.Y(n_2938)
);

AND2x2_ASAP7_75t_L g2939 ( 
.A(n_2681),
.B(n_1821),
.Y(n_2939)
);

INVx2_ASAP7_75t_L g2940 ( 
.A(n_2736),
.Y(n_2940)
);

INVx5_ASAP7_75t_L g2941 ( 
.A(n_2865),
.Y(n_2941)
);

INVx5_ASAP7_75t_L g2942 ( 
.A(n_2865),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2740),
.Y(n_2943)
);

CKINVDCx6p67_ASAP7_75t_R g2944 ( 
.A(n_2731),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_SL g2945 ( 
.A(n_2819),
.B(n_1517),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2605),
.B(n_1910),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_SL g2947 ( 
.A(n_2821),
.B(n_1527),
.Y(n_2947)
);

AO21x2_ASAP7_75t_L g2948 ( 
.A1(n_2839),
.A2(n_1941),
.B(n_1917),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2750),
.Y(n_2949)
);

INVx1_ASAP7_75t_SL g2950 ( 
.A(n_2838),
.Y(n_2950)
);

AND2x2_ASAP7_75t_L g2951 ( 
.A(n_2702),
.B(n_1828),
.Y(n_2951)
);

INVx2_ASAP7_75t_L g2952 ( 
.A(n_2760),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2714),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2717),
.Y(n_2954)
);

INVx2_ASAP7_75t_L g2955 ( 
.A(n_2765),
.Y(n_2955)
);

INVx2_ASAP7_75t_SL g2956 ( 
.A(n_2769),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2718),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2721),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2724),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2730),
.Y(n_2960)
);

AND3x2_ASAP7_75t_L g2961 ( 
.A(n_2826),
.B(n_1653),
.C(n_1567),
.Y(n_2961)
);

INVx2_ASAP7_75t_L g2962 ( 
.A(n_2766),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2778),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_SL g2964 ( 
.A(n_2723),
.B(n_2591),
.Y(n_2964)
);

NAND3xp33_ASAP7_75t_L g2965 ( 
.A(n_2720),
.B(n_1369),
.C(n_1364),
.Y(n_2965)
);

INVxp67_ASAP7_75t_L g2966 ( 
.A(n_2623),
.Y(n_2966)
);

AO21x2_ASAP7_75t_L g2967 ( 
.A1(n_2711),
.A2(n_1954),
.B(n_1950),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2738),
.Y(n_2968)
);

INVx3_ASAP7_75t_L g2969 ( 
.A(n_2582),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2744),
.Y(n_2970)
);

INVx2_ASAP7_75t_L g2971 ( 
.A(n_2781),
.Y(n_2971)
);

BUFx3_ASAP7_75t_L g2972 ( 
.A(n_2662),
.Y(n_2972)
);

INVx2_ASAP7_75t_L g2973 ( 
.A(n_2788),
.Y(n_2973)
);

AND2x2_ASAP7_75t_SL g2974 ( 
.A(n_2859),
.B(n_2445),
.Y(n_2974)
);

NAND3xp33_ASAP7_75t_L g2975 ( 
.A(n_2868),
.B(n_1374),
.C(n_1372),
.Y(n_2975)
);

NAND3xp33_ASAP7_75t_L g2976 ( 
.A(n_2786),
.B(n_1376),
.C(n_1375),
.Y(n_2976)
);

INVx2_ASAP7_75t_SL g2977 ( 
.A(n_2770),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2746),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2752),
.Y(n_2979)
);

NAND3xp33_ASAP7_75t_L g2980 ( 
.A(n_2866),
.B(n_2672),
.C(n_2879),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_SL g2981 ( 
.A(n_2723),
.B(n_1536),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2638),
.B(n_1968),
.Y(n_2982)
);

INVx2_ASAP7_75t_L g2983 ( 
.A(n_2789),
.Y(n_2983)
);

INVx2_ASAP7_75t_L g2984 ( 
.A(n_2792),
.Y(n_2984)
);

OAI22xp33_ASAP7_75t_SL g2985 ( 
.A1(n_2858),
.A2(n_1973),
.B1(n_1987),
.B2(n_1971),
.Y(n_2985)
);

INVx2_ASAP7_75t_L g2986 ( 
.A(n_2817),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2818),
.Y(n_2987)
);

INVx2_ASAP7_75t_L g2988 ( 
.A(n_2824),
.Y(n_2988)
);

NOR2xp33_ASAP7_75t_L g2989 ( 
.A(n_2861),
.B(n_2453),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2753),
.Y(n_2990)
);

INVx2_ASAP7_75t_SL g2991 ( 
.A(n_2581),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2639),
.B(n_2003),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2832),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2848),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2849),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2660),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2644),
.B(n_2024),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2755),
.Y(n_2998)
);

BUFx10_ASAP7_75t_L g2999 ( 
.A(n_2874),
.Y(n_2999)
);

AOI22xp33_ASAP7_75t_SL g3000 ( 
.A1(n_2771),
.A2(n_2569),
.B1(n_1836),
.B2(n_2007),
.Y(n_3000)
);

NAND2xp33_ASAP7_75t_L g3001 ( 
.A(n_2712),
.B(n_1540),
.Y(n_3001)
);

AOI22xp33_ASAP7_75t_L g3002 ( 
.A1(n_2698),
.A2(n_2044),
.B1(n_2067),
.B2(n_2047),
.Y(n_3002)
);

AOI21x1_ASAP7_75t_L g3003 ( 
.A1(n_2816),
.A2(n_1476),
.B(n_1461),
.Y(n_3003)
);

BUFx4f_ASAP7_75t_L g3004 ( 
.A(n_2874),
.Y(n_3004)
);

AOI22xp33_ASAP7_75t_L g3005 ( 
.A1(n_2645),
.A2(n_1336),
.B1(n_1741),
.B2(n_1738),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2665),
.Y(n_3006)
);

AND2x4_ASAP7_75t_L g3007 ( 
.A(n_2579),
.B(n_1491),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2758),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2655),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2658),
.B(n_1556),
.Y(n_3010)
);

NOR2xp33_ASAP7_75t_L g3011 ( 
.A(n_2722),
.B(n_2458),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2684),
.Y(n_3012)
);

AND2x2_ASAP7_75t_L g3013 ( 
.A(n_2708),
.B(n_1883),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_2671),
.Y(n_3014)
);

INVx2_ASAP7_75t_L g3015 ( 
.A(n_2676),
.Y(n_3015)
);

BUFx3_ASAP7_75t_L g3016 ( 
.A(n_2662),
.Y(n_3016)
);

INVx3_ASAP7_75t_L g3017 ( 
.A(n_2582),
.Y(n_3017)
);

OAI22x1_ASAP7_75t_L g3018 ( 
.A1(n_2656),
.A2(n_2513),
.B1(n_1379),
.B2(n_1383),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_SL g3019 ( 
.A(n_2862),
.B(n_1563),
.Y(n_3019)
);

NAND2xp33_ASAP7_75t_L g3020 ( 
.A(n_2812),
.B(n_1573),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2813),
.Y(n_3021)
);

AOI22xp5_ASAP7_75t_L g3022 ( 
.A1(n_2863),
.A2(n_1575),
.B1(n_1589),
.B2(n_1577),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2675),
.B(n_1596),
.Y(n_3023)
);

INVx3_ASAP7_75t_L g3024 ( 
.A(n_2587),
.Y(n_3024)
);

INVx2_ASAP7_75t_L g3025 ( 
.A(n_2801),
.Y(n_3025)
);

INVx2_ASAP7_75t_L g3026 ( 
.A(n_2810),
.Y(n_3026)
);

OAI22xp33_ASAP7_75t_L g3027 ( 
.A1(n_2846),
.A2(n_2019),
.B1(n_2020),
.B2(n_2015),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2814),
.Y(n_3028)
);

BUFx6f_ASAP7_75t_L g3029 ( 
.A(n_2587),
.Y(n_3029)
);

INVx2_ASAP7_75t_L g3030 ( 
.A(n_2822),
.Y(n_3030)
);

INVx4_ASAP7_75t_L g3031 ( 
.A(n_2669),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_SL g3032 ( 
.A(n_2732),
.B(n_1604),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2829),
.Y(n_3033)
);

INVx2_ASAP7_75t_L g3034 ( 
.A(n_2830),
.Y(n_3034)
);

NOR2xp33_ASAP7_75t_L g3035 ( 
.A(n_2747),
.B(n_1378),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2833),
.Y(n_3036)
);

CKINVDCx5p33_ASAP7_75t_R g3037 ( 
.A(n_2688),
.Y(n_3037)
);

INVx2_ASAP7_75t_L g3038 ( 
.A(n_2836),
.Y(n_3038)
);

INVx2_ASAP7_75t_L g3039 ( 
.A(n_2840),
.Y(n_3039)
);

BUFx6f_ASAP7_75t_L g3040 ( 
.A(n_2589),
.Y(n_3040)
);

AOI22xp5_ASAP7_75t_L g3041 ( 
.A1(n_2860),
.A2(n_1607),
.B1(n_1630),
.B2(n_1619),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2844),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2852),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2854),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_SL g3045 ( 
.A(n_2733),
.B(n_2812),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_L g3046 ( 
.A(n_2741),
.B(n_2649),
.Y(n_3046)
);

INVx1_ASAP7_75t_SL g3047 ( 
.A(n_2697),
.Y(n_3047)
);

NAND2xp33_ASAP7_75t_R g3048 ( 
.A(n_2761),
.B(n_1639),
.Y(n_3048)
);

BUFx6f_ASAP7_75t_L g3049 ( 
.A(n_2589),
.Y(n_3049)
);

INVx2_ASAP7_75t_L g3050 ( 
.A(n_2793),
.Y(n_3050)
);

INVx2_ASAP7_75t_SL g3051 ( 
.A(n_2725),
.Y(n_3051)
);

CKINVDCx14_ASAP7_75t_R g3052 ( 
.A(n_2648),
.Y(n_3052)
);

NAND3xp33_ASAP7_75t_L g3053 ( 
.A(n_2692),
.B(n_1392),
.C(n_1384),
.Y(n_3053)
);

INVx3_ASAP7_75t_L g3054 ( 
.A(n_2600),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_2794),
.Y(n_3055)
);

INVx2_ASAP7_75t_L g3056 ( 
.A(n_2795),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2805),
.Y(n_3057)
);

NOR2xp33_ASAP7_75t_L g3058 ( 
.A(n_2610),
.B(n_1395),
.Y(n_3058)
);

AND2x6_ASAP7_75t_L g3059 ( 
.A(n_2757),
.B(n_1428),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2800),
.Y(n_3060)
);

INVx5_ASAP7_75t_L g3061 ( 
.A(n_2586),
.Y(n_3061)
);

INVx2_ASAP7_75t_L g3062 ( 
.A(n_2803),
.Y(n_3062)
);

INVx8_ASAP7_75t_L g3063 ( 
.A(n_2586),
.Y(n_3063)
);

BUFx2_ASAP7_75t_L g3064 ( 
.A(n_2653),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2806),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_SL g3066 ( 
.A(n_2828),
.B(n_1650),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2693),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2774),
.Y(n_3068)
);

INVx4_ASAP7_75t_L g3069 ( 
.A(n_2669),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2785),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2776),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_SL g3072 ( 
.A(n_2828),
.B(n_1656),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_2785),
.Y(n_3073)
);

OAI21xp5_ASAP7_75t_L g3074 ( 
.A1(n_2827),
.A2(n_1660),
.B(n_1659),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_SL g3075 ( 
.A(n_2834),
.B(n_1661),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2779),
.Y(n_3076)
);

BUFx3_ASAP7_75t_L g3077 ( 
.A(n_2670),
.Y(n_3077)
);

NAND3xp33_ASAP7_75t_L g3078 ( 
.A(n_2743),
.B(n_1397),
.C(n_1396),
.Y(n_3078)
);

BUFx6f_ASAP7_75t_L g3079 ( 
.A(n_2600),
.Y(n_3079)
);

AOI22xp33_ASAP7_75t_L g3080 ( 
.A1(n_2791),
.A2(n_1336),
.B1(n_1880),
.B2(n_1855),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2780),
.Y(n_3081)
);

INVx2_ASAP7_75t_L g3082 ( 
.A(n_2787),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2767),
.Y(n_3083)
);

NOR2xp33_ASAP7_75t_R g3084 ( 
.A(n_2871),
.B(n_1665),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_L g3085 ( 
.A(n_2651),
.B(n_1678),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2787),
.Y(n_3086)
);

CKINVDCx5p33_ASAP7_75t_R g3087 ( 
.A(n_2763),
.Y(n_3087)
);

INVx2_ASAP7_75t_L g3088 ( 
.A(n_2797),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2797),
.Y(n_3089)
);

AOI21x1_ASAP7_75t_L g3090 ( 
.A1(n_2654),
.A2(n_1510),
.B(n_1496),
.Y(n_3090)
);

CKINVDCx5p33_ASAP7_75t_R g3091 ( 
.A(n_2881),
.Y(n_3091)
);

BUFx6f_ASAP7_75t_SL g3092 ( 
.A(n_2745),
.Y(n_3092)
);

CKINVDCx20_ASAP7_75t_R g3093 ( 
.A(n_2608),
.Y(n_3093)
);

INVx3_ASAP7_75t_L g3094 ( 
.A(n_2626),
.Y(n_3094)
);

AO22x2_ASAP7_75t_L g3095 ( 
.A1(n_2807),
.A2(n_1521),
.B1(n_1522),
.B2(n_1514),
.Y(n_3095)
);

NOR2xp33_ASAP7_75t_L g3096 ( 
.A(n_2687),
.B(n_1400),
.Y(n_3096)
);

INVx2_ASAP7_75t_L g3097 ( 
.A(n_2757),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2604),
.B(n_1681),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2677),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2578),
.Y(n_3100)
);

NOR2xp33_ASAP7_75t_L g3101 ( 
.A(n_2864),
.B(n_1402),
.Y(n_3101)
);

BUFx6f_ASAP7_75t_L g3102 ( 
.A(n_2626),
.Y(n_3102)
);

INVxp67_ASAP7_75t_SL g3103 ( 
.A(n_2636),
.Y(n_3103)
);

AOI22xp33_ASAP7_75t_L g3104 ( 
.A1(n_2809),
.A2(n_1336),
.B1(n_1904),
.B2(n_1892),
.Y(n_3104)
);

NOR2x1p5_ASAP7_75t_L g3105 ( 
.A(n_2872),
.B(n_1404),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2599),
.Y(n_3106)
);

INVxp33_ASAP7_75t_L g3107 ( 
.A(n_2727),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_SL g3108 ( 
.A(n_2834),
.B(n_1684),
.Y(n_3108)
);

BUFx2_ASAP7_75t_L g3109 ( 
.A(n_2748),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_2768),
.Y(n_3110)
);

AOI22xp33_ASAP7_75t_SL g3111 ( 
.A1(n_2857),
.A2(n_2050),
.B1(n_2059),
.B2(n_1336),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_SL g3112 ( 
.A(n_2845),
.B(n_1688),
.Y(n_3112)
);

INVxp33_ASAP7_75t_L g3113 ( 
.A(n_2754),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2601),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2609),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2613),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2768),
.Y(n_3117)
);

NAND2xp33_ASAP7_75t_L g3118 ( 
.A(n_2845),
.B(n_1690),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2614),
.Y(n_3119)
);

XNOR2x2_ASAP7_75t_SL g3120 ( 
.A(n_2825),
.B(n_1524),
.Y(n_3120)
);

BUFx6f_ASAP7_75t_L g3121 ( 
.A(n_2636),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_SL g3122 ( 
.A(n_2728),
.B(n_2734),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2618),
.Y(n_3123)
);

INVx2_ASAP7_75t_L g3124 ( 
.A(n_2580),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_2625),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_2583),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2615),
.B(n_1692),
.Y(n_3127)
);

OAI22xp33_ASAP7_75t_L g3128 ( 
.A1(n_2835),
.A2(n_1531),
.B1(n_1538),
.B2(n_1526),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_3046),
.B(n_2843),
.Y(n_3129)
);

NOR2x1p5_ASAP7_75t_L g3130 ( 
.A(n_2944),
.B(n_2831),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_SL g3131 ( 
.A(n_2913),
.B(n_2728),
.Y(n_3131)
);

AND2x4_ASAP7_75t_L g3132 ( 
.A(n_2941),
.B(n_2584),
.Y(n_3132)
);

INVx5_ASAP7_75t_L g3133 ( 
.A(n_2999),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2892),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2893),
.Y(n_3135)
);

INVx2_ASAP7_75t_L g3136 ( 
.A(n_2895),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_2914),
.B(n_2811),
.Y(n_3137)
);

BUFx3_ASAP7_75t_L g3138 ( 
.A(n_2886),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_SL g3139 ( 
.A(n_2980),
.B(n_2734),
.Y(n_3139)
);

INVx3_ASAP7_75t_L g3140 ( 
.A(n_2886),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_2929),
.B(n_2823),
.Y(n_3141)
);

NOR2xp33_ASAP7_75t_L g3142 ( 
.A(n_2966),
.B(n_2611),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_2899),
.B(n_2904),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2894),
.Y(n_3144)
);

AND2x2_ASAP7_75t_L g3145 ( 
.A(n_2905),
.B(n_2837),
.Y(n_3145)
);

AND2x4_ASAP7_75t_L g3146 ( 
.A(n_2941),
.B(n_2588),
.Y(n_3146)
);

INVx3_ASAP7_75t_L g3147 ( 
.A(n_3029),
.Y(n_3147)
);

AND2x2_ASAP7_75t_L g3148 ( 
.A(n_2939),
.B(n_2850),
.Y(n_3148)
);

AOI22xp5_ASAP7_75t_L g3149 ( 
.A1(n_2937),
.A2(n_2737),
.B1(n_2853),
.B2(n_2847),
.Y(n_3149)
);

AND2x2_ASAP7_75t_L g3150 ( 
.A(n_2951),
.B(n_2855),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_2908),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2910),
.Y(n_3152)
);

INVx2_ASAP7_75t_L g3153 ( 
.A(n_2897),
.Y(n_3153)
);

INVx3_ASAP7_75t_L g3154 ( 
.A(n_3029),
.Y(n_3154)
);

OR2x2_ASAP7_75t_L g3155 ( 
.A(n_3047),
.B(n_2616),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_2915),
.Y(n_3156)
);

OR2x6_ASAP7_75t_L g3157 ( 
.A(n_3063),
.B(n_2612),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2919),
.Y(n_3158)
);

INVx2_ASAP7_75t_L g3159 ( 
.A(n_2902),
.Y(n_3159)
);

BUFx6f_ASAP7_75t_L g3160 ( 
.A(n_3040),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2924),
.Y(n_3161)
);

NAND3x1_ASAP7_75t_L g3162 ( 
.A(n_3011),
.B(n_2878),
.C(n_2876),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_SL g3163 ( 
.A(n_2956),
.B(n_2977),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2925),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_2938),
.Y(n_3165)
);

NOR2xp33_ASAP7_75t_L g3166 ( 
.A(n_3107),
.B(n_2650),
.Y(n_3166)
);

INVx3_ASAP7_75t_L g3167 ( 
.A(n_3040),
.Y(n_3167)
);

INVx2_ASAP7_75t_L g3168 ( 
.A(n_2909),
.Y(n_3168)
);

INVx2_ASAP7_75t_L g3169 ( 
.A(n_2911),
.Y(n_3169)
);

AND2x6_ASAP7_75t_L g3170 ( 
.A(n_2887),
.B(n_2869),
.Y(n_3170)
);

BUFx3_ASAP7_75t_L g3171 ( 
.A(n_3049),
.Y(n_3171)
);

AND3x4_ASAP7_75t_L g3172 ( 
.A(n_2972),
.B(n_2607),
.C(n_2595),
.Y(n_3172)
);

AND2x6_ASAP7_75t_L g3173 ( 
.A(n_2900),
.B(n_2882),
.Y(n_3173)
);

CKINVDCx16_ASAP7_75t_R g3174 ( 
.A(n_3093),
.Y(n_3174)
);

NOR2xp33_ASAP7_75t_L g3175 ( 
.A(n_3113),
.B(n_2668),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2953),
.Y(n_3176)
);

AOI22xp5_ASAP7_75t_L g3177 ( 
.A1(n_2937),
.A2(n_2764),
.B1(n_2690),
.B2(n_2696),
.Y(n_3177)
);

NAND2x1p5_ASAP7_75t_L g3178 ( 
.A(n_2942),
.B(n_3031),
.Y(n_3178)
);

BUFx4f_ASAP7_75t_L g3179 ( 
.A(n_2907),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2954),
.Y(n_3180)
);

BUFx6f_ASAP7_75t_L g3181 ( 
.A(n_3049),
.Y(n_3181)
);

INVx2_ASAP7_75t_L g3182 ( 
.A(n_2912),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_L g3183 ( 
.A(n_2918),
.B(n_2775),
.Y(n_3183)
);

BUFx6f_ASAP7_75t_L g3184 ( 
.A(n_3079),
.Y(n_3184)
);

INVx2_ASAP7_75t_L g3185 ( 
.A(n_2921),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2957),
.Y(n_3186)
);

AOI22xp5_ASAP7_75t_L g3187 ( 
.A1(n_2937),
.A2(n_2802),
.B1(n_2703),
.B2(n_2799),
.Y(n_3187)
);

AND2x4_ASAP7_75t_L g3188 ( 
.A(n_2942),
.B(n_2596),
.Y(n_3188)
);

INVxp67_ASAP7_75t_L g3189 ( 
.A(n_3109),
.Y(n_3189)
);

BUFx3_ASAP7_75t_L g3190 ( 
.A(n_3079),
.Y(n_3190)
);

NOR2xp33_ASAP7_75t_L g3191 ( 
.A(n_2906),
.B(n_2674),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_L g3192 ( 
.A(n_2896),
.B(n_2783),
.Y(n_3192)
);

INVx2_ASAP7_75t_SL g3193 ( 
.A(n_3051),
.Y(n_3193)
);

NAND2x1p5_ASAP7_75t_L g3194 ( 
.A(n_3069),
.B(n_2637),
.Y(n_3194)
);

INVx4_ASAP7_75t_L g3195 ( 
.A(n_3102),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2958),
.Y(n_3196)
);

AND2x2_ASAP7_75t_L g3197 ( 
.A(n_3013),
.B(n_2772),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_L g3198 ( 
.A(n_2946),
.B(n_2798),
.Y(n_3198)
);

INVxp67_ASAP7_75t_L g3199 ( 
.A(n_3064),
.Y(n_3199)
);

INVx2_ASAP7_75t_L g3200 ( 
.A(n_2922),
.Y(n_3200)
);

INVx5_ASAP7_75t_L g3201 ( 
.A(n_3102),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_2959),
.Y(n_3202)
);

INVx2_ASAP7_75t_L g3203 ( 
.A(n_2927),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_3009),
.Y(n_3204)
);

AND2x4_ASAP7_75t_L g3205 ( 
.A(n_3016),
.B(n_2602),
.Y(n_3205)
);

INVx2_ASAP7_75t_L g3206 ( 
.A(n_2928),
.Y(n_3206)
);

NOR2xp33_ASAP7_75t_SL g3207 ( 
.A(n_3037),
.B(n_3004),
.Y(n_3207)
);

INVx2_ASAP7_75t_L g3208 ( 
.A(n_2931),
.Y(n_3208)
);

AND2x4_ASAP7_75t_L g3209 ( 
.A(n_3077),
.B(n_2606),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_3021),
.Y(n_3210)
);

INVx4_ASAP7_75t_SL g3211 ( 
.A(n_3092),
.Y(n_3211)
);

NAND3xp33_ASAP7_75t_L g3212 ( 
.A(n_3035),
.B(n_2875),
.C(n_2666),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_3028),
.Y(n_3213)
);

INVx4_ASAP7_75t_L g3214 ( 
.A(n_3121),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_3033),
.Y(n_3215)
);

INVx2_ASAP7_75t_L g3216 ( 
.A(n_2935),
.Y(n_3216)
);

INVx4_ASAP7_75t_L g3217 ( 
.A(n_3121),
.Y(n_3217)
);

INVx3_ASAP7_75t_L g3218 ( 
.A(n_2898),
.Y(n_3218)
);

BUFx3_ASAP7_75t_L g3219 ( 
.A(n_2916),
.Y(n_3219)
);

INVx2_ASAP7_75t_L g3220 ( 
.A(n_2936),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_3101),
.B(n_2790),
.Y(n_3221)
);

INVx2_ASAP7_75t_SL g3222 ( 
.A(n_2950),
.Y(n_3222)
);

INVx2_ASAP7_75t_L g3223 ( 
.A(n_2940),
.Y(n_3223)
);

OR2x2_ASAP7_75t_L g3224 ( 
.A(n_2932),
.B(n_2624),
.Y(n_3224)
);

BUFx6f_ASAP7_75t_L g3225 ( 
.A(n_2901),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_3042),
.Y(n_3226)
);

INVx2_ASAP7_75t_L g3227 ( 
.A(n_2943),
.Y(n_3227)
);

INVx3_ASAP7_75t_L g3228 ( 
.A(n_2920),
.Y(n_3228)
);

OAI22xp5_ASAP7_75t_L g3229 ( 
.A1(n_3097),
.A2(n_2735),
.B1(n_2880),
.B2(n_2851),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_3044),
.Y(n_3230)
);

AND2x2_ASAP7_75t_SL g3231 ( 
.A(n_2926),
.B(n_2686),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_2960),
.Y(n_3232)
);

AND2x2_ASAP7_75t_L g3233 ( 
.A(n_3058),
.B(n_2796),
.Y(n_3233)
);

AND2x4_ASAP7_75t_L g3234 ( 
.A(n_2991),
.B(n_2617),
.Y(n_3234)
);

AND2x4_ASAP7_75t_L g3235 ( 
.A(n_3070),
.B(n_2621),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_2968),
.Y(n_3236)
);

BUFx6f_ASAP7_75t_L g3237 ( 
.A(n_2969),
.Y(n_3237)
);

BUFx10_ASAP7_75t_L g3238 ( 
.A(n_2888),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2970),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_2949),
.Y(n_3240)
);

NAND2xp33_ASAP7_75t_L g3241 ( 
.A(n_3059),
.B(n_2735),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_2978),
.Y(n_3242)
);

NOR2xp33_ASAP7_75t_L g3243 ( 
.A(n_3027),
.B(n_2890),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2979),
.Y(n_3244)
);

AOI22xp5_ASAP7_75t_L g3245 ( 
.A1(n_2933),
.A2(n_2802),
.B1(n_2751),
.B2(n_2804),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_SL g3246 ( 
.A(n_3061),
.B(n_2670),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_2990),
.Y(n_3247)
);

INVxp67_ASAP7_75t_SL g3248 ( 
.A(n_3110),
.Y(n_3248)
);

BUFx6f_ASAP7_75t_L g3249 ( 
.A(n_3017),
.Y(n_3249)
);

AND2x2_ASAP7_75t_L g3250 ( 
.A(n_3096),
.B(n_2635),
.Y(n_3250)
);

INVx4_ASAP7_75t_L g3251 ( 
.A(n_3091),
.Y(n_3251)
);

NOR2xp33_ASAP7_75t_L g3252 ( 
.A(n_3087),
.B(n_2873),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_2998),
.Y(n_3253)
);

AND2x2_ASAP7_75t_L g3254 ( 
.A(n_3061),
.B(n_2641),
.Y(n_3254)
);

INVx2_ASAP7_75t_SL g3255 ( 
.A(n_3007),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_3008),
.Y(n_3256)
);

BUFx3_ASAP7_75t_L g3257 ( 
.A(n_3024),
.Y(n_3257)
);

BUFx2_ASAP7_75t_L g3258 ( 
.A(n_3095),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_3012),
.Y(n_3259)
);

BUFx6f_ASAP7_75t_L g3260 ( 
.A(n_3054),
.Y(n_3260)
);

BUFx6f_ASAP7_75t_L g3261 ( 
.A(n_3094),
.Y(n_3261)
);

INVx4_ASAP7_75t_L g3262 ( 
.A(n_2934),
.Y(n_3262)
);

AND2x2_ASAP7_75t_L g3263 ( 
.A(n_2964),
.B(n_2627),
.Y(n_3263)
);

NOR2xp33_ASAP7_75t_L g3264 ( 
.A(n_2930),
.B(n_2598),
.Y(n_3264)
);

AO22x2_ASAP7_75t_L g3265 ( 
.A1(n_3120),
.A2(n_1545),
.B1(n_1548),
.B2(n_1539),
.Y(n_3265)
);

BUFx3_ASAP7_75t_L g3266 ( 
.A(n_3073),
.Y(n_3266)
);

BUFx6f_ASAP7_75t_L g3267 ( 
.A(n_3082),
.Y(n_3267)
);

INVx3_ASAP7_75t_L g3268 ( 
.A(n_3088),
.Y(n_3268)
);

AND2x4_ASAP7_75t_L g3269 ( 
.A(n_3103),
.B(n_2619),
.Y(n_3269)
);

NAND2x1p5_ASAP7_75t_L g3270 ( 
.A(n_3122),
.B(n_2637),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_2952),
.Y(n_3271)
);

INVx2_ASAP7_75t_L g3272 ( 
.A(n_2955),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_2962),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_L g3274 ( 
.A(n_3085),
.B(n_2715),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_2963),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_2971),
.Y(n_3276)
);

AND2x4_ASAP7_75t_L g3277 ( 
.A(n_3086),
.B(n_2631),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_2973),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_2983),
.Y(n_3279)
);

INVxp67_ASAP7_75t_L g3280 ( 
.A(n_3032),
.Y(n_3280)
);

NAND3x1_ASAP7_75t_L g3281 ( 
.A(n_2989),
.B(n_2884),
.C(n_2883),
.Y(n_3281)
);

INVx3_ASAP7_75t_L g3282 ( 
.A(n_3062),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_2984),
.Y(n_3283)
);

NOR2xp33_ASAP7_75t_L g3284 ( 
.A(n_2975),
.B(n_2630),
.Y(n_3284)
);

BUFx4f_ASAP7_75t_L g3285 ( 
.A(n_3063),
.Y(n_3285)
);

INVx2_ASAP7_75t_L g3286 ( 
.A(n_2996),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_3006),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_3098),
.B(n_2716),
.Y(n_3288)
);

INVx4_ASAP7_75t_L g3289 ( 
.A(n_2917),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_3014),
.Y(n_3290)
);

INVx2_ASAP7_75t_L g3291 ( 
.A(n_3136),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_L g3292 ( 
.A(n_3129),
.B(n_3030),
.Y(n_3292)
);

AND2x2_ASAP7_75t_L g3293 ( 
.A(n_3145),
.B(n_3148),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_SL g3294 ( 
.A(n_3221),
.B(n_3150),
.Y(n_3294)
);

INVx2_ASAP7_75t_L g3295 ( 
.A(n_3153),
.Y(n_3295)
);

OR2x6_ASAP7_75t_L g3296 ( 
.A(n_3222),
.B(n_3219),
.Y(n_3296)
);

CKINVDCx11_ASAP7_75t_R g3297 ( 
.A(n_3211),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_SL g3298 ( 
.A(n_3183),
.B(n_3111),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_SL g3299 ( 
.A(n_3192),
.B(n_3022),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_3143),
.B(n_3034),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_3134),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_SL g3302 ( 
.A(n_3198),
.B(n_3243),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_SL g3303 ( 
.A(n_3224),
.B(n_3193),
.Y(n_3303)
);

NOR2xp67_ASAP7_75t_L g3304 ( 
.A(n_3133),
.B(n_2885),
.Y(n_3304)
);

NAND2xp5_ASAP7_75t_L g3305 ( 
.A(n_3274),
.B(n_3036),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_3288),
.B(n_3038),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_3135),
.Y(n_3307)
);

BUFx5_ASAP7_75t_L g3308 ( 
.A(n_3144),
.Y(n_3308)
);

INVx2_ASAP7_75t_L g3309 ( 
.A(n_3159),
.Y(n_3309)
);

INVx4_ASAP7_75t_L g3310 ( 
.A(n_3133),
.Y(n_3310)
);

CKINVDCx5p33_ASAP7_75t_R g3311 ( 
.A(n_3174),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_3151),
.B(n_3039),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_SL g3313 ( 
.A(n_3155),
.B(n_3099),
.Y(n_3313)
);

INVx3_ASAP7_75t_L g3314 ( 
.A(n_3195),
.Y(n_3314)
);

BUFx6f_ASAP7_75t_L g3315 ( 
.A(n_3160),
.Y(n_3315)
);

NOR2xp33_ASAP7_75t_L g3316 ( 
.A(n_3199),
.B(n_2947),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_L g3317 ( 
.A(n_3152),
.B(n_3043),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_SL g3318 ( 
.A(n_3233),
.B(n_3045),
.Y(n_3318)
);

OAI22xp5_ASAP7_75t_L g3319 ( 
.A1(n_3280),
.A2(n_3117),
.B1(n_2903),
.B2(n_3023),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_SL g3320 ( 
.A(n_3264),
.B(n_3197),
.Y(n_3320)
);

INVx3_ASAP7_75t_L g3321 ( 
.A(n_3214),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_3156),
.B(n_3015),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_3158),
.B(n_3050),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_L g3324 ( 
.A(n_3161),
.B(n_3055),
.Y(n_3324)
);

NOR2xp33_ASAP7_75t_L g3325 ( 
.A(n_3189),
.B(n_2976),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3164),
.Y(n_3326)
);

O2A1O1Ixp33_ASAP7_75t_L g3327 ( 
.A1(n_3139),
.A2(n_2985),
.B(n_3019),
.C(n_3128),
.Y(n_3327)
);

INVx2_ASAP7_75t_L g3328 ( 
.A(n_3168),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_SL g3329 ( 
.A(n_3250),
.B(n_3041),
.Y(n_3329)
);

OAI221xp5_ASAP7_75t_L g3330 ( 
.A1(n_3212),
.A2(n_3000),
.B1(n_2965),
.B2(n_3078),
.C(n_3053),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_3165),
.B(n_3056),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_SL g3332 ( 
.A(n_3207),
.B(n_3010),
.Y(n_3332)
);

INVx1_ASAP7_75t_L g3333 ( 
.A(n_3176),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3180),
.Y(n_3334)
);

AND2x2_ASAP7_75t_L g3335 ( 
.A(n_3142),
.B(n_2974),
.Y(n_3335)
);

BUFx6f_ASAP7_75t_L g3336 ( 
.A(n_3160),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_SL g3337 ( 
.A(n_3282),
.B(n_3057),
.Y(n_3337)
);

AOI22xp5_ASAP7_75t_L g3338 ( 
.A1(n_3284),
.A2(n_3048),
.B1(n_2945),
.B2(n_3001),
.Y(n_3338)
);

NOR2xp33_ASAP7_75t_L g3339 ( 
.A(n_3252),
.B(n_3166),
.Y(n_3339)
);

INVx2_ASAP7_75t_L g3340 ( 
.A(n_3169),
.Y(n_3340)
);

INVxp67_ASAP7_75t_L g3341 ( 
.A(n_3175),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_3186),
.B(n_2986),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3196),
.Y(n_3343)
);

INVx3_ASAP7_75t_L g3344 ( 
.A(n_3217),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_L g3345 ( 
.A(n_3202),
.B(n_2987),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_L g3346 ( 
.A(n_3204),
.B(n_3210),
.Y(n_3346)
);

INVx2_ASAP7_75t_SL g3347 ( 
.A(n_3201),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_L g3348 ( 
.A(n_3213),
.B(n_2988),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_SL g3349 ( 
.A(n_3231),
.B(n_3065),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_3215),
.Y(n_3350)
);

BUFx6f_ASAP7_75t_L g3351 ( 
.A(n_3181),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3226),
.Y(n_3352)
);

INVx2_ASAP7_75t_SL g3353 ( 
.A(n_3201),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_3230),
.Y(n_3354)
);

INVx8_ASAP7_75t_L g3355 ( 
.A(n_3181),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3232),
.Y(n_3356)
);

AND2x4_ASAP7_75t_L g3357 ( 
.A(n_3255),
.B(n_3089),
.Y(n_3357)
);

AOI22xp5_ASAP7_75t_L g3358 ( 
.A1(n_3263),
.A2(n_3068),
.B1(n_3071),
.B2(n_3067),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_SL g3359 ( 
.A(n_3191),
.B(n_2993),
.Y(n_3359)
);

INVx2_ASAP7_75t_L g3360 ( 
.A(n_3182),
.Y(n_3360)
);

AOI22xp5_ASAP7_75t_L g3361 ( 
.A1(n_3229),
.A2(n_3131),
.B1(n_3187),
.B2(n_3177),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3236),
.Y(n_3362)
);

AND2x4_ASAP7_75t_L g3363 ( 
.A(n_3257),
.B(n_3100),
.Y(n_3363)
);

INVx2_ASAP7_75t_L g3364 ( 
.A(n_3185),
.Y(n_3364)
);

NOR2xp33_ASAP7_75t_L g3365 ( 
.A(n_3238),
.B(n_3076),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_3239),
.B(n_2994),
.Y(n_3366)
);

AOI22xp33_ASAP7_75t_L g3367 ( 
.A1(n_3286),
.A2(n_3081),
.B1(n_3083),
.B2(n_2995),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_L g3368 ( 
.A(n_3242),
.B(n_2982),
.Y(n_3368)
);

INVx4_ASAP7_75t_L g3369 ( 
.A(n_3184),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_L g3370 ( 
.A(n_3244),
.B(n_2992),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_3247),
.B(n_2997),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3253),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_3256),
.B(n_3127),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_3259),
.B(n_3137),
.Y(n_3374)
);

NOR2xp33_ASAP7_75t_SL g3375 ( 
.A(n_3251),
.B(n_2756),
.Y(n_3375)
);

OR2x6_ASAP7_75t_L g3376 ( 
.A(n_3157),
.B(n_2782),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_L g3377 ( 
.A(n_3141),
.B(n_3060),
.Y(n_3377)
);

BUFx6f_ASAP7_75t_L g3378 ( 
.A(n_3138),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_3287),
.B(n_3002),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_L g3380 ( 
.A(n_3290),
.B(n_3025),
.Y(n_3380)
);

AOI21xp5_ASAP7_75t_L g3381 ( 
.A1(n_3248),
.A2(n_3074),
.B(n_3072),
.Y(n_3381)
);

INVx2_ASAP7_75t_L g3382 ( 
.A(n_3200),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_SL g3383 ( 
.A(n_3245),
.B(n_3149),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_3271),
.B(n_3026),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_3273),
.B(n_3059),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_SL g3386 ( 
.A(n_3203),
.B(n_3206),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_3275),
.B(n_3059),
.Y(n_3387)
);

NOR2xp33_ASAP7_75t_L g3388 ( 
.A(n_3163),
.B(n_3052),
.Y(n_3388)
);

NAND3xp33_ASAP7_75t_SL g3389 ( 
.A(n_3172),
.B(n_3084),
.C(n_2657),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_3276),
.B(n_2967),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_3278),
.B(n_3066),
.Y(n_3391)
);

OAI22xp5_ASAP7_75t_L g3392 ( 
.A1(n_3208),
.A2(n_3104),
.B1(n_3080),
.B2(n_3075),
.Y(n_3392)
);

AOI22xp33_ASAP7_75t_L g3393 ( 
.A1(n_3216),
.A2(n_3005),
.B1(n_2948),
.B2(n_3106),
.Y(n_3393)
);

INVx2_ASAP7_75t_L g3394 ( 
.A(n_3220),
.Y(n_3394)
);

AND2x2_ASAP7_75t_L g3395 ( 
.A(n_3265),
.B(n_3105),
.Y(n_3395)
);

NOR2xp33_ASAP7_75t_L g3396 ( 
.A(n_3266),
.B(n_2981),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_3279),
.B(n_3108),
.Y(n_3397)
);

AOI22xp33_ASAP7_75t_L g3398 ( 
.A1(n_3223),
.A2(n_3240),
.B1(n_3272),
.B2(n_3227),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3283),
.B(n_3112),
.Y(n_3399)
);

NOR2xp67_ASAP7_75t_L g3400 ( 
.A(n_3262),
.B(n_3114),
.Y(n_3400)
);

AOI22xp33_ASAP7_75t_SL g3401 ( 
.A1(n_3173),
.A2(n_3258),
.B1(n_3170),
.B2(n_3179),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3268),
.B(n_3124),
.Y(n_3402)
);

INVx2_ASAP7_75t_SL g3403 ( 
.A(n_3171),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_3235),
.Y(n_3404)
);

AND2x2_ASAP7_75t_L g3405 ( 
.A(n_3269),
.B(n_3018),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_3270),
.B(n_3126),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_3267),
.B(n_2889),
.Y(n_3407)
);

BUFx2_ASAP7_75t_L g3408 ( 
.A(n_3190),
.Y(n_3408)
);

INVx2_ASAP7_75t_SL g3409 ( 
.A(n_3225),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_L g3410 ( 
.A(n_3218),
.B(n_2891),
.Y(n_3410)
);

AOI22xp33_ASAP7_75t_L g3411 ( 
.A1(n_3173),
.A2(n_3116),
.B1(n_3119),
.B2(n_3115),
.Y(n_3411)
);

NOR2xp33_ASAP7_75t_SL g3412 ( 
.A(n_3285),
.B(n_2820),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_SL g3413 ( 
.A(n_3225),
.B(n_3123),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_SL g3414 ( 
.A(n_3237),
.B(n_3125),
.Y(n_3414)
);

INVx2_ASAP7_75t_L g3415 ( 
.A(n_3228),
.Y(n_3415)
);

INVx2_ASAP7_75t_SL g3416 ( 
.A(n_3237),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_3254),
.B(n_2751),
.Y(n_3417)
);

AOI22xp5_ASAP7_75t_L g3418 ( 
.A1(n_3241),
.A2(n_3234),
.B1(n_3118),
.B2(n_3020),
.Y(n_3418)
);

AND2x2_ASAP7_75t_SL g3419 ( 
.A(n_3289),
.B(n_2685),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_3140),
.B(n_2773),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_3277),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_SL g3422 ( 
.A(n_3249),
.B(n_2685),
.Y(n_3422)
);

AOI22xp5_ASAP7_75t_L g3423 ( 
.A1(n_3170),
.A2(n_2808),
.B1(n_2777),
.B2(n_2629),
.Y(n_3423)
);

BUFx6f_ASAP7_75t_L g3424 ( 
.A(n_3260),
.Y(n_3424)
);

AOI22xp33_ASAP7_75t_L g3425 ( 
.A1(n_3205),
.A2(n_1336),
.B1(n_1431),
.B2(n_1428),
.Y(n_3425)
);

AOI22xp5_ASAP7_75t_L g3426 ( 
.A1(n_3339),
.A2(n_3281),
.B1(n_3162),
.B2(n_3209),
.Y(n_3426)
);

BUFx6f_ASAP7_75t_L g3427 ( 
.A(n_3315),
.Y(n_3427)
);

HB1xp67_ASAP7_75t_L g3428 ( 
.A(n_3296),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_3301),
.Y(n_3429)
);

INVx2_ASAP7_75t_L g3430 ( 
.A(n_3307),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_3326),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3333),
.Y(n_3432)
);

BUFx6f_ASAP7_75t_L g3433 ( 
.A(n_3315),
.Y(n_3433)
);

NAND2xp5_ASAP7_75t_L g3434 ( 
.A(n_3300),
.B(n_3147),
.Y(n_3434)
);

INVx3_ASAP7_75t_L g3435 ( 
.A(n_3310),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3292),
.B(n_3154),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_3302),
.B(n_3167),
.Y(n_3437)
);

HB1xp67_ASAP7_75t_L g3438 ( 
.A(n_3296),
.Y(n_3438)
);

INVx3_ASAP7_75t_SL g3439 ( 
.A(n_3311),
.Y(n_3439)
);

INVx1_ASAP7_75t_SL g3440 ( 
.A(n_3408),
.Y(n_3440)
);

INVx2_ASAP7_75t_L g3441 ( 
.A(n_3334),
.Y(n_3441)
);

HB1xp67_ASAP7_75t_L g3442 ( 
.A(n_3293),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_3343),
.Y(n_3443)
);

INVx2_ASAP7_75t_L g3444 ( 
.A(n_3350),
.Y(n_3444)
);

BUFx3_ASAP7_75t_L g3445 ( 
.A(n_3355),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3305),
.B(n_3249),
.Y(n_3446)
);

INVx2_ASAP7_75t_SL g3447 ( 
.A(n_3355),
.Y(n_3447)
);

INVxp67_ASAP7_75t_L g3448 ( 
.A(n_3378),
.Y(n_3448)
);

INVx2_ASAP7_75t_L g3449 ( 
.A(n_3352),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_3354),
.Y(n_3450)
);

INVx3_ASAP7_75t_L g3451 ( 
.A(n_3378),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3356),
.Y(n_3452)
);

INVx2_ASAP7_75t_L g3453 ( 
.A(n_3362),
.Y(n_3453)
);

AOI22xp5_ASAP7_75t_L g3454 ( 
.A1(n_3335),
.A2(n_2628),
.B1(n_3146),
.B2(n_3132),
.Y(n_3454)
);

INVx4_ASAP7_75t_L g3455 ( 
.A(n_3336),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3372),
.Y(n_3456)
);

AND2x6_ASAP7_75t_L g3457 ( 
.A(n_3336),
.B(n_3261),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3346),
.Y(n_3458)
);

INVx4_ASAP7_75t_L g3459 ( 
.A(n_3351),
.Y(n_3459)
);

INVx2_ASAP7_75t_L g3460 ( 
.A(n_3291),
.Y(n_3460)
);

INVx1_ASAP7_75t_SL g3461 ( 
.A(n_3351),
.Y(n_3461)
);

INVx3_ASAP7_75t_L g3462 ( 
.A(n_3424),
.Y(n_3462)
);

INVx2_ASAP7_75t_L g3463 ( 
.A(n_3295),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_SL g3464 ( 
.A(n_3341),
.B(n_3178),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_L g3465 ( 
.A(n_3306),
.B(n_3188),
.Y(n_3465)
);

AND2x4_ASAP7_75t_L g3466 ( 
.A(n_3369),
.B(n_3130),
.Y(n_3466)
);

INVx1_ASAP7_75t_L g3467 ( 
.A(n_3342),
.Y(n_3467)
);

OAI22xp5_ASAP7_75t_SL g3468 ( 
.A1(n_3401),
.A2(n_2729),
.B1(n_3194),
.B2(n_1410),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3345),
.Y(n_3469)
);

BUFx6f_ASAP7_75t_L g3470 ( 
.A(n_3424),
.Y(n_3470)
);

BUFx3_ASAP7_75t_L g3471 ( 
.A(n_3347),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3348),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3366),
.Y(n_3473)
);

INVx3_ASAP7_75t_L g3474 ( 
.A(n_3314),
.Y(n_3474)
);

INVx3_ASAP7_75t_L g3475 ( 
.A(n_3321),
.Y(n_3475)
);

INVx3_ASAP7_75t_SL g3476 ( 
.A(n_3376),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3312),
.Y(n_3477)
);

INVx2_ASAP7_75t_L g3478 ( 
.A(n_3309),
.Y(n_3478)
);

INVx4_ASAP7_75t_L g3479 ( 
.A(n_3344),
.Y(n_3479)
);

INVx4_ASAP7_75t_L g3480 ( 
.A(n_3297),
.Y(n_3480)
);

INVx2_ASAP7_75t_L g3481 ( 
.A(n_3328),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3317),
.Y(n_3482)
);

INVx2_ASAP7_75t_SL g3483 ( 
.A(n_3403),
.Y(n_3483)
);

BUFx6f_ASAP7_75t_L g3484 ( 
.A(n_3353),
.Y(n_3484)
);

BUFx3_ASAP7_75t_L g3485 ( 
.A(n_3409),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_L g3486 ( 
.A(n_3374),
.B(n_3246),
.Y(n_3486)
);

HB1xp67_ASAP7_75t_L g3487 ( 
.A(n_3416),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3322),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_SL g3489 ( 
.A(n_3320),
.B(n_2695),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_SL g3490 ( 
.A(n_3316),
.B(n_2695),
.Y(n_3490)
);

AOI22xp5_ASAP7_75t_L g3491 ( 
.A1(n_3298),
.A2(n_2646),
.B1(n_2640),
.B2(n_2706),
.Y(n_3491)
);

OR2x6_ASAP7_75t_L g3492 ( 
.A(n_3376),
.B(n_2877),
.Y(n_3492)
);

INVx2_ASAP7_75t_L g3493 ( 
.A(n_3340),
.Y(n_3493)
);

AND2x4_ASAP7_75t_L g3494 ( 
.A(n_3363),
.B(n_2923),
.Y(n_3494)
);

BUFx6f_ASAP7_75t_L g3495 ( 
.A(n_3419),
.Y(n_3495)
);

BUFx6f_ASAP7_75t_L g3496 ( 
.A(n_3357),
.Y(n_3496)
);

INVx5_ASAP7_75t_L g3497 ( 
.A(n_3405),
.Y(n_3497)
);

AOI22xp33_ASAP7_75t_L g3498 ( 
.A1(n_3330),
.A2(n_2961),
.B1(n_1550),
.B2(n_1554),
.Y(n_3498)
);

INVx4_ASAP7_75t_L g3499 ( 
.A(n_3415),
.Y(n_3499)
);

AOI22xp33_ASAP7_75t_L g3500 ( 
.A1(n_3294),
.A2(n_1559),
.B1(n_1565),
.B2(n_1549),
.Y(n_3500)
);

AND2x2_ASAP7_75t_L g3501 ( 
.A(n_3395),
.B(n_2856),
.Y(n_3501)
);

INVx3_ASAP7_75t_L g3502 ( 
.A(n_3421),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_3373),
.B(n_2707),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_SL g3504 ( 
.A(n_3325),
.B(n_2870),
.Y(n_3504)
);

HB1xp67_ASAP7_75t_L g3505 ( 
.A(n_3404),
.Y(n_3505)
);

INVx3_ASAP7_75t_L g3506 ( 
.A(n_3360),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3323),
.Y(n_3507)
);

INVx2_ASAP7_75t_SL g3508 ( 
.A(n_3407),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_L g3509 ( 
.A(n_3368),
.B(n_1694),
.Y(n_3509)
);

AND2x2_ASAP7_75t_L g3510 ( 
.A(n_3303),
.B(n_3090),
.Y(n_3510)
);

BUFx6f_ASAP7_75t_L g3511 ( 
.A(n_3422),
.Y(n_3511)
);

NOR2xp33_ASAP7_75t_L g3512 ( 
.A(n_3329),
.B(n_2841),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_L g3513 ( 
.A(n_3370),
.B(n_1695),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_3371),
.B(n_1697),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3324),
.Y(n_3515)
);

INVx3_ASAP7_75t_L g3516 ( 
.A(n_3364),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_L g3517 ( 
.A(n_3377),
.B(n_1709),
.Y(n_3517)
);

INVx2_ASAP7_75t_SL g3518 ( 
.A(n_3313),
.Y(n_3518)
);

AND2x2_ASAP7_75t_SL g3519 ( 
.A(n_3412),
.B(n_1428),
.Y(n_3519)
);

AO22x1_ASAP7_75t_L g3520 ( 
.A1(n_3365),
.A2(n_1415),
.B1(n_1419),
.B2(n_1407),
.Y(n_3520)
);

INVx3_ASAP7_75t_L g3521 ( 
.A(n_3382),
.Y(n_3521)
);

OAI21xp5_ASAP7_75t_L g3522 ( 
.A1(n_3299),
.A2(n_3003),
.B(n_2680),
.Y(n_3522)
);

INVx2_ASAP7_75t_L g3523 ( 
.A(n_3394),
.Y(n_3523)
);

BUFx3_ASAP7_75t_L g3524 ( 
.A(n_3388),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3331),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_3384),
.Y(n_3526)
);

BUFx6f_ASAP7_75t_L g3527 ( 
.A(n_3410),
.Y(n_3527)
);

INVx3_ASAP7_75t_L g3528 ( 
.A(n_3308),
.Y(n_3528)
);

INVx3_ASAP7_75t_L g3529 ( 
.A(n_3308),
.Y(n_3529)
);

BUFx2_ASAP7_75t_L g3530 ( 
.A(n_3420),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3380),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_SL g3532 ( 
.A(n_3338),
.B(n_1713),
.Y(n_3532)
);

OAI22xp5_ASAP7_75t_L g3533 ( 
.A1(n_3426),
.A2(n_3411),
.B1(n_3361),
.B2(n_3358),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_3430),
.Y(n_3534)
);

A2O1A1Ixp33_ASAP7_75t_L g3535 ( 
.A1(n_3512),
.A2(n_3327),
.B(n_3383),
.C(n_3381),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_SL g3536 ( 
.A(n_3527),
.B(n_3308),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3441),
.Y(n_3537)
);

NOR3xp33_ASAP7_75t_SL g3538 ( 
.A(n_3504),
.B(n_3389),
.C(n_3332),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3458),
.B(n_3349),
.Y(n_3539)
);

AOI21xp5_ASAP7_75t_L g3540 ( 
.A1(n_3522),
.A2(n_3319),
.B(n_3392),
.Y(n_3540)
);

A2O1A1Ixp33_ASAP7_75t_L g3541 ( 
.A1(n_3498),
.A2(n_3396),
.B(n_3318),
.C(n_3418),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_3444),
.Y(n_3542)
);

OA22x2_ASAP7_75t_L g3543 ( 
.A1(n_3454),
.A2(n_3417),
.B1(n_3414),
.B2(n_3413),
.Y(n_3543)
);

AND2x2_ASAP7_75t_L g3544 ( 
.A(n_3442),
.B(n_3530),
.Y(n_3544)
);

AOI21xp5_ASAP7_75t_L g3545 ( 
.A1(n_3532),
.A2(n_3390),
.B(n_3391),
.Y(n_3545)
);

O2A1O1Ixp5_ASAP7_75t_SL g3546 ( 
.A1(n_3489),
.A2(n_3359),
.B(n_3386),
.C(n_3337),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_3477),
.B(n_3397),
.Y(n_3547)
);

INVx2_ASAP7_75t_L g3548 ( 
.A(n_3449),
.Y(n_3548)
);

A2O1A1Ixp33_ASAP7_75t_L g3549 ( 
.A1(n_3482),
.A2(n_3399),
.B(n_3379),
.C(n_3423),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3453),
.Y(n_3550)
);

INVx2_ASAP7_75t_SL g3551 ( 
.A(n_3470),
.Y(n_3551)
);

AOI21xp5_ASAP7_75t_L g3552 ( 
.A1(n_3528),
.A2(n_3393),
.B(n_3387),
.Y(n_3552)
);

A2O1A1Ixp33_ASAP7_75t_L g3553 ( 
.A1(n_3488),
.A2(n_3385),
.B(n_3400),
.C(n_3367),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_3429),
.Y(n_3554)
);

BUFx6f_ASAP7_75t_L g3555 ( 
.A(n_3470),
.Y(n_3555)
);

BUFx2_ASAP7_75t_L g3556 ( 
.A(n_3495),
.Y(n_3556)
);

O2A1O1Ixp33_ASAP7_75t_SL g3557 ( 
.A1(n_3464),
.A2(n_3406),
.B(n_3402),
.C(n_1578),
.Y(n_3557)
);

NOR2xp33_ASAP7_75t_L g3558 ( 
.A(n_3524),
.B(n_3375),
.Y(n_3558)
);

AND2x4_ASAP7_75t_L g3559 ( 
.A(n_3451),
.B(n_3304),
.Y(n_3559)
);

O2A1O1Ixp33_ASAP7_75t_L g3560 ( 
.A1(n_3490),
.A2(n_1579),
.B(n_1591),
.C(n_1569),
.Y(n_3560)
);

OAI21xp33_ASAP7_75t_L g3561 ( 
.A1(n_3519),
.A2(n_3425),
.B(n_3398),
.Y(n_3561)
);

INVx2_ASAP7_75t_L g3562 ( 
.A(n_3460),
.Y(n_3562)
);

NAND2x1p5_ASAP7_75t_L g3563 ( 
.A(n_3479),
.B(n_3308),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_3463),
.Y(n_3564)
);

NOR2xp33_ASAP7_75t_R g3565 ( 
.A(n_3462),
.B(n_1715),
.Y(n_3565)
);

BUFx6f_ASAP7_75t_L g3566 ( 
.A(n_3427),
.Y(n_3566)
);

OAI22xp5_ASAP7_75t_L g3567 ( 
.A1(n_3486),
.A2(n_1446),
.B1(n_1447),
.B2(n_1421),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_SL g3568 ( 
.A(n_3527),
.B(n_1723),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_L g3569 ( 
.A(n_3507),
.B(n_1449),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_SL g3570 ( 
.A(n_3518),
.B(n_1727),
.Y(n_3570)
);

INVx2_ASAP7_75t_SL g3571 ( 
.A(n_3427),
.Y(n_3571)
);

A2O1A1Ixp33_ASAP7_75t_L g3572 ( 
.A1(n_3515),
.A2(n_1601),
.B(n_1602),
.C(n_1600),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3525),
.B(n_1452),
.Y(n_3573)
);

AOI21xp5_ASAP7_75t_L g3574 ( 
.A1(n_3529),
.A2(n_2691),
.B(n_2632),
.Y(n_3574)
);

AOI21xp5_ASAP7_75t_L g3575 ( 
.A1(n_3517),
.A2(n_1441),
.B(n_1431),
.Y(n_3575)
);

AOI21xp5_ASAP7_75t_L g3576 ( 
.A1(n_3467),
.A2(n_1441),
.B(n_1431),
.Y(n_3576)
);

BUFx12f_ASAP7_75t_L g3577 ( 
.A(n_3480),
.Y(n_3577)
);

NOR2xp33_ASAP7_75t_SL g3578 ( 
.A(n_3439),
.B(n_1733),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_L g3579 ( 
.A(n_3469),
.B(n_1456),
.Y(n_3579)
);

OAI221xp5_ASAP7_75t_L g3580 ( 
.A1(n_3500),
.A2(n_1610),
.B1(n_1616),
.B2(n_1606),
.C(n_1605),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3472),
.B(n_1457),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_SL g3582 ( 
.A(n_3465),
.B(n_3473),
.Y(n_3582)
);

AOI222xp33_ASAP7_75t_L g3583 ( 
.A1(n_3520),
.A2(n_1463),
.B1(n_1459),
.B2(n_1471),
.C1(n_1464),
.C2(n_1462),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_L g3584 ( 
.A(n_3526),
.B(n_1472),
.Y(n_3584)
);

A2O1A1Ixp33_ASAP7_75t_L g3585 ( 
.A1(n_3437),
.A2(n_1624),
.B(n_1642),
.C(n_1622),
.Y(n_3585)
);

AOI21xp5_ASAP7_75t_L g3586 ( 
.A1(n_3531),
.A2(n_1488),
.B(n_1441),
.Y(n_3586)
);

INVx4_ASAP7_75t_L g3587 ( 
.A(n_3457),
.Y(n_3587)
);

INVx2_ASAP7_75t_L g3588 ( 
.A(n_3478),
.Y(n_3588)
);

AOI21xp5_ASAP7_75t_L g3589 ( 
.A1(n_3509),
.A2(n_1571),
.B(n_1488),
.Y(n_3589)
);

AND2x2_ASAP7_75t_L g3590 ( 
.A(n_3508),
.B(n_1645),
.Y(n_3590)
);

BUFx12f_ASAP7_75t_L g3591 ( 
.A(n_3466),
.Y(n_3591)
);

AND2x4_ASAP7_75t_L g3592 ( 
.A(n_3448),
.B(n_1648),
.Y(n_3592)
);

OAI21xp5_ASAP7_75t_L g3593 ( 
.A1(n_3513),
.A2(n_1657),
.B(n_1654),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_L g3594 ( 
.A(n_3434),
.B(n_1473),
.Y(n_3594)
);

AOI21x1_ASAP7_75t_L g3595 ( 
.A1(n_3510),
.A2(n_1672),
.B(n_1666),
.Y(n_3595)
);

INVx1_ASAP7_75t_L g3596 ( 
.A(n_3431),
.Y(n_3596)
);

AND2x2_ASAP7_75t_L g3597 ( 
.A(n_3501),
.B(n_1675),
.Y(n_3597)
);

AOI22xp33_ASAP7_75t_L g3598 ( 
.A1(n_3495),
.A2(n_1687),
.B1(n_1701),
.B2(n_1682),
.Y(n_3598)
);

OAI22xp5_ASAP7_75t_L g3599 ( 
.A1(n_3436),
.A2(n_1477),
.B1(n_1478),
.B2(n_1475),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_SL g3600 ( 
.A(n_3497),
.B(n_1739),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3432),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3443),
.Y(n_3602)
);

A2O1A1Ixp33_ASAP7_75t_L g3603 ( 
.A1(n_3514),
.A2(n_1708),
.B(n_1710),
.C(n_1705),
.Y(n_3603)
);

BUFx8_ASAP7_75t_L g3604 ( 
.A(n_3457),
.Y(n_3604)
);

NOR2xp33_ASAP7_75t_L g3605 ( 
.A(n_3440),
.B(n_1743),
.Y(n_3605)
);

AOI21xp5_ASAP7_75t_L g3606 ( 
.A1(n_3503),
.A2(n_1571),
.B(n_1488),
.Y(n_3606)
);

CKINVDCx8_ASAP7_75t_R g3607 ( 
.A(n_3433),
.Y(n_3607)
);

INVx1_ASAP7_75t_L g3608 ( 
.A(n_3450),
.Y(n_3608)
);

AOI21xp5_ASAP7_75t_L g3609 ( 
.A1(n_3446),
.A2(n_1901),
.B(n_1571),
.Y(n_3609)
);

OR2x6_ASAP7_75t_L g3610 ( 
.A(n_3445),
.B(n_1901),
.Y(n_3610)
);

NOR2xp33_ASAP7_75t_L g3611 ( 
.A(n_3499),
.B(n_1745),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_L g3612 ( 
.A(n_3505),
.B(n_1479),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3452),
.Y(n_3613)
);

INVx2_ASAP7_75t_L g3614 ( 
.A(n_3481),
.Y(n_3614)
);

NAND2x1p5_ASAP7_75t_L g3615 ( 
.A(n_3455),
.B(n_1901),
.Y(n_3615)
);

AOI21xp5_ASAP7_75t_L g3616 ( 
.A1(n_3492),
.A2(n_1751),
.B(n_1748),
.Y(n_3616)
);

INVx2_ASAP7_75t_L g3617 ( 
.A(n_3493),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_SL g3618 ( 
.A(n_3497),
.B(n_3496),
.Y(n_3618)
);

BUFx6f_ASAP7_75t_L g3619 ( 
.A(n_3433),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3456),
.Y(n_3620)
);

AOI21xp5_ASAP7_75t_L g3621 ( 
.A1(n_3523),
.A2(n_1759),
.B(n_1757),
.Y(n_3621)
);

OAI22xp5_ASAP7_75t_L g3622 ( 
.A1(n_3502),
.A2(n_1489),
.B1(n_1490),
.B2(n_1486),
.Y(n_3622)
);

AO21x1_ASAP7_75t_L g3623 ( 
.A1(n_3491),
.A2(n_1716),
.B(n_1714),
.Y(n_3623)
);

OAI21xp33_ASAP7_75t_SL g3624 ( 
.A1(n_3521),
.A2(n_1720),
.B(n_1717),
.Y(n_3624)
);

INVxp67_ASAP7_75t_L g3625 ( 
.A(n_3487),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_L g3626 ( 
.A(n_3506),
.B(n_1492),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3516),
.Y(n_3627)
);

AO32x2_ASAP7_75t_L g3628 ( 
.A1(n_3468),
.A2(n_2),
.A3(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_3628)
);

INVx3_ASAP7_75t_L g3629 ( 
.A(n_3484),
.Y(n_3629)
);

NOR2xp33_ASAP7_75t_L g3630 ( 
.A(n_3496),
.B(n_1762),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3511),
.Y(n_3631)
);

NOR2xp33_ASAP7_75t_R g3632 ( 
.A(n_3447),
.B(n_1772),
.Y(n_3632)
);

INVx6_ASAP7_75t_L g3633 ( 
.A(n_3459),
.Y(n_3633)
);

AOI21xp5_ASAP7_75t_L g3634 ( 
.A1(n_3474),
.A2(n_1787),
.B(n_1782),
.Y(n_3634)
);

NAND2x1p5_ASAP7_75t_L g3635 ( 
.A(n_3485),
.B(n_1721),
.Y(n_3635)
);

NAND3xp33_ASAP7_75t_L g3636 ( 
.A(n_3428),
.B(n_1494),
.C(n_1493),
.Y(n_3636)
);

CKINVDCx5p33_ASAP7_75t_R g3637 ( 
.A(n_3476),
.Y(n_3637)
);

NOR3xp33_ASAP7_75t_SL g3638 ( 
.A(n_3438),
.B(n_1499),
.C(n_1498),
.Y(n_3638)
);

NOR2xp33_ASAP7_75t_R g3639 ( 
.A(n_3435),
.B(n_1790),
.Y(n_3639)
);

A2O1A1Ixp33_ASAP7_75t_L g3640 ( 
.A1(n_3511),
.A2(n_1730),
.B(n_1731),
.C(n_1729),
.Y(n_3640)
);

AOI21xp5_ASAP7_75t_L g3641 ( 
.A1(n_3475),
.A2(n_1800),
.B(n_1797),
.Y(n_3641)
);

AOI21xp5_ASAP7_75t_L g3642 ( 
.A1(n_3483),
.A2(n_1805),
.B(n_1802),
.Y(n_3642)
);

OR2x6_ASAP7_75t_L g3643 ( 
.A(n_3484),
.B(n_3494),
.Y(n_3643)
);

INVx2_ASAP7_75t_L g3644 ( 
.A(n_3471),
.Y(n_3644)
);

OAI21xp5_ASAP7_75t_L g3645 ( 
.A1(n_3461),
.A2(n_1746),
.B(n_1740),
.Y(n_3645)
);

BUFx12f_ASAP7_75t_L g3646 ( 
.A(n_3604),
.Y(n_3646)
);

INVx1_ASAP7_75t_L g3647 ( 
.A(n_3554),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_L g3648 ( 
.A(n_3582),
.B(n_1502),
.Y(n_3648)
);

O2A1O1Ixp33_ASAP7_75t_L g3649 ( 
.A1(n_3593),
.A2(n_1767),
.B(n_1769),
.C(n_1756),
.Y(n_3649)
);

BUFx12f_ASAP7_75t_L g3650 ( 
.A(n_3637),
.Y(n_3650)
);

BUFx6f_ASAP7_75t_L g3651 ( 
.A(n_3555),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_3596),
.Y(n_3652)
);

AOI22xp5_ASAP7_75t_L g3653 ( 
.A1(n_3533),
.A2(n_1515),
.B1(n_1516),
.B2(n_1513),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_3601),
.Y(n_3654)
);

AOI22xp33_ASAP7_75t_SL g3655 ( 
.A1(n_3645),
.A2(n_3543),
.B1(n_3558),
.B2(n_3540),
.Y(n_3655)
);

BUFx3_ASAP7_75t_L g3656 ( 
.A(n_3607),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3602),
.Y(n_3657)
);

BUFx6f_ASAP7_75t_L g3658 ( 
.A(n_3555),
.Y(n_3658)
);

CKINVDCx5p33_ASAP7_75t_R g3659 ( 
.A(n_3577),
.Y(n_3659)
);

INVx2_ASAP7_75t_L g3660 ( 
.A(n_3534),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_3547),
.B(n_3544),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3608),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3539),
.B(n_1518),
.Y(n_3663)
);

INVx2_ASAP7_75t_L g3664 ( 
.A(n_3542),
.Y(n_3664)
);

OR2x6_ASAP7_75t_SL g3665 ( 
.A(n_3636),
.B(n_1520),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_L g3666 ( 
.A(n_3549),
.B(n_3548),
.Y(n_3666)
);

INVx2_ASAP7_75t_L g3667 ( 
.A(n_3562),
.Y(n_3667)
);

BUFx6f_ASAP7_75t_L g3668 ( 
.A(n_3566),
.Y(n_3668)
);

INVx2_ASAP7_75t_SL g3669 ( 
.A(n_3633),
.Y(n_3669)
);

NOR2xp33_ASAP7_75t_L g3670 ( 
.A(n_3556),
.B(n_1827),
.Y(n_3670)
);

BUFx3_ASAP7_75t_L g3671 ( 
.A(n_3566),
.Y(n_3671)
);

OR2x6_ASAP7_75t_L g3672 ( 
.A(n_3618),
.B(n_1774),
.Y(n_3672)
);

AOI22xp33_ASAP7_75t_L g3673 ( 
.A1(n_3623),
.A2(n_1791),
.B1(n_1794),
.B2(n_1776),
.Y(n_3673)
);

INVx4_ASAP7_75t_L g3674 ( 
.A(n_3587),
.Y(n_3674)
);

AOI22xp33_ASAP7_75t_L g3675 ( 
.A1(n_3561),
.A2(n_1809),
.B1(n_1810),
.B2(n_1796),
.Y(n_3675)
);

NAND2x1p5_ASAP7_75t_L g3676 ( 
.A(n_3536),
.B(n_1814),
.Y(n_3676)
);

AOI22xp5_ASAP7_75t_L g3677 ( 
.A1(n_3538),
.A2(n_1529),
.B1(n_1532),
.B2(n_1525),
.Y(n_3677)
);

INVx2_ASAP7_75t_L g3678 ( 
.A(n_3564),
.Y(n_3678)
);

AND2x4_ASAP7_75t_L g3679 ( 
.A(n_3644),
.B(n_961),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3613),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_3620),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_3537),
.B(n_1534),
.Y(n_3682)
);

CKINVDCx5p33_ASAP7_75t_R g3683 ( 
.A(n_3591),
.Y(n_3683)
);

OAI22xp33_ASAP7_75t_L g3684 ( 
.A1(n_3610),
.A2(n_1537),
.B1(n_1541),
.B2(n_1535),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3550),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_L g3686 ( 
.A(n_3541),
.B(n_1551),
.Y(n_3686)
);

BUFx12f_ASAP7_75t_L g3687 ( 
.A(n_3619),
.Y(n_3687)
);

INVx2_ASAP7_75t_SL g3688 ( 
.A(n_3633),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_L g3689 ( 
.A(n_3588),
.B(n_1558),
.Y(n_3689)
);

BUFx6f_ASAP7_75t_L g3690 ( 
.A(n_3619),
.Y(n_3690)
);

NOR2xp33_ASAP7_75t_L g3691 ( 
.A(n_3605),
.B(n_1833),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3614),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_L g3693 ( 
.A(n_3617),
.B(n_1560),
.Y(n_3693)
);

CKINVDCx5p33_ASAP7_75t_R g3694 ( 
.A(n_3643),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_3597),
.B(n_1562),
.Y(n_3695)
);

NOR2x1_ASAP7_75t_SL g3696 ( 
.A(n_3595),
.B(n_1815),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_L g3697 ( 
.A(n_3535),
.B(n_1568),
.Y(n_3697)
);

AND2x2_ASAP7_75t_SL g3698 ( 
.A(n_3578),
.B(n_1816),
.Y(n_3698)
);

INVx4_ASAP7_75t_L g3699 ( 
.A(n_3629),
.Y(n_3699)
);

INVx1_ASAP7_75t_SL g3700 ( 
.A(n_3565),
.Y(n_3700)
);

INVx4_ASAP7_75t_L g3701 ( 
.A(n_3643),
.Y(n_3701)
);

CKINVDCx5p33_ASAP7_75t_R g3702 ( 
.A(n_3632),
.Y(n_3702)
);

BUFx2_ASAP7_75t_L g3703 ( 
.A(n_3631),
.Y(n_3703)
);

INVx2_ASAP7_75t_L g3704 ( 
.A(n_3627),
.Y(n_3704)
);

NAND2xp5_ASAP7_75t_SL g3705 ( 
.A(n_3553),
.B(n_1845),
.Y(n_3705)
);

HB1xp67_ASAP7_75t_L g3706 ( 
.A(n_3625),
.Y(n_3706)
);

OR2x2_ASAP7_75t_L g3707 ( 
.A(n_3612),
.B(n_3594),
.Y(n_3707)
);

A2O1A1Ixp33_ASAP7_75t_L g3708 ( 
.A1(n_3603),
.A2(n_3545),
.B(n_3589),
.C(n_3575),
.Y(n_3708)
);

BUFx6f_ASAP7_75t_L g3709 ( 
.A(n_3551),
.Y(n_3709)
);

INVx2_ASAP7_75t_L g3710 ( 
.A(n_3590),
.Y(n_3710)
);

NOR2x1_ASAP7_75t_L g3711 ( 
.A(n_3600),
.B(n_3568),
.Y(n_3711)
);

HB1xp67_ASAP7_75t_L g3712 ( 
.A(n_3563),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3560),
.Y(n_3713)
);

AOI21xp5_ASAP7_75t_L g3714 ( 
.A1(n_3552),
.A2(n_1860),
.B(n_1858),
.Y(n_3714)
);

BUFx6f_ASAP7_75t_SL g3715 ( 
.A(n_3559),
.Y(n_3715)
);

BUFx2_ASAP7_75t_R g3716 ( 
.A(n_3570),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3628),
.Y(n_3717)
);

BUFx6f_ASAP7_75t_L g3718 ( 
.A(n_3571),
.Y(n_3718)
);

OAI22xp5_ASAP7_75t_SL g3719 ( 
.A1(n_3598),
.A2(n_3610),
.B1(n_3635),
.B2(n_3580),
.Y(n_3719)
);

INVx3_ASAP7_75t_L g3720 ( 
.A(n_3592),
.Y(n_3720)
);

XOR2xp5_ASAP7_75t_L g3721 ( 
.A(n_3599),
.B(n_962),
.Y(n_3721)
);

OAI21xp5_ASAP7_75t_L g3722 ( 
.A1(n_3546),
.A2(n_1830),
.B(n_1826),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_L g3723 ( 
.A(n_3569),
.B(n_1572),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3628),
.Y(n_3724)
);

HB1xp67_ASAP7_75t_L g3725 ( 
.A(n_3626),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3585),
.Y(n_3726)
);

INVx2_ASAP7_75t_L g3727 ( 
.A(n_3573),
.Y(n_3727)
);

INVx1_ASAP7_75t_L g3728 ( 
.A(n_3572),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_3579),
.B(n_1574),
.Y(n_3729)
);

CKINVDCx5p33_ASAP7_75t_R g3730 ( 
.A(n_3639),
.Y(n_3730)
);

AOI22xp33_ASAP7_75t_L g3731 ( 
.A1(n_3583),
.A2(n_1834),
.B1(n_1841),
.B2(n_1831),
.Y(n_3731)
);

BUFx6f_ASAP7_75t_L g3732 ( 
.A(n_3630),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_3581),
.B(n_1576),
.Y(n_3733)
);

INVx3_ASAP7_75t_L g3734 ( 
.A(n_3615),
.Y(n_3734)
);

NAND2x1p5_ASAP7_75t_L g3735 ( 
.A(n_3611),
.B(n_1850),
.Y(n_3735)
);

INVx2_ASAP7_75t_SL g3736 ( 
.A(n_3584),
.Y(n_3736)
);

INVx3_ASAP7_75t_L g3737 ( 
.A(n_3638),
.Y(n_3737)
);

INVx2_ASAP7_75t_L g3738 ( 
.A(n_3567),
.Y(n_3738)
);

AND2x2_ASAP7_75t_L g3739 ( 
.A(n_3640),
.B(n_1861),
.Y(n_3739)
);

INVx2_ASAP7_75t_L g3740 ( 
.A(n_3622),
.Y(n_3740)
);

AOI22xp5_ASAP7_75t_L g3741 ( 
.A1(n_3624),
.A2(n_1585),
.B1(n_1586),
.B2(n_1584),
.Y(n_3741)
);

INVx4_ASAP7_75t_L g3742 ( 
.A(n_3557),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3616),
.B(n_3609),
.Y(n_3743)
);

AOI21xp5_ASAP7_75t_L g3744 ( 
.A1(n_3708),
.A2(n_3576),
.B(n_3586),
.Y(n_3744)
);

OAI21x1_ASAP7_75t_L g3745 ( 
.A1(n_3743),
.A2(n_3606),
.B(n_3574),
.Y(n_3745)
);

A2O1A1Ixp33_ASAP7_75t_L g3746 ( 
.A1(n_3655),
.A2(n_3642),
.B(n_3621),
.C(n_3641),
.Y(n_3746)
);

OAI21xp5_ASAP7_75t_L g3747 ( 
.A1(n_3686),
.A2(n_3634),
.B(n_1881),
.Y(n_3747)
);

AND2x4_ASAP7_75t_L g3748 ( 
.A(n_3703),
.B(n_966),
.Y(n_3748)
);

AND2x2_ASAP7_75t_L g3749 ( 
.A(n_3661),
.B(n_3647),
.Y(n_3749)
);

INVx2_ASAP7_75t_SL g3750 ( 
.A(n_3651),
.Y(n_3750)
);

AOI22xp33_ASAP7_75t_L g3751 ( 
.A1(n_3698),
.A2(n_1887),
.B1(n_1894),
.B2(n_1867),
.Y(n_3751)
);

AOI21xp5_ASAP7_75t_L g3752 ( 
.A1(n_3705),
.A2(n_1873),
.B(n_1869),
.Y(n_3752)
);

BUFx2_ASAP7_75t_L g3753 ( 
.A(n_3701),
.Y(n_3753)
);

A2O1A1Ixp33_ASAP7_75t_L g3754 ( 
.A1(n_3653),
.A2(n_1902),
.B(n_1908),
.C(n_1900),
.Y(n_3754)
);

A2O1A1Ixp33_ASAP7_75t_L g3755 ( 
.A1(n_3691),
.A2(n_1923),
.B(n_1924),
.C(n_1916),
.Y(n_3755)
);

INVx3_ASAP7_75t_L g3756 ( 
.A(n_3651),
.Y(n_3756)
);

BUFx2_ASAP7_75t_L g3757 ( 
.A(n_3706),
.Y(n_3757)
);

INVx5_ASAP7_75t_L g3758 ( 
.A(n_3646),
.Y(n_3758)
);

AOI221x1_ASAP7_75t_L g3759 ( 
.A1(n_3717),
.A2(n_1931),
.B1(n_1939),
.B2(n_1936),
.C(n_1927),
.Y(n_3759)
);

OAI21x1_ASAP7_75t_SL g3760 ( 
.A1(n_3696),
.A2(n_1995),
.B(n_1930),
.Y(n_3760)
);

O2A1O1Ixp33_ASAP7_75t_L g3761 ( 
.A1(n_3697),
.A2(n_1959),
.B(n_1964),
.C(n_1942),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3652),
.Y(n_3762)
);

INVx2_ASAP7_75t_L g3763 ( 
.A(n_3685),
.Y(n_3763)
);

BUFx12f_ASAP7_75t_L g3764 ( 
.A(n_3659),
.Y(n_3764)
);

INVx2_ASAP7_75t_L g3765 ( 
.A(n_3654),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_3657),
.Y(n_3766)
);

AND2x2_ASAP7_75t_L g3767 ( 
.A(n_3662),
.B(n_1970),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3680),
.Y(n_3768)
);

BUFx2_ASAP7_75t_L g3769 ( 
.A(n_3694),
.Y(n_3769)
);

OAI21xp5_ASAP7_75t_L g3770 ( 
.A1(n_3714),
.A2(n_1983),
.B(n_1972),
.Y(n_3770)
);

AOI22xp5_ASAP7_75t_L g3771 ( 
.A1(n_3719),
.A2(n_1588),
.B1(n_1592),
.B2(n_1587),
.Y(n_3771)
);

INVx2_ASAP7_75t_L g3772 ( 
.A(n_3681),
.Y(n_3772)
);

NAND3xp33_ASAP7_75t_SL g3773 ( 
.A(n_3735),
.B(n_1597),
.C(n_1595),
.Y(n_3773)
);

OAI221xp5_ASAP7_75t_L g3774 ( 
.A1(n_3731),
.A2(n_1998),
.B1(n_2005),
.B2(n_1994),
.C(n_1989),
.Y(n_3774)
);

OAI22xp5_ASAP7_75t_L g3775 ( 
.A1(n_3736),
.A2(n_3675),
.B1(n_3707),
.B2(n_3721),
.Y(n_3775)
);

CKINVDCx20_ASAP7_75t_R g3776 ( 
.A(n_3730),
.Y(n_3776)
);

AOI21xp5_ASAP7_75t_L g3777 ( 
.A1(n_3666),
.A2(n_1886),
.B(n_1875),
.Y(n_3777)
);

OAI21xp5_ASAP7_75t_L g3778 ( 
.A1(n_3649),
.A2(n_2014),
.B(n_2013),
.Y(n_3778)
);

OAI21x1_ASAP7_75t_L g3779 ( 
.A1(n_3722),
.A2(n_2031),
.B(n_2017),
.Y(n_3779)
);

OAI21x1_ASAP7_75t_L g3780 ( 
.A1(n_3692),
.A2(n_2046),
.B(n_2037),
.Y(n_3780)
);

INVx2_ASAP7_75t_SL g3781 ( 
.A(n_3658),
.Y(n_3781)
);

AND2x2_ASAP7_75t_L g3782 ( 
.A(n_3710),
.B(n_2000),
.Y(n_3782)
);

BUFx3_ASAP7_75t_L g3783 ( 
.A(n_3671),
.Y(n_3783)
);

OAI22xp5_ASAP7_75t_L g3784 ( 
.A1(n_3672),
.A2(n_1599),
.B1(n_1611),
.B2(n_1598),
.Y(n_3784)
);

NOR2xp33_ASAP7_75t_L g3785 ( 
.A(n_3732),
.B(n_1613),
.Y(n_3785)
);

NAND2xp33_ASAP7_75t_SL g3786 ( 
.A(n_3702),
.B(n_3732),
.Y(n_3786)
);

OR2x6_ASAP7_75t_L g3787 ( 
.A(n_3674),
.B(n_2012),
.Y(n_3787)
);

A2O1A1Ixp33_ASAP7_75t_L g3788 ( 
.A1(n_3738),
.A2(n_2021),
.B(n_2018),
.C(n_1617),
.Y(n_3788)
);

A2O1A1Ixp33_ASAP7_75t_L g3789 ( 
.A1(n_3728),
.A2(n_1621),
.B(n_1623),
.C(n_1614),
.Y(n_3789)
);

OAI21x1_ASAP7_75t_L g3790 ( 
.A1(n_3660),
.A2(n_968),
.B(n_967),
.Y(n_3790)
);

NOR2xp33_ASAP7_75t_L g3791 ( 
.A(n_3727),
.B(n_3716),
.Y(n_3791)
);

A2O1A1Ixp33_ASAP7_75t_L g3792 ( 
.A1(n_3726),
.A2(n_1627),
.B(n_1628),
.C(n_1626),
.Y(n_3792)
);

OAI22x1_ASAP7_75t_SL g3793 ( 
.A1(n_3683),
.A2(n_1638),
.B1(n_1641),
.B2(n_1634),
.Y(n_3793)
);

NOR2x1_ASAP7_75t_SL g3794 ( 
.A(n_3724),
.B(n_969),
.Y(n_3794)
);

NOR2xp33_ASAP7_75t_L g3795 ( 
.A(n_3700),
.B(n_1646),
.Y(n_3795)
);

A2O1A1Ixp33_ASAP7_75t_L g3796 ( 
.A1(n_3711),
.A2(n_1655),
.B(n_1662),
.C(n_1647),
.Y(n_3796)
);

INVx1_ASAP7_75t_SL g3797 ( 
.A(n_3656),
.Y(n_3797)
);

OAI21x1_ASAP7_75t_L g3798 ( 
.A1(n_3664),
.A2(n_980),
.B(n_970),
.Y(n_3798)
);

A2O1A1Ixp33_ASAP7_75t_L g3799 ( 
.A1(n_3713),
.A2(n_1669),
.B(n_1670),
.C(n_1667),
.Y(n_3799)
);

BUFx12f_ASAP7_75t_L g3800 ( 
.A(n_3650),
.Y(n_3800)
);

INVx1_ASAP7_75t_L g3801 ( 
.A(n_3704),
.Y(n_3801)
);

AOI21xp5_ASAP7_75t_L g3802 ( 
.A1(n_3725),
.A2(n_3673),
.B(n_3648),
.Y(n_3802)
);

NAND2xp5_ASAP7_75t_L g3803 ( 
.A(n_3667),
.B(n_1671),
.Y(n_3803)
);

BUFx6f_ASAP7_75t_L g3804 ( 
.A(n_3658),
.Y(n_3804)
);

NAND2xp5_ASAP7_75t_L g3805 ( 
.A(n_3678),
.B(n_3663),
.Y(n_3805)
);

O2A1O1Ixp33_ASAP7_75t_L g3806 ( 
.A1(n_3684),
.A2(n_1676),
.B(n_1680),
.C(n_1674),
.Y(n_3806)
);

INVx1_ASAP7_75t_SL g3807 ( 
.A(n_3709),
.Y(n_3807)
);

AO32x2_ASAP7_75t_L g3808 ( 
.A1(n_3742),
.A2(n_6),
.A3(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_3808)
);

O2A1O1Ixp5_ASAP7_75t_L g3809 ( 
.A1(n_3740),
.A2(n_1698),
.B(n_1699),
.C(n_1689),
.Y(n_3809)
);

INVxp67_ASAP7_75t_L g3810 ( 
.A(n_3709),
.Y(n_3810)
);

AOI21xp5_ASAP7_75t_L g3811 ( 
.A1(n_3712),
.A2(n_1912),
.B(n_1889),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_L g3812 ( 
.A(n_3682),
.B(n_1700),
.Y(n_3812)
);

BUFx2_ASAP7_75t_L g3813 ( 
.A(n_3687),
.Y(n_3813)
);

OAI21x1_ASAP7_75t_L g3814 ( 
.A1(n_3676),
.A2(n_982),
.B(n_981),
.Y(n_3814)
);

INVxp67_ASAP7_75t_L g3815 ( 
.A(n_3718),
.Y(n_3815)
);

INVx2_ASAP7_75t_L g3816 ( 
.A(n_3679),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_L g3817 ( 
.A(n_3689),
.B(n_1704),
.Y(n_3817)
);

BUFx10_ASAP7_75t_L g3818 ( 
.A(n_3670),
.Y(n_3818)
);

AOI221xp5_ASAP7_75t_L g3819 ( 
.A1(n_3761),
.A2(n_1711),
.B1(n_1712),
.B2(n_1707),
.C(n_1706),
.Y(n_3819)
);

OAI22xp5_ASAP7_75t_L g3820 ( 
.A1(n_3771),
.A2(n_3665),
.B1(n_3672),
.B2(n_3737),
.Y(n_3820)
);

AOI22xp5_ASAP7_75t_L g3821 ( 
.A1(n_3775),
.A2(n_3739),
.B1(n_3715),
.B2(n_3720),
.Y(n_3821)
);

BUFx12f_ASAP7_75t_L g3822 ( 
.A(n_3764),
.Y(n_3822)
);

HB1xp67_ASAP7_75t_L g3823 ( 
.A(n_3757),
.Y(n_3823)
);

AND2x2_ASAP7_75t_L g3824 ( 
.A(n_3749),
.B(n_3669),
.Y(n_3824)
);

AOI22xp5_ASAP7_75t_L g3825 ( 
.A1(n_3791),
.A2(n_3734),
.B1(n_3677),
.B2(n_3741),
.Y(n_3825)
);

AOI22xp33_ASAP7_75t_L g3826 ( 
.A1(n_3770),
.A2(n_3723),
.B1(n_3733),
.B2(n_3729),
.Y(n_3826)
);

AOI22xp33_ASAP7_75t_L g3827 ( 
.A1(n_3773),
.A2(n_3695),
.B1(n_3699),
.B2(n_3693),
.Y(n_3827)
);

AOI22xp33_ASAP7_75t_L g3828 ( 
.A1(n_3747),
.A2(n_3688),
.B1(n_3718),
.B2(n_1725),
.Y(n_3828)
);

INVx2_ASAP7_75t_L g3829 ( 
.A(n_3765),
.Y(n_3829)
);

AOI22xp5_ASAP7_75t_L g3830 ( 
.A1(n_3746),
.A2(n_3802),
.B1(n_3753),
.B2(n_3786),
.Y(n_3830)
);

OAI222xp33_ASAP7_75t_L g3831 ( 
.A1(n_3805),
.A2(n_1732),
.B1(n_1726),
.B2(n_1734),
.C1(n_1728),
.C2(n_1718),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_3762),
.Y(n_3832)
);

OAI22x1_ASAP7_75t_L g3833 ( 
.A1(n_3766),
.A2(n_1744),
.B1(n_1747),
.B2(n_1742),
.Y(n_3833)
);

BUFx12f_ASAP7_75t_L g3834 ( 
.A(n_3758),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3768),
.Y(n_3835)
);

AND2x4_ASAP7_75t_L g3836 ( 
.A(n_3801),
.B(n_3668),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_3772),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3763),
.Y(n_3838)
);

OAI22xp33_ASAP7_75t_L g3839 ( 
.A1(n_3759),
.A2(n_3690),
.B1(n_3668),
.B2(n_2053),
.Y(n_3839)
);

BUFx10_ASAP7_75t_L g3840 ( 
.A(n_3785),
.Y(n_3840)
);

AOI22xp5_ASAP7_75t_L g3841 ( 
.A1(n_3816),
.A2(n_3690),
.B1(n_1750),
.B2(n_1752),
.Y(n_3841)
);

AOI21xp33_ASAP7_75t_L g3842 ( 
.A1(n_3809),
.A2(n_1754),
.B(n_1749),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3767),
.Y(n_3843)
);

AOI22xp33_ASAP7_75t_L g3844 ( 
.A1(n_3760),
.A2(n_1760),
.B1(n_1761),
.B2(n_1758),
.Y(n_3844)
);

OAI22xp33_ASAP7_75t_L g3845 ( 
.A1(n_3758),
.A2(n_2069),
.B1(n_1765),
.B2(n_1766),
.Y(n_3845)
);

AND2x2_ASAP7_75t_L g3846 ( 
.A(n_3769),
.B(n_4),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_3782),
.Y(n_3847)
);

INVx1_ASAP7_75t_L g3848 ( 
.A(n_3780),
.Y(n_3848)
);

HB1xp67_ASAP7_75t_L g3849 ( 
.A(n_3745),
.Y(n_3849)
);

INVx1_ASAP7_75t_SL g3850 ( 
.A(n_3807),
.Y(n_3850)
);

INVx1_ASAP7_75t_L g3851 ( 
.A(n_3808),
.Y(n_3851)
);

AOI22xp33_ASAP7_75t_L g3852 ( 
.A1(n_3778),
.A2(n_1770),
.B1(n_1775),
.B2(n_1763),
.Y(n_3852)
);

OR2x6_ASAP7_75t_L g3853 ( 
.A(n_3800),
.B(n_986),
.Y(n_3853)
);

AOI22xp33_ASAP7_75t_L g3854 ( 
.A1(n_3777),
.A2(n_1778),
.B1(n_1781),
.B2(n_1777),
.Y(n_3854)
);

HB1xp67_ASAP7_75t_L g3855 ( 
.A(n_3783),
.Y(n_3855)
);

NAND2xp5_ASAP7_75t_L g3856 ( 
.A(n_3803),
.B(n_1783),
.Y(n_3856)
);

AND2x2_ASAP7_75t_L g3857 ( 
.A(n_3797),
.B(n_6),
.Y(n_3857)
);

OAI22xp5_ASAP7_75t_L g3858 ( 
.A1(n_3788),
.A2(n_1785),
.B1(n_1786),
.B2(n_1784),
.Y(n_3858)
);

OAI21xp5_ASAP7_75t_L g3859 ( 
.A1(n_3799),
.A2(n_1789),
.B(n_1788),
.Y(n_3859)
);

OR2x2_ASAP7_75t_L g3860 ( 
.A(n_3810),
.B(n_10),
.Y(n_3860)
);

AOI22xp33_ASAP7_75t_SL g3861 ( 
.A1(n_3794),
.A2(n_1799),
.B1(n_1801),
.B2(n_1795),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_3808),
.Y(n_3862)
);

INVx2_ASAP7_75t_L g3863 ( 
.A(n_3756),
.Y(n_3863)
);

OAI21x1_ASAP7_75t_L g3864 ( 
.A1(n_3744),
.A2(n_989),
.B(n_988),
.Y(n_3864)
);

AOI22xp33_ASAP7_75t_L g3865 ( 
.A1(n_3751),
.A2(n_1807),
.B1(n_1808),
.B2(n_1803),
.Y(n_3865)
);

CKINVDCx6p67_ASAP7_75t_R g3866 ( 
.A(n_3776),
.Y(n_3866)
);

CKINVDCx11_ASAP7_75t_R g3867 ( 
.A(n_3818),
.Y(n_3867)
);

OAI222xp33_ASAP7_75t_L g3868 ( 
.A1(n_3774),
.A2(n_1825),
.B1(n_1813),
.B2(n_1829),
.C1(n_1823),
.C2(n_1812),
.Y(n_3868)
);

AOI22xp33_ASAP7_75t_L g3869 ( 
.A1(n_3795),
.A2(n_1837),
.B1(n_1838),
.B2(n_1835),
.Y(n_3869)
);

OA21x2_ASAP7_75t_L g3870 ( 
.A1(n_3779),
.A2(n_3798),
.B(n_3790),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3750),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3781),
.Y(n_3872)
);

OAI22xp33_ASAP7_75t_L g3873 ( 
.A1(n_3787),
.A2(n_2039),
.B1(n_2042),
.B2(n_2038),
.Y(n_3873)
);

INVx3_ASAP7_75t_L g3874 ( 
.A(n_3804),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3755),
.Y(n_3875)
);

OAI221xp5_ASAP7_75t_L g3876 ( 
.A1(n_3796),
.A2(n_1842),
.B1(n_1846),
.B2(n_1840),
.C(n_1839),
.Y(n_3876)
);

OAI21xp5_ASAP7_75t_L g3877 ( 
.A1(n_3789),
.A2(n_1848),
.B(n_1847),
.Y(n_3877)
);

NAND2x1p5_ASAP7_75t_L g3878 ( 
.A(n_3748),
.B(n_990),
.Y(n_3878)
);

AOI22xp33_ASAP7_75t_L g3879 ( 
.A1(n_3787),
.A2(n_1851),
.B1(n_1852),
.B2(n_1849),
.Y(n_3879)
);

OAI22xp5_ASAP7_75t_L g3880 ( 
.A1(n_3792),
.A2(n_1859),
.B1(n_1865),
.B2(n_1857),
.Y(n_3880)
);

NOR2xp33_ASAP7_75t_L g3881 ( 
.A(n_3815),
.B(n_1866),
.Y(n_3881)
);

OAI22xp33_ASAP7_75t_L g3882 ( 
.A1(n_3813),
.A2(n_3812),
.B1(n_3817),
.B2(n_3811),
.Y(n_3882)
);

INVxp67_ASAP7_75t_SL g3883 ( 
.A(n_3804),
.Y(n_3883)
);

HB1xp67_ASAP7_75t_L g3884 ( 
.A(n_3814),
.Y(n_3884)
);

AOI211xp5_ASAP7_75t_L g3885 ( 
.A1(n_3806),
.A2(n_1871),
.B(n_1874),
.C(n_1870),
.Y(n_3885)
);

AOI221xp5_ASAP7_75t_L g3886 ( 
.A1(n_3754),
.A2(n_2048),
.B1(n_2049),
.B2(n_2045),
.C(n_2043),
.Y(n_3886)
);

AOI21xp33_ASAP7_75t_L g3887 ( 
.A1(n_3784),
.A2(n_1884),
.B(n_1877),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3793),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3752),
.Y(n_3889)
);

AOI22xp33_ASAP7_75t_L g3890 ( 
.A1(n_3770),
.A2(n_1890),
.B1(n_1893),
.B2(n_1888),
.Y(n_3890)
);

AOI22xp5_ASAP7_75t_L g3891 ( 
.A1(n_3771),
.A2(n_1897),
.B1(n_1898),
.B2(n_1896),
.Y(n_3891)
);

AO22x1_ASAP7_75t_L g3892 ( 
.A1(n_3758),
.A2(n_1905),
.B1(n_1906),
.B2(n_1903),
.Y(n_3892)
);

INVx2_ASAP7_75t_L g3893 ( 
.A(n_3765),
.Y(n_3893)
);

INVx2_ASAP7_75t_L g3894 ( 
.A(n_3765),
.Y(n_3894)
);

NAND2xp5_ASAP7_75t_L g3895 ( 
.A(n_3749),
.B(n_1909),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3832),
.Y(n_3896)
);

BUFx2_ASAP7_75t_L g3897 ( 
.A(n_3823),
.Y(n_3897)
);

OAI21x1_ASAP7_75t_L g3898 ( 
.A1(n_3849),
.A2(n_10),
.B(n_11),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3835),
.Y(n_3899)
);

INVx2_ASAP7_75t_L g3900 ( 
.A(n_3829),
.Y(n_3900)
);

AOI22xp33_ASAP7_75t_L g3901 ( 
.A1(n_3889),
.A2(n_3875),
.B1(n_3820),
.B2(n_3882),
.Y(n_3901)
);

INVx2_ASAP7_75t_SL g3902 ( 
.A(n_3855),
.Y(n_3902)
);

BUFx6f_ASAP7_75t_L g3903 ( 
.A(n_3867),
.Y(n_3903)
);

BUFx6f_ASAP7_75t_L g3904 ( 
.A(n_3834),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3837),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_3838),
.Y(n_3906)
);

OR2x2_ASAP7_75t_L g3907 ( 
.A(n_3893),
.B(n_11),
.Y(n_3907)
);

NOR2xp33_ASAP7_75t_L g3908 ( 
.A(n_3847),
.B(n_1911),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_L g3909 ( 
.A(n_3894),
.B(n_1913),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3843),
.Y(n_3910)
);

BUFx10_ASAP7_75t_L g3911 ( 
.A(n_3888),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_3851),
.Y(n_3912)
);

HB1xp67_ASAP7_75t_L g3913 ( 
.A(n_3884),
.Y(n_3913)
);

OAI21x1_ASAP7_75t_L g3914 ( 
.A1(n_3864),
.A2(n_12),
.B(n_13),
.Y(n_3914)
);

AOI22xp33_ASAP7_75t_L g3915 ( 
.A1(n_3839),
.A2(n_2056),
.B1(n_2060),
.B2(n_2055),
.Y(n_3915)
);

AND2x2_ASAP7_75t_L g3916 ( 
.A(n_3824),
.B(n_13),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3862),
.Y(n_3917)
);

INVx2_ASAP7_75t_L g3918 ( 
.A(n_3871),
.Y(n_3918)
);

CKINVDCx5p33_ASAP7_75t_R g3919 ( 
.A(n_3866),
.Y(n_3919)
);

AND2x2_ASAP7_75t_L g3920 ( 
.A(n_3883),
.B(n_14),
.Y(n_3920)
);

OR2x2_ASAP7_75t_L g3921 ( 
.A(n_3850),
.B(n_14),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3872),
.Y(n_3922)
);

BUFx3_ASAP7_75t_L g3923 ( 
.A(n_3822),
.Y(n_3923)
);

AOI21x1_ASAP7_75t_L g3924 ( 
.A1(n_3895),
.A2(n_1929),
.B(n_1914),
.Y(n_3924)
);

CKINVDCx5p33_ASAP7_75t_R g3925 ( 
.A(n_3840),
.Y(n_3925)
);

HB1xp67_ASAP7_75t_L g3926 ( 
.A(n_3836),
.Y(n_3926)
);

INVx2_ASAP7_75t_L g3927 ( 
.A(n_3863),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3848),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3860),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3830),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3870),
.Y(n_3931)
);

INVx1_ASAP7_75t_L g3932 ( 
.A(n_3870),
.Y(n_3932)
);

HB1xp67_ASAP7_75t_L g3933 ( 
.A(n_3874),
.Y(n_3933)
);

INVx3_ASAP7_75t_L g3934 ( 
.A(n_3857),
.Y(n_3934)
);

OAI21x1_ASAP7_75t_L g3935 ( 
.A1(n_3821),
.A2(n_15),
.B(n_16),
.Y(n_3935)
);

BUFx4f_ASAP7_75t_SL g3936 ( 
.A(n_3846),
.Y(n_3936)
);

INVx2_ASAP7_75t_L g3937 ( 
.A(n_3833),
.Y(n_3937)
);

INVx2_ASAP7_75t_L g3938 ( 
.A(n_3856),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3881),
.Y(n_3939)
);

BUFx2_ASAP7_75t_L g3940 ( 
.A(n_3853),
.Y(n_3940)
);

AND2x2_ASAP7_75t_L g3941 ( 
.A(n_3825),
.B(n_15),
.Y(n_3941)
);

AND2x2_ASAP7_75t_L g3942 ( 
.A(n_3853),
.B(n_3878),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3841),
.Y(n_3943)
);

INVx2_ASAP7_75t_L g3944 ( 
.A(n_3892),
.Y(n_3944)
);

AOI21x1_ASAP7_75t_L g3945 ( 
.A1(n_3858),
.A2(n_1937),
.B(n_1932),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3827),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_L g3947 ( 
.A(n_3826),
.B(n_1938),
.Y(n_3947)
);

INVx2_ASAP7_75t_L g3948 ( 
.A(n_3876),
.Y(n_3948)
);

INVx2_ASAP7_75t_L g3949 ( 
.A(n_3880),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3861),
.Y(n_3950)
);

HB1xp67_ASAP7_75t_L g3951 ( 
.A(n_3831),
.Y(n_3951)
);

INVx2_ASAP7_75t_L g3952 ( 
.A(n_3891),
.Y(n_3952)
);

INVx1_ASAP7_75t_L g3953 ( 
.A(n_3844),
.Y(n_3953)
);

INVx1_ASAP7_75t_L g3954 ( 
.A(n_3859),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3877),
.Y(n_3955)
);

INVx3_ASAP7_75t_L g3956 ( 
.A(n_3873),
.Y(n_3956)
);

AOI21x1_ASAP7_75t_L g3957 ( 
.A1(n_3842),
.A2(n_1943),
.B(n_1940),
.Y(n_3957)
);

NAND2xp5_ASAP7_75t_L g3958 ( 
.A(n_3869),
.B(n_3819),
.Y(n_3958)
);

CKINVDCx11_ASAP7_75t_R g3959 ( 
.A(n_3845),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3828),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3879),
.Y(n_3961)
);

INVx2_ASAP7_75t_L g3962 ( 
.A(n_3885),
.Y(n_3962)
);

INVx2_ASAP7_75t_L g3963 ( 
.A(n_3854),
.Y(n_3963)
);

OAI22xp5_ASAP7_75t_L g3964 ( 
.A1(n_3901),
.A2(n_3890),
.B1(n_3852),
.B2(n_3865),
.Y(n_3964)
);

AOI22xp33_ASAP7_75t_L g3965 ( 
.A1(n_3951),
.A2(n_3886),
.B1(n_3887),
.B2(n_1953),
.Y(n_3965)
);

BUFx4f_ASAP7_75t_SL g3966 ( 
.A(n_3903),
.Y(n_3966)
);

AOI211xp5_ASAP7_75t_L g3967 ( 
.A1(n_3954),
.A2(n_3868),
.B(n_1958),
.C(n_1962),
.Y(n_3967)
);

AOI221xp5_ASAP7_75t_L g3968 ( 
.A1(n_3955),
.A2(n_1966),
.B1(n_1967),
.B2(n_1965),
.C(n_1944),
.Y(n_3968)
);

OAI221xp5_ASAP7_75t_L g3969 ( 
.A1(n_3947),
.A2(n_1976),
.B1(n_1977),
.B2(n_1975),
.C(n_1969),
.Y(n_3969)
);

INVx1_ASAP7_75t_L g3970 ( 
.A(n_3896),
.Y(n_3970)
);

OAI211xp5_ASAP7_75t_SL g3971 ( 
.A1(n_3930),
.A2(n_1980),
.B(n_1981),
.C(n_1978),
.Y(n_3971)
);

AOI22xp33_ASAP7_75t_L g3972 ( 
.A1(n_3948),
.A2(n_1990),
.B1(n_1992),
.B2(n_1988),
.Y(n_3972)
);

AOI22xp33_ASAP7_75t_L g3973 ( 
.A1(n_3959),
.A2(n_1999),
.B1(n_2001),
.B2(n_1997),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_L g3974 ( 
.A(n_3897),
.B(n_2006),
.Y(n_3974)
);

INVx2_ASAP7_75t_L g3975 ( 
.A(n_3899),
.Y(n_3975)
);

INVx1_ASAP7_75t_L g3976 ( 
.A(n_3905),
.Y(n_3976)
);

AOI22xp33_ASAP7_75t_L g3977 ( 
.A1(n_3962),
.A2(n_2011),
.B1(n_2022),
.B2(n_2008),
.Y(n_3977)
);

AOI22xp33_ASAP7_75t_L g3978 ( 
.A1(n_3946),
.A2(n_2033),
.B1(n_2036),
.B2(n_2029),
.Y(n_3978)
);

BUFx2_ASAP7_75t_L g3979 ( 
.A(n_3902),
.Y(n_3979)
);

AOI22xp33_ASAP7_75t_L g3980 ( 
.A1(n_3956),
.A2(n_2062),
.B1(n_2066),
.B2(n_2051),
.Y(n_3980)
);

OAI22xp33_ASAP7_75t_L g3981 ( 
.A1(n_3940),
.A2(n_1922),
.B1(n_1926),
.B2(n_1915),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3906),
.Y(n_3982)
);

INVx2_ASAP7_75t_L g3983 ( 
.A(n_3900),
.Y(n_3983)
);

OAI211xp5_ASAP7_75t_L g3984 ( 
.A1(n_3941),
.A2(n_1948),
.B(n_1979),
.C(n_1945),
.Y(n_3984)
);

AOI22xp33_ASAP7_75t_SL g3985 ( 
.A1(n_3936),
.A2(n_1984),
.B1(n_1985),
.B2(n_1982),
.Y(n_3985)
);

AND2x2_ASAP7_75t_L g3986 ( 
.A(n_3926),
.B(n_16),
.Y(n_3986)
);

AND2x2_ASAP7_75t_L g3987 ( 
.A(n_3933),
.B(n_3929),
.Y(n_3987)
);

AND2x2_ASAP7_75t_L g3988 ( 
.A(n_3912),
.B(n_17),
.Y(n_3988)
);

INVx2_ASAP7_75t_L g3989 ( 
.A(n_3918),
.Y(n_3989)
);

AND2x2_ASAP7_75t_L g3990 ( 
.A(n_3917),
.B(n_17),
.Y(n_3990)
);

CKINVDCx6p67_ASAP7_75t_R g3991 ( 
.A(n_3903),
.Y(n_3991)
);

AOI22xp33_ASAP7_75t_L g3992 ( 
.A1(n_3949),
.A2(n_1993),
.B1(n_2002),
.B2(n_1986),
.Y(n_3992)
);

OAI22xp5_ASAP7_75t_SL g3993 ( 
.A1(n_3919),
.A2(n_2025),
.B1(n_2027),
.B2(n_2004),
.Y(n_3993)
);

INVx1_ASAP7_75t_L g3994 ( 
.A(n_3928),
.Y(n_3994)
);

INVx1_ASAP7_75t_L g3995 ( 
.A(n_3910),
.Y(n_3995)
);

AOI22xp5_ASAP7_75t_L g3996 ( 
.A1(n_3944),
.A2(n_2035),
.B1(n_2040),
.B2(n_2030),
.Y(n_3996)
);

AOI22xp33_ASAP7_75t_L g3997 ( 
.A1(n_3950),
.A2(n_2054),
.B1(n_20),
.B2(n_18),
.Y(n_3997)
);

OAI211xp5_ASAP7_75t_SL g3998 ( 
.A1(n_3961),
.A2(n_20),
.B(n_18),
.C(n_19),
.Y(n_3998)
);

NOR3xp33_ASAP7_75t_L g3999 ( 
.A(n_3958),
.B(n_21),
.C(n_22),
.Y(n_3999)
);

NOR2x1_ASAP7_75t_SL g4000 ( 
.A(n_3931),
.B(n_3932),
.Y(n_4000)
);

OR2x2_ASAP7_75t_L g4001 ( 
.A(n_3913),
.B(n_21),
.Y(n_4001)
);

AO31x2_ASAP7_75t_L g4002 ( 
.A1(n_3922),
.A2(n_24),
.A3(n_22),
.B(n_23),
.Y(n_4002)
);

OAI22xp5_ASAP7_75t_L g4003 ( 
.A1(n_3953),
.A2(n_26),
.B1(n_23),
.B2(n_25),
.Y(n_4003)
);

A2O1A1Ixp33_ASAP7_75t_L g4004 ( 
.A1(n_3935),
.A2(n_35),
.B(n_43),
.C(n_26),
.Y(n_4004)
);

INVx3_ASAP7_75t_L g4005 ( 
.A(n_3904),
.Y(n_4005)
);

AOI21xp33_ASAP7_75t_L g4006 ( 
.A1(n_3937),
.A2(n_27),
.B(n_28),
.Y(n_4006)
);

INVx2_ASAP7_75t_L g4007 ( 
.A(n_3927),
.Y(n_4007)
);

INVx2_ASAP7_75t_L g4008 ( 
.A(n_3907),
.Y(n_4008)
);

AND2x6_ASAP7_75t_SL g4009 ( 
.A(n_3939),
.B(n_28),
.Y(n_4009)
);

AOI22xp33_ASAP7_75t_L g4010 ( 
.A1(n_3963),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_4010)
);

AOI22xp33_ASAP7_75t_L g4011 ( 
.A1(n_3952),
.A2(n_32),
.B1(n_29),
.B2(n_31),
.Y(n_4011)
);

INVx1_ASAP7_75t_L g4012 ( 
.A(n_3909),
.Y(n_4012)
);

INVx4_ASAP7_75t_L g4013 ( 
.A(n_3925),
.Y(n_4013)
);

OAI22xp33_ASAP7_75t_L g4014 ( 
.A1(n_3938),
.A2(n_36),
.B1(n_32),
.B2(n_34),
.Y(n_4014)
);

AOI33xp33_ASAP7_75t_L g4015 ( 
.A1(n_3960),
.A2(n_38),
.A3(n_40),
.B1(n_36),
.B2(n_37),
.B3(n_39),
.Y(n_4015)
);

INVx1_ASAP7_75t_L g4016 ( 
.A(n_3934),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_3921),
.Y(n_4017)
);

OAI211xp5_ASAP7_75t_L g4018 ( 
.A1(n_3915),
.A2(n_41),
.B(n_38),
.C(n_40),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_3920),
.B(n_41),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_3898),
.Y(n_4020)
);

AOI22xp33_ASAP7_75t_SL g4021 ( 
.A1(n_3942),
.A2(n_45),
.B1(n_42),
.B2(n_43),
.Y(n_4021)
);

OAI22xp5_ASAP7_75t_L g4022 ( 
.A1(n_3943),
.A2(n_46),
.B1(n_42),
.B2(n_45),
.Y(n_4022)
);

INVx1_ASAP7_75t_L g4023 ( 
.A(n_3916),
.Y(n_4023)
);

A2O1A1Ixp33_ASAP7_75t_L g4024 ( 
.A1(n_3914),
.A2(n_56),
.B(n_64),
.C(n_47),
.Y(n_4024)
);

AOI22xp33_ASAP7_75t_L g4025 ( 
.A1(n_3904),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_4025)
);

OR2x6_ASAP7_75t_L g4026 ( 
.A(n_3923),
.B(n_48),
.Y(n_4026)
);

OAI211xp5_ASAP7_75t_L g4027 ( 
.A1(n_3924),
.A2(n_52),
.B(n_49),
.C(n_51),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_3908),
.Y(n_4028)
);

AOI22xp33_ASAP7_75t_L g4029 ( 
.A1(n_3911),
.A2(n_55),
.B1(n_52),
.B2(n_54),
.Y(n_4029)
);

OAI22xp5_ASAP7_75t_L g4030 ( 
.A1(n_3945),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_4030)
);

OAI22xp5_ASAP7_75t_L g4031 ( 
.A1(n_3957),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_4031)
);

INVx2_ASAP7_75t_L g4032 ( 
.A(n_3897),
.Y(n_4032)
);

NAND3xp33_ASAP7_75t_L g4033 ( 
.A(n_3954),
.B(n_59),
.C(n_60),
.Y(n_4033)
);

OAI22xp5_ASAP7_75t_L g4034 ( 
.A1(n_3901),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_4034)
);

AO22x1_ASAP7_75t_L g4035 ( 
.A1(n_3930),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_4035)
);

INVx1_ASAP7_75t_L g4036 ( 
.A(n_3896),
.Y(n_4036)
);

AOI221xp5_ASAP7_75t_L g4037 ( 
.A1(n_3951),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.C(n_66),
.Y(n_4037)
);

AND2x2_ASAP7_75t_L g4038 ( 
.A(n_3926),
.B(n_65),
.Y(n_4038)
);

BUFx4f_ASAP7_75t_SL g4039 ( 
.A(n_3903),
.Y(n_4039)
);

AOI22xp33_ASAP7_75t_L g4040 ( 
.A1(n_3951),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_4040)
);

HB1xp67_ASAP7_75t_L g4041 ( 
.A(n_3913),
.Y(n_4041)
);

AOI22xp33_ASAP7_75t_SL g4042 ( 
.A1(n_3951),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_4042)
);

AND2x2_ASAP7_75t_L g4043 ( 
.A(n_3926),
.B(n_69),
.Y(n_4043)
);

AOI21xp33_ASAP7_75t_SL g4044 ( 
.A1(n_3951),
.A2(n_70),
.B(n_71),
.Y(n_4044)
);

INVx2_ASAP7_75t_L g4045 ( 
.A(n_3897),
.Y(n_4045)
);

AND2x4_ASAP7_75t_L g4046 ( 
.A(n_3897),
.B(n_70),
.Y(n_4046)
);

OR2x2_ASAP7_75t_L g4047 ( 
.A(n_3897),
.B(n_71),
.Y(n_4047)
);

AND2x4_ASAP7_75t_SL g4048 ( 
.A(n_3903),
.B(n_73),
.Y(n_4048)
);

AOI22xp33_ASAP7_75t_L g4049 ( 
.A1(n_3951),
.A2(n_78),
.B1(n_75),
.B2(n_77),
.Y(n_4049)
);

INVx2_ASAP7_75t_L g4050 ( 
.A(n_3897),
.Y(n_4050)
);

AOI22xp33_ASAP7_75t_L g4051 ( 
.A1(n_3951),
.A2(n_78),
.B1(n_75),
.B2(n_77),
.Y(n_4051)
);

OAI22xp5_ASAP7_75t_L g4052 ( 
.A1(n_3901),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_4052)
);

OAI211xp5_ASAP7_75t_L g4053 ( 
.A1(n_3951),
.A2(n_83),
.B(n_80),
.C(n_81),
.Y(n_4053)
);

INVx3_ASAP7_75t_L g4054 ( 
.A(n_3904),
.Y(n_4054)
);

AOI22xp33_ASAP7_75t_L g4055 ( 
.A1(n_3951),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_4055)
);

AOI21x1_ASAP7_75t_L g4056 ( 
.A1(n_3946),
.A2(n_85),
.B(n_86),
.Y(n_4056)
);

OAI211xp5_ASAP7_75t_L g4057 ( 
.A1(n_3951),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_4057)
);

AOI22xp33_ASAP7_75t_L g4058 ( 
.A1(n_3951),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_4058)
);

AND2x2_ASAP7_75t_L g4059 ( 
.A(n_3926),
.B(n_90),
.Y(n_4059)
);

INVx1_ASAP7_75t_L g4060 ( 
.A(n_3896),
.Y(n_4060)
);

INVx3_ASAP7_75t_L g4061 ( 
.A(n_3904),
.Y(n_4061)
);

OAI221xp5_ASAP7_75t_L g4062 ( 
.A1(n_3901),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.C(n_95),
.Y(n_4062)
);

AOI22xp33_ASAP7_75t_L g4063 ( 
.A1(n_3951),
.A2(n_96),
.B1(n_91),
.B2(n_95),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_3896),
.Y(n_4064)
);

AOI22xp33_ASAP7_75t_L g4065 ( 
.A1(n_3951),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_4065)
);

OA21x2_ASAP7_75t_L g4066 ( 
.A1(n_3931),
.A2(n_99),
.B(n_100),
.Y(n_4066)
);

AOI22xp33_ASAP7_75t_L g4067 ( 
.A1(n_3951),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_4067)
);

AOI22xp33_ASAP7_75t_L g4068 ( 
.A1(n_3951),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_4068)
);

BUFx2_ASAP7_75t_L g4069 ( 
.A(n_3897),
.Y(n_4069)
);

AOI221xp5_ASAP7_75t_L g4070 ( 
.A1(n_3951),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.C(n_109),
.Y(n_4070)
);

AOI22xp33_ASAP7_75t_L g4071 ( 
.A1(n_3951),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_4071)
);

AOI22xp33_ASAP7_75t_SL g4072 ( 
.A1(n_3951),
.A2(n_112),
.B1(n_110),
.B2(n_111),
.Y(n_4072)
);

AOI22xp33_ASAP7_75t_L g4073 ( 
.A1(n_3951),
.A2(n_114),
.B1(n_111),
.B2(n_113),
.Y(n_4073)
);

AOI22xp33_ASAP7_75t_L g4074 ( 
.A1(n_3951),
.A2(n_116),
.B1(n_113),
.B2(n_114),
.Y(n_4074)
);

OAI22xp5_ASAP7_75t_L g4075 ( 
.A1(n_3901),
.A2(n_119),
.B1(n_116),
.B2(n_117),
.Y(n_4075)
);

AOI22xp5_ASAP7_75t_L g4076 ( 
.A1(n_3951),
.A2(n_121),
.B1(n_117),
.B2(n_120),
.Y(n_4076)
);

AOI22xp33_ASAP7_75t_L g4077 ( 
.A1(n_3951),
.A2(n_125),
.B1(n_120),
.B2(n_122),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_3896),
.Y(n_4078)
);

AOI22xp33_ASAP7_75t_L g4079 ( 
.A1(n_3951),
.A2(n_126),
.B1(n_122),
.B2(n_125),
.Y(n_4079)
);

OAI22xp5_ASAP7_75t_L g4080 ( 
.A1(n_3901),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_4080)
);

AOI221xp5_ASAP7_75t_L g4081 ( 
.A1(n_3951),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.C(n_130),
.Y(n_4081)
);

AND2x2_ASAP7_75t_L g4082 ( 
.A(n_4069),
.B(n_129),
.Y(n_4082)
);

INVx1_ASAP7_75t_L g4083 ( 
.A(n_3976),
.Y(n_4083)
);

INVx2_ASAP7_75t_L g4084 ( 
.A(n_4000),
.Y(n_4084)
);

INVx2_ASAP7_75t_L g4085 ( 
.A(n_4007),
.Y(n_4085)
);

OAI211xp5_ASAP7_75t_SL g4086 ( 
.A1(n_3973),
.A2(n_132),
.B(n_130),
.C(n_131),
.Y(n_4086)
);

NAND2xp5_ASAP7_75t_L g4087 ( 
.A(n_4020),
.B(n_133),
.Y(n_4087)
);

AND2x2_ASAP7_75t_L g4088 ( 
.A(n_3979),
.B(n_133),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_3982),
.Y(n_4089)
);

INVx1_ASAP7_75t_L g4090 ( 
.A(n_3970),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_4036),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_4060),
.Y(n_4092)
);

AOI22xp33_ASAP7_75t_L g4093 ( 
.A1(n_3999),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_4064),
.Y(n_4094)
);

AND2x2_ASAP7_75t_L g4095 ( 
.A(n_4032),
.B(n_136),
.Y(n_4095)
);

HB1xp67_ASAP7_75t_L g4096 ( 
.A(n_4041),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_4012),
.B(n_137),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_4078),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_L g4099 ( 
.A(n_4008),
.B(n_138),
.Y(n_4099)
);

INVxp67_ASAP7_75t_L g4100 ( 
.A(n_4045),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3994),
.Y(n_4101)
);

OR2x2_ASAP7_75t_L g4102 ( 
.A(n_4017),
.B(n_138),
.Y(n_4102)
);

BUFx2_ASAP7_75t_L g4103 ( 
.A(n_4050),
.Y(n_4103)
);

AND2x2_ASAP7_75t_L g4104 ( 
.A(n_3987),
.B(n_139),
.Y(n_4104)
);

AND2x2_ASAP7_75t_L g4105 ( 
.A(n_4016),
.B(n_139),
.Y(n_4105)
);

AND2x2_ASAP7_75t_L g4106 ( 
.A(n_4023),
.B(n_140),
.Y(n_4106)
);

AND2x2_ASAP7_75t_L g4107 ( 
.A(n_3983),
.B(n_140),
.Y(n_4107)
);

INVx1_ASAP7_75t_L g4108 ( 
.A(n_3975),
.Y(n_4108)
);

HB1xp67_ASAP7_75t_L g4109 ( 
.A(n_4066),
.Y(n_4109)
);

AND2x2_ASAP7_75t_L g4110 ( 
.A(n_3989),
.B(n_141),
.Y(n_4110)
);

AND2x2_ASAP7_75t_L g4111 ( 
.A(n_3988),
.B(n_141),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_3995),
.Y(n_4112)
);

INVxp67_ASAP7_75t_SL g4113 ( 
.A(n_4066),
.Y(n_4113)
);

AND2x2_ASAP7_75t_L g4114 ( 
.A(n_3990),
.B(n_142),
.Y(n_4114)
);

AND2x2_ASAP7_75t_L g4115 ( 
.A(n_4046),
.B(n_142),
.Y(n_4115)
);

NAND2xp5_ASAP7_75t_L g4116 ( 
.A(n_3986),
.B(n_143),
.Y(n_4116)
);

AND2x2_ASAP7_75t_L g4117 ( 
.A(n_4038),
.B(n_145),
.Y(n_4117)
);

OR2x2_ASAP7_75t_L g4118 ( 
.A(n_4047),
.B(n_145),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_4002),
.Y(n_4119)
);

INVx5_ASAP7_75t_SL g4120 ( 
.A(n_3991),
.Y(n_4120)
);

INVx1_ASAP7_75t_L g4121 ( 
.A(n_4002),
.Y(n_4121)
);

OAI221xp5_ASAP7_75t_L g4122 ( 
.A1(n_4076),
.A2(n_149),
.B1(n_146),
.B2(n_148),
.C(n_150),
.Y(n_4122)
);

INVxp67_ASAP7_75t_R g4123 ( 
.A(n_3966),
.Y(n_4123)
);

BUFx6f_ASAP7_75t_L g4124 ( 
.A(n_4005),
.Y(n_4124)
);

INVx2_ASAP7_75t_L g4125 ( 
.A(n_4001),
.Y(n_4125)
);

AND2x4_ASAP7_75t_L g4126 ( 
.A(n_4054),
.B(n_146),
.Y(n_4126)
);

AND2x2_ASAP7_75t_L g4127 ( 
.A(n_4043),
.B(n_148),
.Y(n_4127)
);

OR2x2_ASAP7_75t_L g4128 ( 
.A(n_3974),
.B(n_149),
.Y(n_4128)
);

NAND2xp5_ASAP7_75t_L g4129 ( 
.A(n_4059),
.B(n_150),
.Y(n_4129)
);

OR2x6_ASAP7_75t_L g4130 ( 
.A(n_4026),
.B(n_151),
.Y(n_4130)
);

INVx2_ASAP7_75t_L g4131 ( 
.A(n_4061),
.Y(n_4131)
);

INVx2_ASAP7_75t_L g4132 ( 
.A(n_4002),
.Y(n_4132)
);

INVx2_ASAP7_75t_L g4133 ( 
.A(n_4056),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_SL g4134 ( 
.A(n_4013),
.B(n_151),
.Y(n_4134)
);

HB1xp67_ASAP7_75t_L g4135 ( 
.A(n_4019),
.Y(n_4135)
);

INVx2_ASAP7_75t_L g4136 ( 
.A(n_4028),
.Y(n_4136)
);

AOI22xp33_ASAP7_75t_L g4137 ( 
.A1(n_4037),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_4033),
.Y(n_4138)
);

AND2x2_ASAP7_75t_L g4139 ( 
.A(n_4026),
.B(n_152),
.Y(n_4139)
);

INVx2_ASAP7_75t_L g4140 ( 
.A(n_4009),
.Y(n_4140)
);

HB1xp67_ASAP7_75t_L g4141 ( 
.A(n_4035),
.Y(n_4141)
);

NOR2x1_ASAP7_75t_SL g4142 ( 
.A(n_4053),
.B(n_153),
.Y(n_4142)
);

AND2x2_ASAP7_75t_L g4143 ( 
.A(n_4048),
.B(n_154),
.Y(n_4143)
);

AND2x4_ASAP7_75t_L g4144 ( 
.A(n_4004),
.B(n_4024),
.Y(n_4144)
);

AND2x2_ASAP7_75t_L g4145 ( 
.A(n_4044),
.B(n_155),
.Y(n_4145)
);

INVx2_ASAP7_75t_L g4146 ( 
.A(n_4039),
.Y(n_4146)
);

AND2x2_ASAP7_75t_L g4147 ( 
.A(n_3980),
.B(n_157),
.Y(n_4147)
);

INVx2_ASAP7_75t_L g4148 ( 
.A(n_3996),
.Y(n_4148)
);

OR2x2_ASAP7_75t_L g4149 ( 
.A(n_4006),
.B(n_157),
.Y(n_4149)
);

NOR2xp33_ASAP7_75t_L g4150 ( 
.A(n_3984),
.B(n_3969),
.Y(n_4150)
);

OR2x2_ASAP7_75t_L g4151 ( 
.A(n_4003),
.B(n_158),
.Y(n_4151)
);

INVx2_ASAP7_75t_L g4152 ( 
.A(n_4030),
.Y(n_4152)
);

INVx3_ASAP7_75t_L g4153 ( 
.A(n_3981),
.Y(n_4153)
);

BUFx3_ASAP7_75t_L g4154 ( 
.A(n_3993),
.Y(n_4154)
);

INVx2_ASAP7_75t_L g4155 ( 
.A(n_4031),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_4015),
.Y(n_4156)
);

INVx2_ASAP7_75t_L g4157 ( 
.A(n_4062),
.Y(n_4157)
);

INVx1_ASAP7_75t_L g4158 ( 
.A(n_4057),
.Y(n_4158)
);

INVx2_ASAP7_75t_L g4159 ( 
.A(n_4034),
.Y(n_4159)
);

AND2x2_ASAP7_75t_L g4160 ( 
.A(n_4021),
.B(n_158),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_4014),
.Y(n_4161)
);

INVx2_ASAP7_75t_L g4162 ( 
.A(n_4052),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_4027),
.Y(n_4163)
);

BUFx3_ASAP7_75t_L g4164 ( 
.A(n_4075),
.Y(n_4164)
);

BUFx2_ASAP7_75t_L g4165 ( 
.A(n_4070),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_4022),
.Y(n_4166)
);

INVx3_ASAP7_75t_L g4167 ( 
.A(n_4042),
.Y(n_4167)
);

INVx2_ASAP7_75t_L g4168 ( 
.A(n_4080),
.Y(n_4168)
);

AND2x2_ASAP7_75t_L g4169 ( 
.A(n_4072),
.B(n_159),
.Y(n_4169)
);

BUFx2_ASAP7_75t_L g4170 ( 
.A(n_4081),
.Y(n_4170)
);

INVxp67_ASAP7_75t_R g4171 ( 
.A(n_3964),
.Y(n_4171)
);

INVx2_ASAP7_75t_L g4172 ( 
.A(n_3998),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_4018),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4040),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_L g4175 ( 
.A(n_3972),
.B(n_160),
.Y(n_4175)
);

OR2x2_ASAP7_75t_L g4176 ( 
.A(n_4049),
.B(n_161),
.Y(n_4176)
);

INVx2_ASAP7_75t_L g4177 ( 
.A(n_3971),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_4051),
.Y(n_4178)
);

AND2x2_ASAP7_75t_L g4179 ( 
.A(n_4055),
.B(n_4058),
.Y(n_4179)
);

INVx2_ASAP7_75t_L g4180 ( 
.A(n_4063),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_4065),
.Y(n_4181)
);

OR2x2_ASAP7_75t_L g4182 ( 
.A(n_4067),
.B(n_162),
.Y(n_4182)
);

NOR2x1_ASAP7_75t_SL g4183 ( 
.A(n_3985),
.B(n_162),
.Y(n_4183)
);

BUFx3_ASAP7_75t_L g4184 ( 
.A(n_4025),
.Y(n_4184)
);

BUFx6f_ASAP7_75t_L g4185 ( 
.A(n_3977),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_4068),
.Y(n_4186)
);

OR2x2_ASAP7_75t_L g4187 ( 
.A(n_4071),
.B(n_4073),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_4074),
.Y(n_4188)
);

INVx2_ASAP7_75t_L g4189 ( 
.A(n_4077),
.Y(n_4189)
);

AND2x2_ASAP7_75t_L g4190 ( 
.A(n_4079),
.B(n_163),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_L g4191 ( 
.A(n_3997),
.B(n_164),
.Y(n_4191)
);

OR2x2_ASAP7_75t_L g4192 ( 
.A(n_4010),
.B(n_165),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_L g4193 ( 
.A(n_3978),
.B(n_165),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_4011),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_L g4195 ( 
.A(n_3968),
.B(n_166),
.Y(n_4195)
);

INVx2_ASAP7_75t_L g4196 ( 
.A(n_3992),
.Y(n_4196)
);

OR2x2_ASAP7_75t_L g4197 ( 
.A(n_4029),
.B(n_166),
.Y(n_4197)
);

NOR2xp33_ASAP7_75t_R g4198 ( 
.A(n_3965),
.B(n_169),
.Y(n_4198)
);

INVx1_ASAP7_75t_SL g4199 ( 
.A(n_3967),
.Y(n_4199)
);

INVx2_ASAP7_75t_L g4200 ( 
.A(n_4000),
.Y(n_4200)
);

INVx2_ASAP7_75t_L g4201 ( 
.A(n_4000),
.Y(n_4201)
);

HB1xp67_ASAP7_75t_L g4202 ( 
.A(n_4041),
.Y(n_4202)
);

INVx2_ASAP7_75t_L g4203 ( 
.A(n_4000),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_3976),
.Y(n_4204)
);

AND2x2_ASAP7_75t_L g4205 ( 
.A(n_4069),
.B(n_168),
.Y(n_4205)
);

INVx2_ASAP7_75t_L g4206 ( 
.A(n_4000),
.Y(n_4206)
);

HB1xp67_ASAP7_75t_L g4207 ( 
.A(n_4041),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_4020),
.B(n_170),
.Y(n_4208)
);

HB1xp67_ASAP7_75t_L g4209 ( 
.A(n_4041),
.Y(n_4209)
);

AND2x2_ASAP7_75t_L g4210 ( 
.A(n_4069),
.B(n_171),
.Y(n_4210)
);

AND2x2_ASAP7_75t_L g4211 ( 
.A(n_4069),
.B(n_171),
.Y(n_4211)
);

NAND2xp5_ASAP7_75t_L g4212 ( 
.A(n_4020),
.B(n_172),
.Y(n_4212)
);

INVx2_ASAP7_75t_L g4213 ( 
.A(n_4000),
.Y(n_4213)
);

AND2x2_ASAP7_75t_L g4214 ( 
.A(n_4069),
.B(n_173),
.Y(n_4214)
);

AND2x2_ASAP7_75t_L g4215 ( 
.A(n_4069),
.B(n_173),
.Y(n_4215)
);

AND2x4_ASAP7_75t_L g4216 ( 
.A(n_4069),
.B(n_174),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_L g4217 ( 
.A(n_4020),
.B(n_174),
.Y(n_4217)
);

NAND2xp5_ASAP7_75t_L g4218 ( 
.A(n_4020),
.B(n_175),
.Y(n_4218)
);

INVx2_ASAP7_75t_L g4219 ( 
.A(n_4000),
.Y(n_4219)
);

AND2x2_ASAP7_75t_L g4220 ( 
.A(n_4069),
.B(n_175),
.Y(n_4220)
);

INVx2_ASAP7_75t_L g4221 ( 
.A(n_4000),
.Y(n_4221)
);

AOI221xp5_ASAP7_75t_L g4222 ( 
.A1(n_3999),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.C(n_179),
.Y(n_4222)
);

AO21x2_ASAP7_75t_L g4223 ( 
.A1(n_4000),
.A2(n_176),
.B(n_177),
.Y(n_4223)
);

AND2x2_ASAP7_75t_L g4224 ( 
.A(n_4069),
.B(n_178),
.Y(n_4224)
);

NAND2xp5_ASAP7_75t_L g4225 ( 
.A(n_4020),
.B(n_179),
.Y(n_4225)
);

AOI22xp5_ASAP7_75t_L g4226 ( 
.A1(n_3999),
.A2(n_183),
.B1(n_180),
.B2(n_181),
.Y(n_4226)
);

HB1xp67_ASAP7_75t_L g4227 ( 
.A(n_4041),
.Y(n_4227)
);

AND2x2_ASAP7_75t_L g4228 ( 
.A(n_4069),
.B(n_180),
.Y(n_4228)
);

NAND2xp5_ASAP7_75t_L g4229 ( 
.A(n_4020),
.B(n_181),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_3976),
.Y(n_4230)
);

AOI22xp5_ASAP7_75t_L g4231 ( 
.A1(n_3999),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.Y(n_4231)
);

NAND2x1p5_ASAP7_75t_L g4232 ( 
.A(n_4069),
.B(n_184),
.Y(n_4232)
);

AND2x2_ASAP7_75t_L g4233 ( 
.A(n_4069),
.B(n_185),
.Y(n_4233)
);

AND2x2_ASAP7_75t_L g4234 ( 
.A(n_4069),
.B(n_186),
.Y(n_4234)
);

INVx1_ASAP7_75t_L g4235 ( 
.A(n_3976),
.Y(n_4235)
);

AND2x2_ASAP7_75t_L g4236 ( 
.A(n_4069),
.B(n_186),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_3976),
.Y(n_4237)
);

INVx2_ASAP7_75t_L g4238 ( 
.A(n_4000),
.Y(n_4238)
);

AOI22xp33_ASAP7_75t_L g4239 ( 
.A1(n_3999),
.A2(n_191),
.B1(n_189),
.B2(n_190),
.Y(n_4239)
);

NAND2xp5_ASAP7_75t_L g4240 ( 
.A(n_4020),
.B(n_191),
.Y(n_4240)
);

NOR2xp33_ASAP7_75t_L g4241 ( 
.A(n_3991),
.B(n_193),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_3976),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_3976),
.Y(n_4243)
);

INVx1_ASAP7_75t_L g4244 ( 
.A(n_4083),
.Y(n_4244)
);

INVx2_ASAP7_75t_L g4245 ( 
.A(n_4131),
.Y(n_4245)
);

AOI31xp33_ASAP7_75t_L g4246 ( 
.A1(n_4141),
.A2(n_196),
.A3(n_194),
.B(n_195),
.Y(n_4246)
);

AND2x2_ASAP7_75t_L g4247 ( 
.A(n_4135),
.B(n_194),
.Y(n_4247)
);

NAND4xp25_ASAP7_75t_L g4248 ( 
.A(n_4165),
.B(n_197),
.C(n_198),
.D(n_196),
.Y(n_4248)
);

INVx1_ASAP7_75t_L g4249 ( 
.A(n_4089),
.Y(n_4249)
);

AOI22xp33_ASAP7_75t_L g4250 ( 
.A1(n_4170),
.A2(n_199),
.B1(n_195),
.B2(n_197),
.Y(n_4250)
);

AND2x2_ASAP7_75t_L g4251 ( 
.A(n_4103),
.B(n_199),
.Y(n_4251)
);

OA21x2_ASAP7_75t_L g4252 ( 
.A1(n_4113),
.A2(n_200),
.B(n_201),
.Y(n_4252)
);

AND2x2_ASAP7_75t_L g4253 ( 
.A(n_4136),
.B(n_200),
.Y(n_4253)
);

INVx2_ASAP7_75t_L g4254 ( 
.A(n_4124),
.Y(n_4254)
);

AND2x2_ASAP7_75t_L g4255 ( 
.A(n_4125),
.B(n_4100),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_4090),
.Y(n_4256)
);

NAND3xp33_ASAP7_75t_L g4257 ( 
.A(n_4222),
.B(n_202),
.C(n_203),
.Y(n_4257)
);

AOI33xp33_ASAP7_75t_L g4258 ( 
.A1(n_4158),
.A2(n_206),
.A3(n_208),
.B1(n_204),
.B2(n_205),
.B3(n_207),
.Y(n_4258)
);

NAND2xp5_ASAP7_75t_L g4259 ( 
.A(n_4138),
.B(n_4152),
.Y(n_4259)
);

OAI221xp5_ASAP7_75t_L g4260 ( 
.A1(n_4167),
.A2(n_207),
.B1(n_204),
.B2(n_206),
.C(n_209),
.Y(n_4260)
);

INVx2_ASAP7_75t_L g4261 ( 
.A(n_4124),
.Y(n_4261)
);

OAI33xp33_ASAP7_75t_L g4262 ( 
.A1(n_4156),
.A2(n_211),
.A3(n_213),
.B1(n_209),
.B2(n_210),
.B3(n_212),
.Y(n_4262)
);

OA21x2_ASAP7_75t_L g4263 ( 
.A1(n_4084),
.A2(n_210),
.B(n_211),
.Y(n_4263)
);

OAI211xp5_ASAP7_75t_SL g4264 ( 
.A1(n_4199),
.A2(n_215),
.B(n_213),
.C(n_214),
.Y(n_4264)
);

OAI211xp5_ASAP7_75t_L g4265 ( 
.A1(n_4226),
.A2(n_217),
.B(n_215),
.C(n_216),
.Y(n_4265)
);

OAI221xp5_ASAP7_75t_L g4266 ( 
.A1(n_4140),
.A2(n_221),
.B1(n_218),
.B2(n_219),
.C(n_222),
.Y(n_4266)
);

AND2x2_ASAP7_75t_L g4267 ( 
.A(n_4096),
.B(n_218),
.Y(n_4267)
);

AOI221xp5_ASAP7_75t_L g4268 ( 
.A1(n_4144),
.A2(n_224),
.B1(n_221),
.B2(n_223),
.C(n_225),
.Y(n_4268)
);

HB1xp67_ASAP7_75t_L g4269 ( 
.A(n_4202),
.Y(n_4269)
);

INVx1_ASAP7_75t_L g4270 ( 
.A(n_4091),
.Y(n_4270)
);

AOI21xp5_ASAP7_75t_L g4271 ( 
.A1(n_4171),
.A2(n_225),
.B(n_226),
.Y(n_4271)
);

OAI33xp33_ASAP7_75t_L g4272 ( 
.A1(n_4163),
.A2(n_4121),
.A3(n_4119),
.B1(n_4173),
.B2(n_4161),
.B3(n_4174),
.Y(n_4272)
);

AOI22xp33_ASAP7_75t_L g4273 ( 
.A1(n_4164),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_L g4274 ( 
.A(n_4155),
.B(n_227),
.Y(n_4274)
);

AOI221xp5_ASAP7_75t_L g4275 ( 
.A1(n_4157),
.A2(n_4109),
.B1(n_4122),
.B2(n_4181),
.C(n_4178),
.Y(n_4275)
);

OAI22xp5_ASAP7_75t_L g4276 ( 
.A1(n_4231),
.A2(n_231),
.B1(n_229),
.B2(n_230),
.Y(n_4276)
);

AOI22xp5_ASAP7_75t_L g4277 ( 
.A1(n_4172),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_4277)
);

AOI22xp33_ASAP7_75t_L g4278 ( 
.A1(n_4179),
.A2(n_234),
.B1(n_232),
.B2(n_233),
.Y(n_4278)
);

AND2x2_ASAP7_75t_L g4279 ( 
.A(n_4207),
.B(n_4209),
.Y(n_4279)
);

INVx4_ASAP7_75t_R g4280 ( 
.A(n_4123),
.Y(n_4280)
);

AOI21xp33_ASAP7_75t_L g4281 ( 
.A1(n_4150),
.A2(n_4187),
.B(n_4195),
.Y(n_4281)
);

AND2x2_ASAP7_75t_L g4282 ( 
.A(n_4227),
.B(n_233),
.Y(n_4282)
);

BUFx3_ASAP7_75t_L g4283 ( 
.A(n_4146),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_4092),
.Y(n_4284)
);

HB1xp67_ASAP7_75t_L g4285 ( 
.A(n_4223),
.Y(n_4285)
);

AOI22xp5_ASAP7_75t_L g4286 ( 
.A1(n_4137),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.Y(n_4286)
);

NAND3xp33_ASAP7_75t_SL g4287 ( 
.A(n_4093),
.B(n_235),
.C(n_236),
.Y(n_4287)
);

INVxp67_ASAP7_75t_L g4288 ( 
.A(n_4142),
.Y(n_4288)
);

OAI221xp5_ASAP7_75t_L g4289 ( 
.A1(n_4239),
.A2(n_239),
.B1(n_237),
.B2(n_238),
.C(n_240),
.Y(n_4289)
);

NOR2xp33_ASAP7_75t_L g4290 ( 
.A(n_4120),
.B(n_4154),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4094),
.Y(n_4291)
);

NAND3xp33_ASAP7_75t_L g4292 ( 
.A(n_4133),
.B(n_239),
.C(n_240),
.Y(n_4292)
);

NAND2xp5_ASAP7_75t_L g4293 ( 
.A(n_4159),
.B(n_241),
.Y(n_4293)
);

NOR2xp33_ASAP7_75t_L g4294 ( 
.A(n_4120),
.B(n_241),
.Y(n_4294)
);

INVx3_ASAP7_75t_L g4295 ( 
.A(n_4216),
.Y(n_4295)
);

BUFx2_ASAP7_75t_L g4296 ( 
.A(n_4200),
.Y(n_4296)
);

AND2x2_ASAP7_75t_L g4297 ( 
.A(n_4201),
.B(n_242),
.Y(n_4297)
);

HB1xp67_ASAP7_75t_L g4298 ( 
.A(n_4132),
.Y(n_4298)
);

NOR2xp33_ASAP7_75t_L g4299 ( 
.A(n_4153),
.B(n_243),
.Y(n_4299)
);

INVx2_ASAP7_75t_L g4300 ( 
.A(n_4203),
.Y(n_4300)
);

NAND3xp33_ASAP7_75t_L g4301 ( 
.A(n_4191),
.B(n_243),
.C(n_244),
.Y(n_4301)
);

INVx2_ASAP7_75t_L g4302 ( 
.A(n_4206),
.Y(n_4302)
);

INVx1_ASAP7_75t_L g4303 ( 
.A(n_4098),
.Y(n_4303)
);

OAI221xp5_ASAP7_75t_L g4304 ( 
.A1(n_4186),
.A2(n_246),
.B1(n_244),
.B2(n_245),
.C(n_247),
.Y(n_4304)
);

BUFx2_ASAP7_75t_L g4305 ( 
.A(n_4213),
.Y(n_4305)
);

OAI211xp5_ASAP7_75t_L g4306 ( 
.A1(n_4198),
.A2(n_248),
.B(n_245),
.C(n_247),
.Y(n_4306)
);

INVx1_ASAP7_75t_L g4307 ( 
.A(n_4101),
.Y(n_4307)
);

OAI31xp33_ASAP7_75t_SL g4308 ( 
.A1(n_4134),
.A2(n_4188),
.A3(n_4189),
.B(n_4180),
.Y(n_4308)
);

INVx2_ASAP7_75t_L g4309 ( 
.A(n_4219),
.Y(n_4309)
);

INVx2_ASAP7_75t_L g4310 ( 
.A(n_4221),
.Y(n_4310)
);

NOR2x1_ASAP7_75t_L g4311 ( 
.A(n_4130),
.B(n_248),
.Y(n_4311)
);

INVx2_ASAP7_75t_SL g4312 ( 
.A(n_4088),
.Y(n_4312)
);

AOI222xp33_ASAP7_75t_SL g4313 ( 
.A1(n_4166),
.A2(n_251),
.B1(n_254),
.B2(n_249),
.C1(n_250),
.C2(n_253),
.Y(n_4313)
);

NAND4xp25_ASAP7_75t_L g4314 ( 
.A(n_4184),
.B(n_251),
.C(n_253),
.D(n_250),
.Y(n_4314)
);

AOI22xp33_ASAP7_75t_L g4315 ( 
.A1(n_4162),
.A2(n_256),
.B1(n_249),
.B2(n_255),
.Y(n_4315)
);

OAI22xp5_ASAP7_75t_L g4316 ( 
.A1(n_4168),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.Y(n_4316)
);

INVx4_ASAP7_75t_L g4317 ( 
.A(n_4130),
.Y(n_4317)
);

INVx2_ASAP7_75t_L g4318 ( 
.A(n_4238),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_4112),
.Y(n_4319)
);

NAND3xp33_ASAP7_75t_L g4320 ( 
.A(n_4185),
.B(n_257),
.C(n_258),
.Y(n_4320)
);

OAI22xp5_ASAP7_75t_L g4321 ( 
.A1(n_4232),
.A2(n_261),
.B1(n_258),
.B2(n_259),
.Y(n_4321)
);

OAI33xp33_ASAP7_75t_L g4322 ( 
.A1(n_4194),
.A2(n_263),
.A3(n_265),
.B1(n_259),
.B2(n_262),
.B3(n_264),
.Y(n_4322)
);

INVx2_ASAP7_75t_L g4323 ( 
.A(n_4085),
.Y(n_4323)
);

INVx5_ASAP7_75t_L g4324 ( 
.A(n_4139),
.Y(n_4324)
);

OAI33xp33_ASAP7_75t_L g4325 ( 
.A1(n_4087),
.A2(n_267),
.A3(n_269),
.B1(n_263),
.B2(n_266),
.B3(n_268),
.Y(n_4325)
);

OAI33xp33_ASAP7_75t_L g4326 ( 
.A1(n_4208),
.A2(n_271),
.A3(n_273),
.B1(n_268),
.B2(n_270),
.B3(n_272),
.Y(n_4326)
);

AOI22xp33_ASAP7_75t_SL g4327 ( 
.A1(n_4183),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.Y(n_4327)
);

HB1xp67_ASAP7_75t_L g4328 ( 
.A(n_4108),
.Y(n_4328)
);

OR2x2_ASAP7_75t_L g4329 ( 
.A(n_4212),
.B(n_274),
.Y(n_4329)
);

AND2x2_ASAP7_75t_L g4330 ( 
.A(n_4104),
.B(n_4106),
.Y(n_4330)
);

INVx2_ASAP7_75t_L g4331 ( 
.A(n_4204),
.Y(n_4331)
);

INVx2_ASAP7_75t_L g4332 ( 
.A(n_4230),
.Y(n_4332)
);

AND2x2_ASAP7_75t_L g4333 ( 
.A(n_4095),
.B(n_275),
.Y(n_4333)
);

AND2x4_ASAP7_75t_SL g4334 ( 
.A(n_4126),
.B(n_275),
.Y(n_4334)
);

AOI22xp33_ASAP7_75t_L g4335 ( 
.A1(n_4185),
.A2(n_279),
.B1(n_277),
.B2(n_278),
.Y(n_4335)
);

BUFx2_ASAP7_75t_L g4336 ( 
.A(n_4082),
.Y(n_4336)
);

AND2x4_ASAP7_75t_SL g4337 ( 
.A(n_4205),
.B(n_278),
.Y(n_4337)
);

AND2x2_ASAP7_75t_L g4338 ( 
.A(n_4210),
.B(n_279),
.Y(n_4338)
);

AOI22xp33_ASAP7_75t_SL g4339 ( 
.A1(n_4169),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_4339)
);

OAI22xp5_ASAP7_75t_L g4340 ( 
.A1(n_4151),
.A2(n_4218),
.B1(n_4229),
.B2(n_4217),
.Y(n_4340)
);

OR2x2_ASAP7_75t_L g4341 ( 
.A(n_4225),
.B(n_280),
.Y(n_4341)
);

AND2x2_ASAP7_75t_L g4342 ( 
.A(n_4211),
.B(n_282),
.Y(n_4342)
);

OAI22xp33_ASAP7_75t_L g4343 ( 
.A1(n_4197),
.A2(n_286),
.B1(n_283),
.B2(n_284),
.Y(n_4343)
);

AOI221xp5_ASAP7_75t_L g4344 ( 
.A1(n_4240),
.A2(n_287),
.B1(n_284),
.B2(n_286),
.C(n_288),
.Y(n_4344)
);

BUFx6f_ASAP7_75t_L g4345 ( 
.A(n_4143),
.Y(n_4345)
);

AND2x2_ASAP7_75t_L g4346 ( 
.A(n_4214),
.B(n_289),
.Y(n_4346)
);

NAND4xp25_ASAP7_75t_SL g4347 ( 
.A(n_4160),
.B(n_4176),
.C(n_4182),
.D(n_4145),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_SL g4348 ( 
.A(n_4148),
.B(n_290),
.Y(n_4348)
);

INVx2_ASAP7_75t_SL g4349 ( 
.A(n_4215),
.Y(n_4349)
);

OAI22xp33_ASAP7_75t_L g4350 ( 
.A1(n_4192),
.A2(n_292),
.B1(n_290),
.B2(n_291),
.Y(n_4350)
);

NAND2xp5_ASAP7_75t_L g4351 ( 
.A(n_4110),
.B(n_291),
.Y(n_4351)
);

INVx2_ASAP7_75t_L g4352 ( 
.A(n_4235),
.Y(n_4352)
);

NAND2xp5_ASAP7_75t_L g4353 ( 
.A(n_4107),
.B(n_292),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_SL g4354 ( 
.A(n_4097),
.B(n_4220),
.Y(n_4354)
);

INVx5_ASAP7_75t_L g4355 ( 
.A(n_4224),
.Y(n_4355)
);

AOI22xp33_ASAP7_75t_L g4356 ( 
.A1(n_4196),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_4356)
);

NAND3xp33_ASAP7_75t_L g4357 ( 
.A(n_4193),
.B(n_293),
.C(n_295),
.Y(n_4357)
);

OAI321xp33_ASAP7_75t_L g4358 ( 
.A1(n_4086),
.A2(n_299),
.A3(n_301),
.B1(n_296),
.B2(n_297),
.C(n_300),
.Y(n_4358)
);

AOI221xp5_ASAP7_75t_L g4359 ( 
.A1(n_4175),
.A2(n_301),
.B1(n_296),
.B2(n_299),
.C(n_302),
.Y(n_4359)
);

AND2x2_ASAP7_75t_L g4360 ( 
.A(n_4228),
.B(n_303),
.Y(n_4360)
);

AOI22xp33_ASAP7_75t_L g4361 ( 
.A1(n_4177),
.A2(n_305),
.B1(n_303),
.B2(n_304),
.Y(n_4361)
);

AOI21xp33_ASAP7_75t_L g4362 ( 
.A1(n_4149),
.A2(n_305),
.B(n_306),
.Y(n_4362)
);

AOI22xp33_ASAP7_75t_L g4363 ( 
.A1(n_4190),
.A2(n_310),
.B1(n_307),
.B2(n_308),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_4237),
.Y(n_4364)
);

AND2x2_ASAP7_75t_L g4365 ( 
.A(n_4233),
.B(n_4234),
.Y(n_4365)
);

AOI22xp33_ASAP7_75t_L g4366 ( 
.A1(n_4147),
.A2(n_312),
.B1(n_310),
.B2(n_311),
.Y(n_4366)
);

NAND2x1p5_ASAP7_75t_SL g4367 ( 
.A(n_4236),
.B(n_311),
.Y(n_4367)
);

OAI31xp33_ASAP7_75t_L g4368 ( 
.A1(n_4241),
.A2(n_315),
.A3(n_312),
.B(n_313),
.Y(n_4368)
);

INVx2_ASAP7_75t_L g4369 ( 
.A(n_4242),
.Y(n_4369)
);

INVx4_ASAP7_75t_L g4370 ( 
.A(n_4115),
.Y(n_4370)
);

AND2x4_ASAP7_75t_L g4371 ( 
.A(n_4105),
.B(n_313),
.Y(n_4371)
);

OAI211xp5_ASAP7_75t_L g4372 ( 
.A1(n_4099),
.A2(n_317),
.B(n_315),
.C(n_316),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_L g4373 ( 
.A(n_4102),
.B(n_317),
.Y(n_4373)
);

NAND2xp5_ASAP7_75t_SL g4374 ( 
.A(n_4118),
.B(n_318),
.Y(n_4374)
);

OAI211xp5_ASAP7_75t_SL g4375 ( 
.A1(n_4128),
.A2(n_321),
.B(n_319),
.C(n_320),
.Y(n_4375)
);

AND2x2_ASAP7_75t_L g4376 ( 
.A(n_4243),
.B(n_320),
.Y(n_4376)
);

OAI322xp33_ASAP7_75t_L g4377 ( 
.A1(n_4116),
.A2(n_327),
.A3(n_326),
.B1(n_324),
.B2(n_322),
.C1(n_323),
.C2(n_325),
.Y(n_4377)
);

OAI22xp33_ASAP7_75t_L g4378 ( 
.A1(n_4129),
.A2(n_4127),
.B1(n_4117),
.B2(n_4114),
.Y(n_4378)
);

AND2x2_ASAP7_75t_L g4379 ( 
.A(n_4111),
.B(n_322),
.Y(n_4379)
);

AOI221xp5_ASAP7_75t_L g4380 ( 
.A1(n_4165),
.A2(n_325),
.B1(n_323),
.B2(n_324),
.C(n_328),
.Y(n_4380)
);

INVx2_ASAP7_75t_SL g4381 ( 
.A(n_4146),
.Y(n_4381)
);

OAI321xp33_ASAP7_75t_L g4382 ( 
.A1(n_4165),
.A2(n_330),
.A3(n_334),
.B1(n_328),
.B2(n_329),
.C(n_333),
.Y(n_4382)
);

INVx2_ASAP7_75t_L g4383 ( 
.A(n_4131),
.Y(n_4383)
);

OR2x6_ASAP7_75t_L g4384 ( 
.A(n_4130),
.B(n_329),
.Y(n_4384)
);

NAND3xp33_ASAP7_75t_L g4385 ( 
.A(n_4222),
.B(n_333),
.C(n_335),
.Y(n_4385)
);

OAI21xp5_ASAP7_75t_L g4386 ( 
.A1(n_4165),
.A2(n_336),
.B(n_337),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_4083),
.Y(n_4387)
);

INVx2_ASAP7_75t_L g4388 ( 
.A(n_4131),
.Y(n_4388)
);

AOI21xp5_ASAP7_75t_L g4389 ( 
.A1(n_4171),
.A2(n_336),
.B(n_337),
.Y(n_4389)
);

INVx8_ASAP7_75t_L g4390 ( 
.A(n_4130),
.Y(n_4390)
);

BUFx6f_ASAP7_75t_L g4391 ( 
.A(n_4146),
.Y(n_4391)
);

AND2x2_ASAP7_75t_L g4392 ( 
.A(n_4135),
.B(n_338),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_4083),
.Y(n_4393)
);

OAI22xp5_ASAP7_75t_L g4394 ( 
.A1(n_4141),
.A2(n_340),
.B1(n_338),
.B2(n_339),
.Y(n_4394)
);

INVx2_ASAP7_75t_L g4395 ( 
.A(n_4131),
.Y(n_4395)
);

AOI22xp5_ASAP7_75t_L g4396 ( 
.A1(n_4165),
.A2(n_342),
.B1(n_339),
.B2(n_341),
.Y(n_4396)
);

OAI33xp33_ASAP7_75t_L g4397 ( 
.A1(n_4158),
.A2(n_345),
.A3(n_347),
.B1(n_341),
.B2(n_343),
.B3(n_346),
.Y(n_4397)
);

OAI21xp33_ASAP7_75t_L g4398 ( 
.A1(n_4141),
.A2(n_345),
.B(n_346),
.Y(n_4398)
);

NOR2xp33_ASAP7_75t_L g4399 ( 
.A(n_4140),
.B(n_348),
.Y(n_4399)
);

OAI211xp5_ASAP7_75t_L g4400 ( 
.A1(n_4141),
.A2(n_351),
.B(n_349),
.C(n_350),
.Y(n_4400)
);

NAND2xp5_ASAP7_75t_L g4401 ( 
.A(n_4141),
.B(n_350),
.Y(n_4401)
);

INVx2_ASAP7_75t_L g4402 ( 
.A(n_4131),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_4083),
.Y(n_4403)
);

NAND2xp5_ASAP7_75t_L g4404 ( 
.A(n_4141),
.B(n_351),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_4083),
.Y(n_4405)
);

OAI33xp33_ASAP7_75t_L g4406 ( 
.A1(n_4158),
.A2(n_355),
.A3(n_357),
.B1(n_352),
.B2(n_353),
.B3(n_356),
.Y(n_4406)
);

AOI221xp5_ASAP7_75t_L g4407 ( 
.A1(n_4165),
.A2(n_356),
.B1(n_352),
.B2(n_353),
.C(n_358),
.Y(n_4407)
);

INVx2_ASAP7_75t_L g4408 ( 
.A(n_4131),
.Y(n_4408)
);

AOI221xp5_ASAP7_75t_L g4409 ( 
.A1(n_4165),
.A2(n_361),
.B1(n_359),
.B2(n_360),
.C(n_362),
.Y(n_4409)
);

AND2x2_ASAP7_75t_L g4410 ( 
.A(n_4135),
.B(n_359),
.Y(n_4410)
);

AOI22xp33_ASAP7_75t_L g4411 ( 
.A1(n_4165),
.A2(n_364),
.B1(n_362),
.B2(n_363),
.Y(n_4411)
);

NAND3xp33_ASAP7_75t_L g4412 ( 
.A(n_4222),
.B(n_363),
.C(n_365),
.Y(n_4412)
);

NOR3xp33_ASAP7_75t_L g4413 ( 
.A(n_4165),
.B(n_366),
.C(n_367),
.Y(n_4413)
);

OAI221xp5_ASAP7_75t_L g4414 ( 
.A1(n_4165),
.A2(n_369),
.B1(n_367),
.B2(n_368),
.C(n_370),
.Y(n_4414)
);

AOI22xp33_ASAP7_75t_L g4415 ( 
.A1(n_4165),
.A2(n_373),
.B1(n_370),
.B2(n_371),
.Y(n_4415)
);

AOI21xp33_ASAP7_75t_L g4416 ( 
.A1(n_4113),
.A2(n_374),
.B(n_375),
.Y(n_4416)
);

INVx1_ASAP7_75t_L g4417 ( 
.A(n_4083),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_4083),
.Y(n_4418)
);

AOI22xp33_ASAP7_75t_L g4419 ( 
.A1(n_4165),
.A2(n_377),
.B1(n_375),
.B2(n_376),
.Y(n_4419)
);

AOI21xp5_ASAP7_75t_L g4420 ( 
.A1(n_4171),
.A2(n_376),
.B(n_377),
.Y(n_4420)
);

NAND2xp5_ASAP7_75t_L g4421 ( 
.A(n_4141),
.B(n_378),
.Y(n_4421)
);

INVx5_ASAP7_75t_SL g4422 ( 
.A(n_4130),
.Y(n_4422)
);

INVx4_ASAP7_75t_L g4423 ( 
.A(n_4130),
.Y(n_4423)
);

NAND2xp5_ASAP7_75t_L g4424 ( 
.A(n_4141),
.B(n_378),
.Y(n_4424)
);

INVx4_ASAP7_75t_R g4425 ( 
.A(n_4123),
.Y(n_4425)
);

AOI22xp33_ASAP7_75t_L g4426 ( 
.A1(n_4165),
.A2(n_382),
.B1(n_379),
.B2(n_381),
.Y(n_4426)
);

AOI22xp33_ASAP7_75t_L g4427 ( 
.A1(n_4165),
.A2(n_383),
.B1(n_379),
.B2(n_381),
.Y(n_4427)
);

AOI22xp33_ASAP7_75t_L g4428 ( 
.A1(n_4165),
.A2(n_385),
.B1(n_383),
.B2(n_384),
.Y(n_4428)
);

OR2x6_ASAP7_75t_L g4429 ( 
.A(n_4130),
.B(n_385),
.Y(n_4429)
);

OAI221xp5_ASAP7_75t_L g4430 ( 
.A1(n_4165),
.A2(n_388),
.B1(n_386),
.B2(n_387),
.C(n_389),
.Y(n_4430)
);

OR2x2_ASAP7_75t_L g4431 ( 
.A(n_4096),
.B(n_386),
.Y(n_4431)
);

INVx1_ASAP7_75t_L g4432 ( 
.A(n_4083),
.Y(n_4432)
);

OAI31xp33_ASAP7_75t_SL g4433 ( 
.A1(n_4113),
.A2(n_391),
.A3(n_393),
.B(n_390),
.Y(n_4433)
);

AND2x2_ASAP7_75t_L g4434 ( 
.A(n_4135),
.B(n_387),
.Y(n_4434)
);

OAI22xp5_ASAP7_75t_L g4435 ( 
.A1(n_4141),
.A2(n_394),
.B1(n_390),
.B2(n_391),
.Y(n_4435)
);

AND2x2_ASAP7_75t_L g4436 ( 
.A(n_4135),
.B(n_395),
.Y(n_4436)
);

AND2x2_ASAP7_75t_L g4437 ( 
.A(n_4135),
.B(n_395),
.Y(n_4437)
);

AOI221xp5_ASAP7_75t_L g4438 ( 
.A1(n_4165),
.A2(n_398),
.B1(n_396),
.B2(n_397),
.C(n_400),
.Y(n_4438)
);

INVx1_ASAP7_75t_L g4439 ( 
.A(n_4269),
.Y(n_4439)
);

INVxp67_ASAP7_75t_L g4440 ( 
.A(n_4336),
.Y(n_4440)
);

INVx2_ASAP7_75t_L g4441 ( 
.A(n_4283),
.Y(n_4441)
);

INVx1_ASAP7_75t_L g4442 ( 
.A(n_4298),
.Y(n_4442)
);

INVx2_ASAP7_75t_L g4443 ( 
.A(n_4391),
.Y(n_4443)
);

INVx3_ASAP7_75t_L g4444 ( 
.A(n_4391),
.Y(n_4444)
);

OR2x2_ASAP7_75t_L g4445 ( 
.A(n_4259),
.B(n_4279),
.Y(n_4445)
);

NAND2xp5_ASAP7_75t_L g4446 ( 
.A(n_4288),
.B(n_396),
.Y(n_4446)
);

OR2x2_ASAP7_75t_L g4447 ( 
.A(n_4349),
.B(n_400),
.Y(n_4447)
);

INVxp67_ASAP7_75t_SL g4448 ( 
.A(n_4285),
.Y(n_4448)
);

OR2x2_ASAP7_75t_L g4449 ( 
.A(n_4312),
.B(n_401),
.Y(n_4449)
);

NAND2xp5_ASAP7_75t_L g4450 ( 
.A(n_4355),
.B(n_401),
.Y(n_4450)
);

INVx1_ASAP7_75t_L g4451 ( 
.A(n_4328),
.Y(n_4451)
);

AND2x2_ASAP7_75t_L g4452 ( 
.A(n_4355),
.B(n_402),
.Y(n_4452)
);

NAND2xp5_ASAP7_75t_L g4453 ( 
.A(n_4355),
.B(n_4398),
.Y(n_4453)
);

INVx1_ASAP7_75t_L g4454 ( 
.A(n_4331),
.Y(n_4454)
);

INVx1_ASAP7_75t_L g4455 ( 
.A(n_4332),
.Y(n_4455)
);

INVx1_ASAP7_75t_L g4456 ( 
.A(n_4352),
.Y(n_4456)
);

INVx1_ASAP7_75t_L g4457 ( 
.A(n_4369),
.Y(n_4457)
);

INVx2_ASAP7_75t_L g4458 ( 
.A(n_4345),
.Y(n_4458)
);

NAND2xp5_ASAP7_75t_L g4459 ( 
.A(n_4324),
.B(n_402),
.Y(n_4459)
);

AND2x2_ASAP7_75t_L g4460 ( 
.A(n_4317),
.B(n_404),
.Y(n_4460)
);

AND2x2_ASAP7_75t_L g4461 ( 
.A(n_4423),
.B(n_404),
.Y(n_4461)
);

NAND2xp5_ASAP7_75t_SL g4462 ( 
.A(n_4324),
.B(n_405),
.Y(n_4462)
);

OR2x2_ASAP7_75t_L g4463 ( 
.A(n_4255),
.B(n_406),
.Y(n_4463)
);

NAND2xp5_ASAP7_75t_L g4464 ( 
.A(n_4324),
.B(n_406),
.Y(n_4464)
);

INVx2_ASAP7_75t_L g4465 ( 
.A(n_4345),
.Y(n_4465)
);

BUFx2_ASAP7_75t_L g4466 ( 
.A(n_4390),
.Y(n_4466)
);

AND2x2_ASAP7_75t_L g4467 ( 
.A(n_4381),
.B(n_407),
.Y(n_4467)
);

HB1xp67_ASAP7_75t_L g4468 ( 
.A(n_4263),
.Y(n_4468)
);

INVx2_ASAP7_75t_L g4469 ( 
.A(n_4390),
.Y(n_4469)
);

AND2x2_ASAP7_75t_L g4470 ( 
.A(n_4254),
.B(n_407),
.Y(n_4470)
);

INVx1_ASAP7_75t_L g4471 ( 
.A(n_4244),
.Y(n_4471)
);

INVx1_ASAP7_75t_L g4472 ( 
.A(n_4249),
.Y(n_4472)
);

INVx2_ASAP7_75t_L g4473 ( 
.A(n_4295),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_4256),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_4270),
.Y(n_4475)
);

INVx2_ASAP7_75t_L g4476 ( 
.A(n_4370),
.Y(n_4476)
);

AND2x2_ASAP7_75t_L g4477 ( 
.A(n_4261),
.B(n_409),
.Y(n_4477)
);

INVx2_ASAP7_75t_L g4478 ( 
.A(n_4296),
.Y(n_4478)
);

AND2x2_ASAP7_75t_L g4479 ( 
.A(n_4305),
.B(n_409),
.Y(n_4479)
);

INVx2_ASAP7_75t_L g4480 ( 
.A(n_4422),
.Y(n_4480)
);

INVx2_ASAP7_75t_L g4481 ( 
.A(n_4422),
.Y(n_4481)
);

NAND2xp5_ASAP7_75t_L g4482 ( 
.A(n_4308),
.B(n_410),
.Y(n_4482)
);

AND2x2_ASAP7_75t_L g4483 ( 
.A(n_4365),
.B(n_410),
.Y(n_4483)
);

HB1xp67_ASAP7_75t_SL g4484 ( 
.A(n_4290),
.Y(n_4484)
);

BUFx2_ASAP7_75t_L g4485 ( 
.A(n_4384),
.Y(n_4485)
);

AND2x4_ASAP7_75t_L g4486 ( 
.A(n_4330),
.B(n_4245),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_4284),
.Y(n_4487)
);

AND2x2_ASAP7_75t_L g4488 ( 
.A(n_4383),
.B(n_411),
.Y(n_4488)
);

AND2x2_ASAP7_75t_L g4489 ( 
.A(n_4388),
.B(n_411),
.Y(n_4489)
);

INVx1_ASAP7_75t_L g4490 ( 
.A(n_4291),
.Y(n_4490)
);

AOI22xp33_ASAP7_75t_L g4491 ( 
.A1(n_4275),
.A2(n_414),
.B1(n_412),
.B2(n_413),
.Y(n_4491)
);

INVx2_ASAP7_75t_L g4492 ( 
.A(n_4300),
.Y(n_4492)
);

AND2x2_ASAP7_75t_L g4493 ( 
.A(n_4395),
.B(n_412),
.Y(n_4493)
);

AND2x2_ASAP7_75t_L g4494 ( 
.A(n_4402),
.B(n_413),
.Y(n_4494)
);

OR2x2_ASAP7_75t_L g4495 ( 
.A(n_4408),
.B(n_414),
.Y(n_4495)
);

INVx2_ASAP7_75t_L g4496 ( 
.A(n_4302),
.Y(n_4496)
);

NAND2xp5_ASAP7_75t_L g4497 ( 
.A(n_4246),
.B(n_415),
.Y(n_4497)
);

INVx2_ASAP7_75t_L g4498 ( 
.A(n_4309),
.Y(n_4498)
);

AND2x2_ASAP7_75t_L g4499 ( 
.A(n_4310),
.B(n_415),
.Y(n_4499)
);

AND2x4_ASAP7_75t_L g4500 ( 
.A(n_4297),
.B(n_416),
.Y(n_4500)
);

NAND2xp5_ASAP7_75t_L g4501 ( 
.A(n_4378),
.B(n_416),
.Y(n_4501)
);

OAI221xp5_ASAP7_75t_SL g4502 ( 
.A1(n_4433),
.A2(n_420),
.B1(n_417),
.B2(n_418),
.C(n_421),
.Y(n_4502)
);

INVx2_ASAP7_75t_L g4503 ( 
.A(n_4318),
.Y(n_4503)
);

AND2x2_ASAP7_75t_L g4504 ( 
.A(n_4251),
.B(n_417),
.Y(n_4504)
);

OR2x2_ASAP7_75t_L g4505 ( 
.A(n_4323),
.B(n_418),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4303),
.Y(n_4506)
);

AND2x2_ASAP7_75t_L g4507 ( 
.A(n_4247),
.B(n_420),
.Y(n_4507)
);

AND2x2_ASAP7_75t_L g4508 ( 
.A(n_4392),
.B(n_4410),
.Y(n_4508)
);

AND2x4_ASAP7_75t_L g4509 ( 
.A(n_4311),
.B(n_421),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_4307),
.Y(n_4510)
);

NAND2xp5_ASAP7_75t_L g4511 ( 
.A(n_4401),
.B(n_4404),
.Y(n_4511)
);

AND2x2_ASAP7_75t_L g4512 ( 
.A(n_4434),
.B(n_422),
.Y(n_4512)
);

AOI22xp5_ASAP7_75t_L g4513 ( 
.A1(n_4313),
.A2(n_425),
.B1(n_423),
.B2(n_424),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4319),
.Y(n_4514)
);

AND2x4_ASAP7_75t_L g4515 ( 
.A(n_4267),
.B(n_423),
.Y(n_4515)
);

INVx1_ASAP7_75t_L g4516 ( 
.A(n_4364),
.Y(n_4516)
);

INVx1_ASAP7_75t_L g4517 ( 
.A(n_4387),
.Y(n_4517)
);

INVx3_ASAP7_75t_L g4518 ( 
.A(n_4334),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_L g4519 ( 
.A(n_4421),
.B(n_424),
.Y(n_4519)
);

OR2x2_ASAP7_75t_L g4520 ( 
.A(n_4424),
.B(n_4340),
.Y(n_4520)
);

NAND2x1p5_ASAP7_75t_L g4521 ( 
.A(n_4252),
.B(n_4282),
.Y(n_4521)
);

AND2x2_ASAP7_75t_L g4522 ( 
.A(n_4436),
.B(n_425),
.Y(n_4522)
);

OR2x2_ASAP7_75t_L g4523 ( 
.A(n_4274),
.B(n_426),
.Y(n_4523)
);

OR2x2_ASAP7_75t_L g4524 ( 
.A(n_4293),
.B(n_4354),
.Y(n_4524)
);

OR2x6_ASAP7_75t_L g4525 ( 
.A(n_4384),
.B(n_426),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_4393),
.Y(n_4526)
);

BUFx4f_ASAP7_75t_SL g4527 ( 
.A(n_4371),
.Y(n_4527)
);

HB1xp67_ASAP7_75t_L g4528 ( 
.A(n_4431),
.Y(n_4528)
);

AND2x2_ASAP7_75t_L g4529 ( 
.A(n_4437),
.B(n_427),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_L g4530 ( 
.A(n_4394),
.B(n_428),
.Y(n_4530)
);

INVx2_ASAP7_75t_L g4531 ( 
.A(n_4253),
.Y(n_4531)
);

AND2x2_ASAP7_75t_L g4532 ( 
.A(n_4338),
.B(n_428),
.Y(n_4532)
);

AND2x2_ASAP7_75t_L g4533 ( 
.A(n_4342),
.B(n_429),
.Y(n_4533)
);

NAND2xp5_ASAP7_75t_L g4534 ( 
.A(n_4435),
.B(n_429),
.Y(n_4534)
);

AND2x2_ASAP7_75t_L g4535 ( 
.A(n_4346),
.B(n_430),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_4403),
.Y(n_4536)
);

AND2x2_ASAP7_75t_L g4537 ( 
.A(n_4360),
.B(n_430),
.Y(n_4537)
);

NAND2xp5_ASAP7_75t_SL g4538 ( 
.A(n_4271),
.B(n_431),
.Y(n_4538)
);

INVx1_ASAP7_75t_L g4539 ( 
.A(n_4405),
.Y(n_4539)
);

INVx2_ASAP7_75t_L g4540 ( 
.A(n_4376),
.Y(n_4540)
);

AND2x2_ASAP7_75t_L g4541 ( 
.A(n_4333),
.B(n_431),
.Y(n_4541)
);

INVx2_ASAP7_75t_L g4542 ( 
.A(n_4417),
.Y(n_4542)
);

INVx2_ASAP7_75t_L g4543 ( 
.A(n_4418),
.Y(n_4543)
);

AND2x2_ASAP7_75t_L g4544 ( 
.A(n_4379),
.B(n_432),
.Y(n_4544)
);

INVx3_ASAP7_75t_L g4545 ( 
.A(n_4337),
.Y(n_4545)
);

INVx2_ASAP7_75t_SL g4546 ( 
.A(n_4280),
.Y(n_4546)
);

INVxp67_ASAP7_75t_L g4547 ( 
.A(n_4399),
.Y(n_4547)
);

INVx1_ASAP7_75t_SL g4548 ( 
.A(n_4429),
.Y(n_4548)
);

AND2x2_ASAP7_75t_L g4549 ( 
.A(n_4299),
.B(n_432),
.Y(n_4549)
);

INVx1_ASAP7_75t_L g4550 ( 
.A(n_4432),
.Y(n_4550)
);

OR2x2_ASAP7_75t_L g4551 ( 
.A(n_4367),
.B(n_433),
.Y(n_4551)
);

INVx1_ASAP7_75t_L g4552 ( 
.A(n_4373),
.Y(n_4552)
);

INVx1_ASAP7_75t_L g4553 ( 
.A(n_4329),
.Y(n_4553)
);

BUFx3_ASAP7_75t_L g4554 ( 
.A(n_4429),
.Y(n_4554)
);

NAND2x1p5_ASAP7_75t_L g4555 ( 
.A(n_4348),
.B(n_433),
.Y(n_4555)
);

HB1xp67_ASAP7_75t_L g4556 ( 
.A(n_4347),
.Y(n_4556)
);

INVx1_ASAP7_75t_L g4557 ( 
.A(n_4341),
.Y(n_4557)
);

INVxp67_ASAP7_75t_L g4558 ( 
.A(n_4272),
.Y(n_4558)
);

HB1xp67_ASAP7_75t_L g4559 ( 
.A(n_4374),
.Y(n_4559)
);

INVx2_ASAP7_75t_L g4560 ( 
.A(n_4351),
.Y(n_4560)
);

NAND2xp5_ASAP7_75t_L g4561 ( 
.A(n_4389),
.B(n_434),
.Y(n_4561)
);

INVx2_ASAP7_75t_L g4562 ( 
.A(n_4353),
.Y(n_4562)
);

AND2x2_ASAP7_75t_L g4563 ( 
.A(n_4281),
.B(n_434),
.Y(n_4563)
);

NAND2xp5_ASAP7_75t_L g4564 ( 
.A(n_4420),
.B(n_435),
.Y(n_4564)
);

OR2x2_ASAP7_75t_L g4565 ( 
.A(n_4292),
.B(n_435),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_4400),
.Y(n_4566)
);

INVx1_ASAP7_75t_L g4567 ( 
.A(n_4301),
.Y(n_4567)
);

INVx2_ASAP7_75t_L g4568 ( 
.A(n_4294),
.Y(n_4568)
);

INVx2_ASAP7_75t_L g4569 ( 
.A(n_4320),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_4316),
.Y(n_4570)
);

INVx1_ASAP7_75t_L g4571 ( 
.A(n_4357),
.Y(n_4571)
);

AND2x2_ASAP7_75t_L g4572 ( 
.A(n_4386),
.B(n_436),
.Y(n_4572)
);

INVx1_ASAP7_75t_L g4573 ( 
.A(n_4258),
.Y(n_4573)
);

INVx2_ASAP7_75t_L g4574 ( 
.A(n_4277),
.Y(n_4574)
);

HB1xp67_ASAP7_75t_L g4575 ( 
.A(n_4321),
.Y(n_4575)
);

NAND3xp33_ASAP7_75t_L g4576 ( 
.A(n_4558),
.B(n_4413),
.C(n_4268),
.Y(n_4576)
);

INVx1_ASAP7_75t_L g4577 ( 
.A(n_4439),
.Y(n_4577)
);

NOR3xp33_ASAP7_75t_L g4578 ( 
.A(n_4466),
.B(n_4385),
.C(n_4257),
.Y(n_4578)
);

AOI22xp33_ASAP7_75t_L g4579 ( 
.A1(n_4556),
.A2(n_4412),
.B1(n_4287),
.B2(n_4314),
.Y(n_4579)
);

INVx2_ASAP7_75t_L g4580 ( 
.A(n_4546),
.Y(n_4580)
);

NAND2xp5_ASAP7_75t_L g4581 ( 
.A(n_4548),
.B(n_4339),
.Y(n_4581)
);

INVx2_ASAP7_75t_L g4582 ( 
.A(n_4545),
.Y(n_4582)
);

INVx1_ASAP7_75t_L g4583 ( 
.A(n_4528),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_4448),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4505),
.Y(n_4585)
);

AOI211xp5_ASAP7_75t_SL g4586 ( 
.A1(n_4502),
.A2(n_4382),
.B(n_4358),
.C(n_4306),
.Y(n_4586)
);

HB1xp67_ASAP7_75t_L g4587 ( 
.A(n_4485),
.Y(n_4587)
);

OAI33xp33_ASAP7_75t_L g4588 ( 
.A1(n_4520),
.A2(n_4350),
.A3(n_4343),
.B1(n_4276),
.B2(n_4248),
.B3(n_4264),
.Y(n_4588)
);

NAND2xp5_ASAP7_75t_L g4589 ( 
.A(n_4566),
.B(n_4396),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_4495),
.Y(n_4590)
);

AND2x2_ASAP7_75t_L g4591 ( 
.A(n_4480),
.B(n_4425),
.Y(n_4591)
);

OR2x2_ASAP7_75t_L g4592 ( 
.A(n_4511),
.B(n_4372),
.Y(n_4592)
);

NAND2xp5_ASAP7_75t_L g4593 ( 
.A(n_4508),
.B(n_4368),
.Y(n_4593)
);

AND2x2_ASAP7_75t_L g4594 ( 
.A(n_4481),
.B(n_4362),
.Y(n_4594)
);

NAND2xp5_ASAP7_75t_L g4595 ( 
.A(n_4554),
.B(n_4327),
.Y(n_4595)
);

INVx3_ASAP7_75t_L g4596 ( 
.A(n_4518),
.Y(n_4596)
);

NAND2xp5_ASAP7_75t_L g4597 ( 
.A(n_4478),
.B(n_4344),
.Y(n_4597)
);

AND2x2_ASAP7_75t_L g4598 ( 
.A(n_4469),
.B(n_4273),
.Y(n_4598)
);

AND2x2_ASAP7_75t_L g4599 ( 
.A(n_4441),
.B(n_4315),
.Y(n_4599)
);

INVx1_ASAP7_75t_L g4600 ( 
.A(n_4447),
.Y(n_4600)
);

INVx1_ASAP7_75t_L g4601 ( 
.A(n_4449),
.Y(n_4601)
);

INVx2_ASAP7_75t_L g4602 ( 
.A(n_4527),
.Y(n_4602)
);

INVxp67_ASAP7_75t_SL g4603 ( 
.A(n_4484),
.Y(n_4603)
);

AND2x2_ASAP7_75t_L g4604 ( 
.A(n_4444),
.B(n_4278),
.Y(n_4604)
);

OAI21xp5_ASAP7_75t_L g4605 ( 
.A1(n_4482),
.A2(n_4491),
.B(n_4521),
.Y(n_4605)
);

NOR2xp33_ASAP7_75t_L g4606 ( 
.A(n_4547),
.B(n_4260),
.Y(n_4606)
);

OR2x2_ASAP7_75t_L g4607 ( 
.A(n_4440),
.B(n_4416),
.Y(n_4607)
);

OAI221xp5_ASAP7_75t_L g4608 ( 
.A1(n_4453),
.A2(n_4359),
.B1(n_4409),
.B2(n_4407),
.C(n_4380),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_4442),
.Y(n_4609)
);

BUFx2_ASAP7_75t_L g4610 ( 
.A(n_4452),
.Y(n_4610)
);

AND2x2_ASAP7_75t_L g4611 ( 
.A(n_4443),
.B(n_4335),
.Y(n_4611)
);

INVx2_ASAP7_75t_L g4612 ( 
.A(n_4458),
.Y(n_4612)
);

OAI33xp33_ASAP7_75t_L g4613 ( 
.A1(n_4451),
.A2(n_4375),
.A3(n_4262),
.B1(n_4397),
.B2(n_4406),
.B3(n_4322),
.Y(n_4613)
);

INVx1_ASAP7_75t_L g4614 ( 
.A(n_4553),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_4557),
.Y(n_4615)
);

NAND2xp5_ASAP7_75t_L g4616 ( 
.A(n_4468),
.B(n_4438),
.Y(n_4616)
);

NAND2x1_ASAP7_75t_SL g4617 ( 
.A(n_4509),
.B(n_4559),
.Y(n_4617)
);

HB1xp67_ASAP7_75t_L g4618 ( 
.A(n_4459),
.Y(n_4618)
);

INVx4_ASAP7_75t_L g4619 ( 
.A(n_4525),
.Y(n_4619)
);

AO21x2_ASAP7_75t_L g4620 ( 
.A1(n_4464),
.A2(n_4430),
.B(n_4414),
.Y(n_4620)
);

NOR3xp33_ASAP7_75t_L g4621 ( 
.A(n_4476),
.B(n_4265),
.C(n_4266),
.Y(n_4621)
);

INVx1_ASAP7_75t_SL g4622 ( 
.A(n_4525),
.Y(n_4622)
);

INVx1_ASAP7_75t_L g4623 ( 
.A(n_4454),
.Y(n_4623)
);

AOI22xp33_ASAP7_75t_SL g4624 ( 
.A1(n_4575),
.A2(n_4289),
.B1(n_4304),
.B2(n_4325),
.Y(n_4624)
);

NAND2xp5_ASAP7_75t_L g4625 ( 
.A(n_4486),
.B(n_4366),
.Y(n_4625)
);

OR2x2_ASAP7_75t_L g4626 ( 
.A(n_4445),
.B(n_4363),
.Y(n_4626)
);

INVx1_ASAP7_75t_L g4627 ( 
.A(n_4455),
.Y(n_4627)
);

OAI31xp33_ASAP7_75t_L g4628 ( 
.A1(n_4573),
.A2(n_4411),
.A3(n_4415),
.B(n_4250),
.Y(n_4628)
);

BUFx2_ASAP7_75t_L g4629 ( 
.A(n_4479),
.Y(n_4629)
);

INVx2_ASAP7_75t_SL g4630 ( 
.A(n_4467),
.Y(n_4630)
);

INVxp67_ASAP7_75t_L g4631 ( 
.A(n_4462),
.Y(n_4631)
);

AND2x2_ASAP7_75t_SL g4632 ( 
.A(n_4551),
.B(n_4419),
.Y(n_4632)
);

NAND2xp5_ASAP7_75t_L g4633 ( 
.A(n_4568),
.B(n_4426),
.Y(n_4633)
);

INVx2_ASAP7_75t_L g4634 ( 
.A(n_4465),
.Y(n_4634)
);

INVx1_ASAP7_75t_L g4635 ( 
.A(n_4456),
.Y(n_4635)
);

AND2x4_ASAP7_75t_L g4636 ( 
.A(n_4473),
.B(n_4286),
.Y(n_4636)
);

AOI22xp33_ASAP7_75t_SL g4637 ( 
.A1(n_4567),
.A2(n_4326),
.B1(n_4377),
.B2(n_4427),
.Y(n_4637)
);

AND2x2_ASAP7_75t_L g4638 ( 
.A(n_4540),
.B(n_4428),
.Y(n_4638)
);

INVx1_ASAP7_75t_L g4639 ( 
.A(n_4457),
.Y(n_4639)
);

AOI33xp33_ASAP7_75t_L g4640 ( 
.A1(n_4513),
.A2(n_4571),
.A3(n_4570),
.B1(n_4574),
.B2(n_4569),
.B3(n_4563),
.Y(n_4640)
);

AOI33xp33_ASAP7_75t_L g4641 ( 
.A1(n_4552),
.A2(n_4356),
.A3(n_4361),
.B1(n_438),
.B2(n_440),
.B3(n_436),
.Y(n_4641)
);

AOI211xp5_ASAP7_75t_SL g4642 ( 
.A1(n_4565),
.A2(n_439),
.B(n_437),
.C(n_438),
.Y(n_4642)
);

INVx3_ASAP7_75t_L g4643 ( 
.A(n_4500),
.Y(n_4643)
);

OAI21xp33_ASAP7_75t_L g4644 ( 
.A1(n_4524),
.A2(n_4562),
.B(n_4560),
.Y(n_4644)
);

NAND3xp33_ASAP7_75t_L g4645 ( 
.A(n_4538),
.B(n_442),
.C(n_439),
.Y(n_4645)
);

NOR2xp33_ASAP7_75t_L g4646 ( 
.A(n_4463),
.B(n_437),
.Y(n_4646)
);

INVx1_ASAP7_75t_L g4647 ( 
.A(n_4542),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4543),
.Y(n_4648)
);

AND2x2_ASAP7_75t_L g4649 ( 
.A(n_4531),
.B(n_442),
.Y(n_4649)
);

INVx2_ASAP7_75t_L g4650 ( 
.A(n_4460),
.Y(n_4650)
);

OAI21xp5_ASAP7_75t_SL g4651 ( 
.A1(n_4501),
.A2(n_443),
.B(n_444),
.Y(n_4651)
);

AND2x2_ASAP7_75t_L g4652 ( 
.A(n_4461),
.B(n_445),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_4471),
.Y(n_4653)
);

OAI221xp5_ASAP7_75t_SL g4654 ( 
.A1(n_4497),
.A2(n_448),
.B1(n_446),
.B2(n_447),
.C(n_449),
.Y(n_4654)
);

NAND2xp5_ASAP7_75t_SL g4655 ( 
.A(n_4555),
.B(n_446),
.Y(n_4655)
);

NOR2xp33_ASAP7_75t_R g4656 ( 
.A(n_4504),
.B(n_447),
.Y(n_4656)
);

INVx2_ASAP7_75t_SL g4657 ( 
.A(n_4470),
.Y(n_4657)
);

A2O1A1Ixp33_ASAP7_75t_SL g4658 ( 
.A1(n_4561),
.A2(n_451),
.B(n_448),
.C(n_450),
.Y(n_4658)
);

HB1xp67_ASAP7_75t_L g4659 ( 
.A(n_4450),
.Y(n_4659)
);

INVx2_ASAP7_75t_L g4660 ( 
.A(n_4499),
.Y(n_4660)
);

AND2x2_ASAP7_75t_L g4661 ( 
.A(n_4483),
.B(n_450),
.Y(n_4661)
);

NAND3xp33_ASAP7_75t_L g4662 ( 
.A(n_4492),
.B(n_454),
.C(n_453),
.Y(n_4662)
);

AND2x2_ASAP7_75t_L g4663 ( 
.A(n_4496),
.B(n_452),
.Y(n_4663)
);

INVx2_ASAP7_75t_SL g4664 ( 
.A(n_4477),
.Y(n_4664)
);

OR2x2_ASAP7_75t_L g4665 ( 
.A(n_4498),
.B(n_453),
.Y(n_4665)
);

NAND3xp33_ASAP7_75t_L g4666 ( 
.A(n_4503),
.B(n_458),
.C(n_456),
.Y(n_4666)
);

AOI22xp5_ASAP7_75t_L g4667 ( 
.A1(n_4572),
.A2(n_459),
.B1(n_455),
.B2(n_456),
.Y(n_4667)
);

AND3x1_ASAP7_75t_L g4668 ( 
.A(n_4446),
.B(n_455),
.C(n_459),
.Y(n_4668)
);

AND2x2_ASAP7_75t_L g4669 ( 
.A(n_4591),
.B(n_4515),
.Y(n_4669)
);

AND2x2_ASAP7_75t_L g4670 ( 
.A(n_4603),
.B(n_4507),
.Y(n_4670)
);

INVx1_ASAP7_75t_L g4671 ( 
.A(n_4587),
.Y(n_4671)
);

AND2x2_ASAP7_75t_L g4672 ( 
.A(n_4596),
.B(n_4512),
.Y(n_4672)
);

NOR2xp33_ASAP7_75t_L g4673 ( 
.A(n_4619),
.B(n_4602),
.Y(n_4673)
);

OR2x2_ASAP7_75t_L g4674 ( 
.A(n_4610),
.B(n_4564),
.Y(n_4674)
);

NOR2xp33_ASAP7_75t_L g4675 ( 
.A(n_4622),
.B(n_4519),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_4584),
.Y(n_4676)
);

INVx2_ASAP7_75t_L g4677 ( 
.A(n_4580),
.Y(n_4677)
);

INVx2_ASAP7_75t_L g4678 ( 
.A(n_4582),
.Y(n_4678)
);

NAND2x1p5_ASAP7_75t_L g4679 ( 
.A(n_4668),
.B(n_4488),
.Y(n_4679)
);

AND2x2_ASAP7_75t_L g4680 ( 
.A(n_4629),
.B(n_4643),
.Y(n_4680)
);

AND2x2_ASAP7_75t_L g4681 ( 
.A(n_4650),
.B(n_4522),
.Y(n_4681)
);

NAND2xp5_ASAP7_75t_SL g4682 ( 
.A(n_4631),
.B(n_4530),
.Y(n_4682)
);

AND2x4_ASAP7_75t_L g4683 ( 
.A(n_4630),
.B(n_4489),
.Y(n_4683)
);

NOR2x1_ASAP7_75t_L g4684 ( 
.A(n_4662),
.B(n_4534),
.Y(n_4684)
);

INVx2_ASAP7_75t_L g4685 ( 
.A(n_4617),
.Y(n_4685)
);

INVx2_ASAP7_75t_L g4686 ( 
.A(n_4657),
.Y(n_4686)
);

HB1xp67_ASAP7_75t_L g4687 ( 
.A(n_4656),
.Y(n_4687)
);

NAND2xp5_ASAP7_75t_L g4688 ( 
.A(n_4586),
.B(n_4493),
.Y(n_4688)
);

AND2x2_ASAP7_75t_L g4689 ( 
.A(n_4604),
.B(n_4529),
.Y(n_4689)
);

INVx1_ASAP7_75t_L g4690 ( 
.A(n_4649),
.Y(n_4690)
);

AND2x2_ASAP7_75t_L g4691 ( 
.A(n_4598),
.B(n_4532),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4665),
.Y(n_4692)
);

OR2x2_ASAP7_75t_L g4693 ( 
.A(n_4581),
.B(n_4595),
.Y(n_4693)
);

AND2x2_ASAP7_75t_L g4694 ( 
.A(n_4594),
.B(n_4533),
.Y(n_4694)
);

NAND2xp5_ASAP7_75t_L g4695 ( 
.A(n_4632),
.B(n_4640),
.Y(n_4695)
);

NAND2xp5_ASAP7_75t_L g4696 ( 
.A(n_4637),
.B(n_4494),
.Y(n_4696)
);

INVx1_ASAP7_75t_L g4697 ( 
.A(n_4583),
.Y(n_4697)
);

INVx2_ASAP7_75t_L g4698 ( 
.A(n_4664),
.Y(n_4698)
);

AND2x2_ASAP7_75t_L g4699 ( 
.A(n_4636),
.B(n_4599),
.Y(n_4699)
);

AND2x2_ASAP7_75t_L g4700 ( 
.A(n_4636),
.B(n_4535),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_4663),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4600),
.Y(n_4702)
);

AOI21xp5_ASAP7_75t_L g4703 ( 
.A1(n_4616),
.A2(n_4523),
.B(n_4549),
.Y(n_4703)
);

BUFx2_ASAP7_75t_L g4704 ( 
.A(n_4601),
.Y(n_4704)
);

INVx1_ASAP7_75t_L g4705 ( 
.A(n_4585),
.Y(n_4705)
);

INVx1_ASAP7_75t_L g4706 ( 
.A(n_4590),
.Y(n_4706)
);

HB1xp67_ASAP7_75t_L g4707 ( 
.A(n_4618),
.Y(n_4707)
);

NOR2x1_ASAP7_75t_L g4708 ( 
.A(n_4666),
.B(n_4537),
.Y(n_4708)
);

AOI22xp5_ASAP7_75t_L g4709 ( 
.A1(n_4576),
.A2(n_4517),
.B1(n_4526),
.B2(n_4516),
.Y(n_4709)
);

NOR2xp33_ASAP7_75t_L g4710 ( 
.A(n_4588),
.B(n_4541),
.Y(n_4710)
);

NOR2x1p5_ASAP7_75t_L g4711 ( 
.A(n_4625),
.B(n_4593),
.Y(n_4711)
);

INVx1_ASAP7_75t_SL g4712 ( 
.A(n_4652),
.Y(n_4712)
);

AND2x4_ASAP7_75t_L g4713 ( 
.A(n_4612),
.B(n_4544),
.Y(n_4713)
);

INVx1_ASAP7_75t_L g4714 ( 
.A(n_4659),
.Y(n_4714)
);

AOI21xp33_ASAP7_75t_L g4715 ( 
.A1(n_4605),
.A2(n_4474),
.B(n_4472),
.Y(n_4715)
);

AND2x2_ASAP7_75t_L g4716 ( 
.A(n_4611),
.B(n_4475),
.Y(n_4716)
);

NAND2xp5_ASAP7_75t_L g4717 ( 
.A(n_4624),
.B(n_4487),
.Y(n_4717)
);

OR2x2_ASAP7_75t_L g4718 ( 
.A(n_4592),
.B(n_4490),
.Y(n_4718)
);

INVx1_ASAP7_75t_L g4719 ( 
.A(n_4577),
.Y(n_4719)
);

NOR2xp33_ASAP7_75t_L g4720 ( 
.A(n_4651),
.B(n_4506),
.Y(n_4720)
);

NOR2x1_ASAP7_75t_L g4721 ( 
.A(n_4645),
.B(n_4510),
.Y(n_4721)
);

INVx1_ASAP7_75t_L g4722 ( 
.A(n_4609),
.Y(n_4722)
);

INVx1_ASAP7_75t_L g4723 ( 
.A(n_4614),
.Y(n_4723)
);

INVx1_ASAP7_75t_L g4724 ( 
.A(n_4615),
.Y(n_4724)
);

AND2x2_ASAP7_75t_L g4725 ( 
.A(n_4634),
.B(n_4514),
.Y(n_4725)
);

OR2x2_ASAP7_75t_L g4726 ( 
.A(n_4589),
.B(n_4536),
.Y(n_4726)
);

HB1xp67_ASAP7_75t_L g4727 ( 
.A(n_4660),
.Y(n_4727)
);

INVx1_ASAP7_75t_L g4728 ( 
.A(n_4647),
.Y(n_4728)
);

OA21x2_ASAP7_75t_L g4729 ( 
.A1(n_4579),
.A2(n_4550),
.B(n_4539),
.Y(n_4729)
);

AND2x4_ASAP7_75t_L g4730 ( 
.A(n_4680),
.B(n_4578),
.Y(n_4730)
);

OR2x2_ASAP7_75t_L g4731 ( 
.A(n_4687),
.B(n_4607),
.Y(n_4731)
);

NOR2x1_ASAP7_75t_L g4732 ( 
.A(n_4671),
.B(n_4655),
.Y(n_4732)
);

AOI221xp5_ASAP7_75t_L g4733 ( 
.A1(n_4715),
.A2(n_4608),
.B1(n_4613),
.B2(n_4597),
.C(n_4644),
.Y(n_4733)
);

AOI22xp5_ASAP7_75t_L g4734 ( 
.A1(n_4695),
.A2(n_4621),
.B1(n_4717),
.B2(n_4620),
.Y(n_4734)
);

INVx1_ASAP7_75t_SL g4735 ( 
.A(n_4699),
.Y(n_4735)
);

INVx1_ASAP7_75t_L g4736 ( 
.A(n_4707),
.Y(n_4736)
);

AND2x2_ASAP7_75t_L g4737 ( 
.A(n_4670),
.B(n_4638),
.Y(n_4737)
);

NAND2xp5_ASAP7_75t_L g4738 ( 
.A(n_4700),
.B(n_4642),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4704),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_4727),
.Y(n_4740)
);

OR2x2_ASAP7_75t_L g4741 ( 
.A(n_4712),
.B(n_4626),
.Y(n_4741)
);

AND2x2_ASAP7_75t_L g4742 ( 
.A(n_4669),
.B(n_4661),
.Y(n_4742)
);

NOR2xp33_ASAP7_75t_L g4743 ( 
.A(n_4679),
.B(n_4606),
.Y(n_4743)
);

NAND3xp33_ASAP7_75t_L g4744 ( 
.A(n_4710),
.B(n_4628),
.C(n_4633),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_L g4745 ( 
.A(n_4672),
.B(n_4646),
.Y(n_4745)
);

NAND2xp5_ASAP7_75t_L g4746 ( 
.A(n_4689),
.B(n_4648),
.Y(n_4746)
);

AND2x2_ASAP7_75t_L g4747 ( 
.A(n_4691),
.B(n_4623),
.Y(n_4747)
);

AND2x2_ASAP7_75t_L g4748 ( 
.A(n_4685),
.B(n_4627),
.Y(n_4748)
);

AND2x2_ASAP7_75t_L g4749 ( 
.A(n_4694),
.B(n_4681),
.Y(n_4749)
);

OAI21xp33_ASAP7_75t_L g4750 ( 
.A1(n_4673),
.A2(n_4639),
.B(n_4635),
.Y(n_4750)
);

INVx1_ASAP7_75t_L g4751 ( 
.A(n_4686),
.Y(n_4751)
);

CKINVDCx5p33_ASAP7_75t_R g4752 ( 
.A(n_4675),
.Y(n_4752)
);

INVx2_ASAP7_75t_L g4753 ( 
.A(n_4713),
.Y(n_4753)
);

NAND3xp33_ASAP7_75t_L g4754 ( 
.A(n_4684),
.B(n_4721),
.C(n_4729),
.Y(n_4754)
);

HB1xp67_ASAP7_75t_L g4755 ( 
.A(n_4683),
.Y(n_4755)
);

NAND5xp2_ASAP7_75t_L g4756 ( 
.A(n_4696),
.B(n_4653),
.C(n_4654),
.D(n_4667),
.E(n_4641),
.Y(n_4756)
);

AOI211xp5_ASAP7_75t_L g4757 ( 
.A1(n_4720),
.A2(n_4658),
.B(n_462),
.C(n_460),
.Y(n_4757)
);

AND2x4_ASAP7_75t_L g4758 ( 
.A(n_4677),
.B(n_461),
.Y(n_4758)
);

AND2x2_ASAP7_75t_L g4759 ( 
.A(n_4678),
.B(n_461),
.Y(n_4759)
);

AND2x2_ASAP7_75t_L g4760 ( 
.A(n_4716),
.B(n_462),
.Y(n_4760)
);

INVx2_ASAP7_75t_L g4761 ( 
.A(n_4698),
.Y(n_4761)
);

INVx1_ASAP7_75t_L g4762 ( 
.A(n_4690),
.Y(n_4762)
);

INVx3_ASAP7_75t_L g4763 ( 
.A(n_4725),
.Y(n_4763)
);

AOI22xp33_ASAP7_75t_L g4764 ( 
.A1(n_4711),
.A2(n_465),
.B1(n_463),
.B2(n_464),
.Y(n_4764)
);

INVx1_ASAP7_75t_L g4765 ( 
.A(n_4714),
.Y(n_4765)
);

AND2x2_ASAP7_75t_L g4766 ( 
.A(n_4708),
.B(n_463),
.Y(n_4766)
);

AND2x2_ASAP7_75t_L g4767 ( 
.A(n_4701),
.B(n_464),
.Y(n_4767)
);

INVx1_ASAP7_75t_SL g4768 ( 
.A(n_4674),
.Y(n_4768)
);

INVx2_ASAP7_75t_L g4769 ( 
.A(n_4718),
.Y(n_4769)
);

AND2x4_ASAP7_75t_SL g4770 ( 
.A(n_4692),
.B(n_4676),
.Y(n_4770)
);

AND2x2_ASAP7_75t_L g4771 ( 
.A(n_4702),
.B(n_465),
.Y(n_4771)
);

INVx2_ASAP7_75t_SL g4772 ( 
.A(n_4697),
.Y(n_4772)
);

OR2x2_ASAP7_75t_L g4773 ( 
.A(n_4688),
.B(n_466),
.Y(n_4773)
);

INVx1_ASAP7_75t_L g4774 ( 
.A(n_4705),
.Y(n_4774)
);

AND2x2_ASAP7_75t_L g4775 ( 
.A(n_4706),
.B(n_467),
.Y(n_4775)
);

NAND2xp5_ASAP7_75t_L g4776 ( 
.A(n_4703),
.B(n_468),
.Y(n_4776)
);

NOR2xp33_ASAP7_75t_L g4777 ( 
.A(n_4735),
.B(n_4693),
.Y(n_4777)
);

OA211x2_ASAP7_75t_L g4778 ( 
.A1(n_4743),
.A2(n_4682),
.B(n_4709),
.C(n_4726),
.Y(n_4778)
);

NAND2x1_ASAP7_75t_L g4779 ( 
.A(n_4763),
.B(n_4723),
.Y(n_4779)
);

NAND2xp5_ASAP7_75t_L g4780 ( 
.A(n_4737),
.B(n_4755),
.Y(n_4780)
);

AND2x2_ASAP7_75t_SL g4781 ( 
.A(n_4770),
.B(n_4724),
.Y(n_4781)
);

INVx1_ASAP7_75t_L g4782 ( 
.A(n_4731),
.Y(n_4782)
);

NAND2xp5_ASAP7_75t_L g4783 ( 
.A(n_4749),
.B(n_4730),
.Y(n_4783)
);

NAND3xp33_ASAP7_75t_L g4784 ( 
.A(n_4754),
.B(n_4722),
.C(n_4719),
.Y(n_4784)
);

OR2x2_ASAP7_75t_L g4785 ( 
.A(n_4738),
.B(n_4728),
.Y(n_4785)
);

INVx1_ASAP7_75t_L g4786 ( 
.A(n_4747),
.Y(n_4786)
);

OR2x2_ASAP7_75t_L g4787 ( 
.A(n_4741),
.B(n_469),
.Y(n_4787)
);

INVxp67_ASAP7_75t_L g4788 ( 
.A(n_4732),
.Y(n_4788)
);

INVx1_ASAP7_75t_L g4789 ( 
.A(n_4739),
.Y(n_4789)
);

HB1xp67_ASAP7_75t_L g4790 ( 
.A(n_4740),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_4760),
.Y(n_4791)
);

OR2x2_ASAP7_75t_L g4792 ( 
.A(n_4773),
.B(n_471),
.Y(n_4792)
);

AND2x2_ASAP7_75t_L g4793 ( 
.A(n_4742),
.B(n_471),
.Y(n_4793)
);

NAND2xp5_ASAP7_75t_L g4794 ( 
.A(n_4766),
.B(n_472),
.Y(n_4794)
);

INVxp67_ASAP7_75t_SL g4795 ( 
.A(n_4769),
.Y(n_4795)
);

INVx1_ASAP7_75t_L g4796 ( 
.A(n_4746),
.Y(n_4796)
);

INVx2_ASAP7_75t_L g4797 ( 
.A(n_4753),
.Y(n_4797)
);

INVx1_ASAP7_75t_L g4798 ( 
.A(n_4736),
.Y(n_4798)
);

OR2x2_ASAP7_75t_L g4799 ( 
.A(n_4768),
.B(n_472),
.Y(n_4799)
);

AND2x2_ASAP7_75t_L g4800 ( 
.A(n_4761),
.B(n_474),
.Y(n_4800)
);

AND2x2_ASAP7_75t_L g4801 ( 
.A(n_4751),
.B(n_475),
.Y(n_4801)
);

INVx1_ASAP7_75t_SL g4802 ( 
.A(n_4752),
.Y(n_4802)
);

AND2x4_ASAP7_75t_L g4803 ( 
.A(n_4748),
.B(n_475),
.Y(n_4803)
);

INVx1_ASAP7_75t_L g4804 ( 
.A(n_4767),
.Y(n_4804)
);

NOR2xp33_ASAP7_75t_L g4805 ( 
.A(n_4756),
.B(n_477),
.Y(n_4805)
);

INVxp67_ASAP7_75t_SL g4806 ( 
.A(n_4776),
.Y(n_4806)
);

INVx1_ASAP7_75t_L g4807 ( 
.A(n_4771),
.Y(n_4807)
);

HB1xp67_ASAP7_75t_L g4808 ( 
.A(n_4758),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_4775),
.Y(n_4809)
);

NAND2xp5_ASAP7_75t_L g4810 ( 
.A(n_4734),
.B(n_478),
.Y(n_4810)
);

INVx1_ASAP7_75t_L g4811 ( 
.A(n_4759),
.Y(n_4811)
);

AND2x4_ASAP7_75t_L g4812 ( 
.A(n_4762),
.B(n_478),
.Y(n_4812)
);

OAI22xp33_ASAP7_75t_L g4813 ( 
.A1(n_4744),
.A2(n_482),
.B1(n_479),
.B2(n_481),
.Y(n_4813)
);

NOR2xp67_ASAP7_75t_SL g4814 ( 
.A(n_4765),
.B(n_479),
.Y(n_4814)
);

INVx2_ASAP7_75t_SL g4815 ( 
.A(n_4772),
.Y(n_4815)
);

INVx2_ASAP7_75t_L g4816 ( 
.A(n_4774),
.Y(n_4816)
);

INVx2_ASAP7_75t_L g4817 ( 
.A(n_4745),
.Y(n_4817)
);

OR2x2_ASAP7_75t_L g4818 ( 
.A(n_4764),
.B(n_482),
.Y(n_4818)
);

INVx1_ASAP7_75t_L g4819 ( 
.A(n_4750),
.Y(n_4819)
);

OAI22xp5_ASAP7_75t_L g4820 ( 
.A1(n_4733),
.A2(n_485),
.B1(n_483),
.B2(n_484),
.Y(n_4820)
);

NOR3xp33_ASAP7_75t_L g4821 ( 
.A(n_4757),
.B(n_483),
.C(n_484),
.Y(n_4821)
);

OAI211xp5_ASAP7_75t_L g4822 ( 
.A1(n_4733),
.A2(n_488),
.B(n_486),
.C(n_487),
.Y(n_4822)
);

INVxp67_ASAP7_75t_SL g4823 ( 
.A(n_4754),
.Y(n_4823)
);

NAND2xp5_ASAP7_75t_L g4824 ( 
.A(n_4735),
.B(n_486),
.Y(n_4824)
);

OAI31xp33_ASAP7_75t_SL g4825 ( 
.A1(n_4823),
.A2(n_490),
.A3(n_487),
.B(n_489),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4780),
.Y(n_4826)
);

INVx2_ASAP7_75t_L g4827 ( 
.A(n_4781),
.Y(n_4827)
);

OAI22xp33_ASAP7_75t_L g4828 ( 
.A1(n_4788),
.A2(n_4784),
.B1(n_4819),
.B2(n_4783),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_4808),
.Y(n_4829)
);

NOR2xp33_ASAP7_75t_SL g4830 ( 
.A(n_4777),
.B(n_489),
.Y(n_4830)
);

NOR2xp33_ASAP7_75t_L g4831 ( 
.A(n_4802),
.B(n_490),
.Y(n_4831)
);

INVx1_ASAP7_75t_L g4832 ( 
.A(n_4790),
.Y(n_4832)
);

INVx1_ASAP7_75t_L g4833 ( 
.A(n_4793),
.Y(n_4833)
);

NAND2xp5_ASAP7_75t_L g4834 ( 
.A(n_4782),
.B(n_4786),
.Y(n_4834)
);

NAND4xp75_ASAP7_75t_L g4835 ( 
.A(n_4778),
.B(n_4815),
.C(n_4789),
.D(n_4798),
.Y(n_4835)
);

INVxp67_ASAP7_75t_L g4836 ( 
.A(n_4814),
.Y(n_4836)
);

AND2x2_ASAP7_75t_L g4837 ( 
.A(n_4797),
.B(n_491),
.Y(n_4837)
);

INVx1_ASAP7_75t_L g4838 ( 
.A(n_4787),
.Y(n_4838)
);

INVx2_ASAP7_75t_L g4839 ( 
.A(n_4799),
.Y(n_4839)
);

AND2x2_ASAP7_75t_L g4840 ( 
.A(n_4795),
.B(n_491),
.Y(n_4840)
);

OAI31xp33_ASAP7_75t_L g4841 ( 
.A1(n_4822),
.A2(n_494),
.A3(n_492),
.B(n_493),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_4824),
.Y(n_4842)
);

INVx1_ASAP7_75t_L g4843 ( 
.A(n_4792),
.Y(n_4843)
);

NAND2xp5_ASAP7_75t_L g4844 ( 
.A(n_4805),
.B(n_4803),
.Y(n_4844)
);

INVx1_ASAP7_75t_SL g4845 ( 
.A(n_4779),
.Y(n_4845)
);

AOI211xp5_ASAP7_75t_L g4846 ( 
.A1(n_4813),
.A2(n_495),
.B(n_492),
.C(n_494),
.Y(n_4846)
);

NOR2xp33_ASAP7_75t_L g4847 ( 
.A(n_4791),
.B(n_495),
.Y(n_4847)
);

AND2x2_ASAP7_75t_L g4848 ( 
.A(n_4804),
.B(n_496),
.Y(n_4848)
);

INVx1_ASAP7_75t_SL g4849 ( 
.A(n_4800),
.Y(n_4849)
);

INVx1_ASAP7_75t_L g4850 ( 
.A(n_4801),
.Y(n_4850)
);

NOR2xp67_ASAP7_75t_L g4851 ( 
.A(n_4807),
.B(n_497),
.Y(n_4851)
);

AOI221xp5_ASAP7_75t_L g4852 ( 
.A1(n_4820),
.A2(n_501),
.B1(n_499),
.B2(n_500),
.C(n_502),
.Y(n_4852)
);

OAI21xp5_ASAP7_75t_L g4853 ( 
.A1(n_4810),
.A2(n_499),
.B(n_500),
.Y(n_4853)
);

AND2x2_ASAP7_75t_L g4854 ( 
.A(n_4809),
.B(n_501),
.Y(n_4854)
);

BUFx2_ASAP7_75t_L g4855 ( 
.A(n_4812),
.Y(n_4855)
);

AND2x2_ASAP7_75t_L g4856 ( 
.A(n_4811),
.B(n_4817),
.Y(n_4856)
);

INVx1_ASAP7_75t_L g4857 ( 
.A(n_4794),
.Y(n_4857)
);

HB1xp67_ASAP7_75t_L g4858 ( 
.A(n_4785),
.Y(n_4858)
);

XNOR2xp5_ASAP7_75t_L g4859 ( 
.A(n_4821),
.B(n_502),
.Y(n_4859)
);

INVx2_ASAP7_75t_SL g4860 ( 
.A(n_4816),
.Y(n_4860)
);

NAND2xp33_ASAP7_75t_L g4861 ( 
.A(n_4818),
.B(n_503),
.Y(n_4861)
);

INVx1_ASAP7_75t_L g4862 ( 
.A(n_4796),
.Y(n_4862)
);

HB1xp67_ASAP7_75t_L g4863 ( 
.A(n_4806),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4780),
.Y(n_4864)
);

OR2x2_ASAP7_75t_L g4865 ( 
.A(n_4780),
.B(n_505),
.Y(n_4865)
);

INVx1_ASAP7_75t_L g4866 ( 
.A(n_4780),
.Y(n_4866)
);

INVx2_ASAP7_75t_L g4867 ( 
.A(n_4781),
.Y(n_4867)
);

INVxp67_ASAP7_75t_SL g4868 ( 
.A(n_4788),
.Y(n_4868)
);

AND2x2_ASAP7_75t_L g4869 ( 
.A(n_4782),
.B(n_506),
.Y(n_4869)
);

AND2x2_ASAP7_75t_L g4870 ( 
.A(n_4782),
.B(n_506),
.Y(n_4870)
);

NOR2xp33_ASAP7_75t_SL g4871 ( 
.A(n_4781),
.B(n_507),
.Y(n_4871)
);

INVx2_ASAP7_75t_SL g4872 ( 
.A(n_4781),
.Y(n_4872)
);

NAND2xp5_ASAP7_75t_L g4873 ( 
.A(n_4823),
.B(n_507),
.Y(n_4873)
);

NAND2xp5_ASAP7_75t_L g4874 ( 
.A(n_4823),
.B(n_508),
.Y(n_4874)
);

NAND2xp5_ASAP7_75t_L g4875 ( 
.A(n_4823),
.B(n_508),
.Y(n_4875)
);

OR2x2_ASAP7_75t_L g4876 ( 
.A(n_4780),
.B(n_509),
.Y(n_4876)
);

INVx2_ASAP7_75t_L g4877 ( 
.A(n_4781),
.Y(n_4877)
);

INVx1_ASAP7_75t_L g4878 ( 
.A(n_4780),
.Y(n_4878)
);

INVxp67_ASAP7_75t_L g4879 ( 
.A(n_4780),
.Y(n_4879)
);

NAND2x1_ASAP7_75t_L g4880 ( 
.A(n_4782),
.B(n_509),
.Y(n_4880)
);

NAND2x1p5_ASAP7_75t_L g4881 ( 
.A(n_4802),
.B(n_510),
.Y(n_4881)
);

AND2x2_ASAP7_75t_L g4882 ( 
.A(n_4782),
.B(n_510),
.Y(n_4882)
);

AND2x2_ASAP7_75t_L g4883 ( 
.A(n_4782),
.B(n_511),
.Y(n_4883)
);

NAND5xp2_ASAP7_75t_L g4884 ( 
.A(n_4829),
.B(n_513),
.C(n_511),
.D(n_512),
.E(n_515),
.Y(n_4884)
);

INVx1_ASAP7_75t_L g4885 ( 
.A(n_4881),
.Y(n_4885)
);

XOR2xp5_ASAP7_75t_L g4886 ( 
.A(n_4859),
.B(n_512),
.Y(n_4886)
);

INVx1_ASAP7_75t_L g4887 ( 
.A(n_4880),
.Y(n_4887)
);

INVxp67_ASAP7_75t_L g4888 ( 
.A(n_4871),
.Y(n_4888)
);

OAI21xp5_ASAP7_75t_SL g4889 ( 
.A1(n_4825),
.A2(n_513),
.B(n_515),
.Y(n_4889)
);

NAND2xp5_ASAP7_75t_L g4890 ( 
.A(n_4845),
.B(n_4872),
.Y(n_4890)
);

INVxp67_ASAP7_75t_L g4891 ( 
.A(n_4830),
.Y(n_4891)
);

OR2x2_ASAP7_75t_L g4892 ( 
.A(n_4844),
.B(n_516),
.Y(n_4892)
);

INVx1_ASAP7_75t_L g4893 ( 
.A(n_4851),
.Y(n_4893)
);

OAI221xp5_ASAP7_75t_SL g4894 ( 
.A1(n_4828),
.A2(n_518),
.B1(n_516),
.B2(n_517),
.C(n_519),
.Y(n_4894)
);

NAND2xp5_ASAP7_75t_L g4895 ( 
.A(n_4827),
.B(n_518),
.Y(n_4895)
);

NAND2xp5_ASAP7_75t_L g4896 ( 
.A(n_4867),
.B(n_519),
.Y(n_4896)
);

AOI221xp5_ASAP7_75t_L g4897 ( 
.A1(n_4868),
.A2(n_522),
.B1(n_525),
.B2(n_521),
.C(n_523),
.Y(n_4897)
);

OAI22xp33_ASAP7_75t_L g4898 ( 
.A1(n_4877),
.A2(n_522),
.B1(n_520),
.B2(n_521),
.Y(n_4898)
);

INVx1_ASAP7_75t_L g4899 ( 
.A(n_4855),
.Y(n_4899)
);

INVx1_ASAP7_75t_L g4900 ( 
.A(n_4840),
.Y(n_4900)
);

OA22x2_ASAP7_75t_L g4901 ( 
.A1(n_4836),
.A2(n_4832),
.B1(n_4833),
.B2(n_4849),
.Y(n_4901)
);

OAI22xp33_ASAP7_75t_SL g4902 ( 
.A1(n_4873),
.A2(n_528),
.B1(n_525),
.B2(n_526),
.Y(n_4902)
);

NOR3xp33_ASAP7_75t_SL g4903 ( 
.A(n_4835),
.B(n_4834),
.C(n_4826),
.Y(n_4903)
);

NAND2xp5_ASAP7_75t_L g4904 ( 
.A(n_4869),
.B(n_4870),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4858),
.Y(n_4905)
);

NOR2xp67_ASAP7_75t_L g4906 ( 
.A(n_4863),
.B(n_530),
.Y(n_4906)
);

NAND2xp5_ASAP7_75t_L g4907 ( 
.A(n_4882),
.B(n_530),
.Y(n_4907)
);

NAND2xp5_ASAP7_75t_L g4908 ( 
.A(n_4883),
.B(n_4837),
.Y(n_4908)
);

OAI22xp33_ASAP7_75t_L g4909 ( 
.A1(n_4874),
.A2(n_533),
.B1(n_531),
.B2(n_532),
.Y(n_4909)
);

NAND2xp5_ASAP7_75t_L g4910 ( 
.A(n_4848),
.B(n_531),
.Y(n_4910)
);

NAND2xp5_ASAP7_75t_L g4911 ( 
.A(n_4854),
.B(n_532),
.Y(n_4911)
);

INVxp67_ASAP7_75t_L g4912 ( 
.A(n_4831),
.Y(n_4912)
);

NAND2x1_ASAP7_75t_L g4913 ( 
.A(n_4838),
.B(n_534),
.Y(n_4913)
);

HB1xp67_ASAP7_75t_L g4914 ( 
.A(n_4865),
.Y(n_4914)
);

INVxp67_ASAP7_75t_SL g4915 ( 
.A(n_4875),
.Y(n_4915)
);

NOR2xp67_ASAP7_75t_L g4916 ( 
.A(n_4860),
.B(n_534),
.Y(n_4916)
);

BUFx12f_ASAP7_75t_L g4917 ( 
.A(n_4876),
.Y(n_4917)
);

INVx1_ASAP7_75t_SL g4918 ( 
.A(n_4856),
.Y(n_4918)
);

OAI21xp5_ASAP7_75t_L g4919 ( 
.A1(n_4879),
.A2(n_535),
.B(n_536),
.Y(n_4919)
);

A2O1A1Ixp33_ASAP7_75t_L g4920 ( 
.A1(n_4841),
.A2(n_539),
.B(n_540),
.C(n_537),
.Y(n_4920)
);

AOI321xp33_ASAP7_75t_SL g4921 ( 
.A1(n_4847),
.A2(n_539),
.A3(n_542),
.B1(n_536),
.B2(n_537),
.C(n_541),
.Y(n_4921)
);

INVx1_ASAP7_75t_SL g4922 ( 
.A(n_4839),
.Y(n_4922)
);

OAI22xp5_ASAP7_75t_L g4923 ( 
.A1(n_4864),
.A2(n_543),
.B1(n_541),
.B2(n_542),
.Y(n_4923)
);

INVx1_ASAP7_75t_L g4924 ( 
.A(n_4850),
.Y(n_4924)
);

INVx1_ASAP7_75t_L g4925 ( 
.A(n_4866),
.Y(n_4925)
);

OA21x2_ASAP7_75t_L g4926 ( 
.A1(n_4853),
.A2(n_543),
.B(n_544),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4878),
.Y(n_4927)
);

AOI22xp5_ASAP7_75t_L g4928 ( 
.A1(n_4861),
.A2(n_4857),
.B1(n_4843),
.B2(n_4842),
.Y(n_4928)
);

INVx1_ASAP7_75t_L g4929 ( 
.A(n_4862),
.Y(n_4929)
);

NAND2xp5_ASAP7_75t_SL g4930 ( 
.A(n_4846),
.B(n_545),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4852),
.Y(n_4931)
);

AOI21xp5_ASAP7_75t_L g4932 ( 
.A1(n_4872),
.A2(n_545),
.B(n_546),
.Y(n_4932)
);

INVx1_ASAP7_75t_L g4933 ( 
.A(n_4881),
.Y(n_4933)
);

INVx1_ASAP7_75t_L g4934 ( 
.A(n_4881),
.Y(n_4934)
);

INVx1_ASAP7_75t_L g4935 ( 
.A(n_4881),
.Y(n_4935)
);

OAI22xp5_ASAP7_75t_L g4936 ( 
.A1(n_4835),
.A2(n_548),
.B1(n_546),
.B2(n_547),
.Y(n_4936)
);

INVx1_ASAP7_75t_L g4937 ( 
.A(n_4881),
.Y(n_4937)
);

INVxp67_ASAP7_75t_L g4938 ( 
.A(n_4871),
.Y(n_4938)
);

HB1xp67_ASAP7_75t_L g4939 ( 
.A(n_4851),
.Y(n_4939)
);

OAI222xp33_ASAP7_75t_L g4940 ( 
.A1(n_4845),
.A2(n_551),
.B1(n_553),
.B2(n_549),
.C1(n_550),
.C2(n_552),
.Y(n_4940)
);

O2A1O1Ixp5_ASAP7_75t_L g4941 ( 
.A1(n_4868),
.A2(n_551),
.B(n_549),
.C(n_550),
.Y(n_4941)
);

INVx1_ASAP7_75t_L g4942 ( 
.A(n_4881),
.Y(n_4942)
);

OAI22xp33_ASAP7_75t_L g4943 ( 
.A1(n_4871),
.A2(n_556),
.B1(n_553),
.B2(n_555),
.Y(n_4943)
);

AND2x2_ASAP7_75t_L g4944 ( 
.A(n_4872),
.B(n_558),
.Y(n_4944)
);

AND2x2_ASAP7_75t_L g4945 ( 
.A(n_4872),
.B(n_558),
.Y(n_4945)
);

AOI22xp5_ASAP7_75t_L g4946 ( 
.A1(n_4872),
.A2(n_561),
.B1(n_559),
.B2(n_560),
.Y(n_4946)
);

OAI21xp33_ASAP7_75t_L g4947 ( 
.A1(n_4872),
.A2(n_571),
.B(n_560),
.Y(n_4947)
);

INVx1_ASAP7_75t_L g4948 ( 
.A(n_4881),
.Y(n_4948)
);

AOI21xp5_ASAP7_75t_L g4949 ( 
.A1(n_4872),
.A2(n_561),
.B(n_563),
.Y(n_4949)
);

OAI32xp33_ASAP7_75t_L g4950 ( 
.A1(n_4845),
.A2(n_565),
.A3(n_563),
.B1(n_564),
.B2(n_566),
.Y(n_4950)
);

INVx2_ASAP7_75t_L g4951 ( 
.A(n_4881),
.Y(n_4951)
);

INVx2_ASAP7_75t_L g4952 ( 
.A(n_4881),
.Y(n_4952)
);

NAND2xp5_ASAP7_75t_L g4953 ( 
.A(n_4845),
.B(n_564),
.Y(n_4953)
);

AOI221x1_ASAP7_75t_L g4954 ( 
.A1(n_4832),
.A2(n_570),
.B1(n_573),
.B2(n_569),
.C(n_572),
.Y(n_4954)
);

OAI21xp5_ASAP7_75t_L g4955 ( 
.A1(n_4835),
.A2(n_566),
.B(n_569),
.Y(n_4955)
);

AOI222xp33_ASAP7_75t_L g4956 ( 
.A1(n_4828),
.A2(n_573),
.B1(n_575),
.B2(n_570),
.C1(n_572),
.C2(n_574),
.Y(n_4956)
);

O2A1O1Ixp33_ASAP7_75t_SL g4957 ( 
.A1(n_4845),
.A2(n_577),
.B(n_574),
.C(n_576),
.Y(n_4957)
);

NAND2xp5_ASAP7_75t_L g4958 ( 
.A(n_4845),
.B(n_576),
.Y(n_4958)
);

AND2x2_ASAP7_75t_L g4959 ( 
.A(n_4872),
.B(n_578),
.Y(n_4959)
);

OAI21xp5_ASAP7_75t_L g4960 ( 
.A1(n_4835),
.A2(n_579),
.B(n_580),
.Y(n_4960)
);

INVx1_ASAP7_75t_L g4961 ( 
.A(n_4881),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_4881),
.Y(n_4962)
);

OR2x2_ASAP7_75t_L g4963 ( 
.A(n_4881),
.B(n_581),
.Y(n_4963)
);

AOI22xp5_ASAP7_75t_L g4964 ( 
.A1(n_4872),
.A2(n_584),
.B1(n_581),
.B2(n_582),
.Y(n_4964)
);

NAND2xp5_ASAP7_75t_L g4965 ( 
.A(n_4845),
.B(n_582),
.Y(n_4965)
);

OAI322xp33_ASAP7_75t_L g4966 ( 
.A1(n_4828),
.A2(n_589),
.A3(n_588),
.B1(n_586),
.B2(n_584),
.C1(n_585),
.C2(n_587),
.Y(n_4966)
);

INVxp67_ASAP7_75t_L g4967 ( 
.A(n_4871),
.Y(n_4967)
);

AND2x2_ASAP7_75t_L g4968 ( 
.A(n_4872),
.B(n_587),
.Y(n_4968)
);

NAND2xp5_ASAP7_75t_L g4969 ( 
.A(n_4845),
.B(n_589),
.Y(n_4969)
);

INVxp67_ASAP7_75t_L g4970 ( 
.A(n_4871),
.Y(n_4970)
);

OR2x2_ASAP7_75t_L g4971 ( 
.A(n_4881),
.B(n_590),
.Y(n_4971)
);

NAND3xp33_ASAP7_75t_L g4972 ( 
.A(n_4825),
.B(n_591),
.C(n_592),
.Y(n_4972)
);

INVxp67_ASAP7_75t_SL g4973 ( 
.A(n_4881),
.Y(n_4973)
);

OAI221xp5_ASAP7_75t_L g4974 ( 
.A1(n_4872),
.A2(n_594),
.B1(n_592),
.B2(n_593),
.C(n_595),
.Y(n_4974)
);

OAI221xp5_ASAP7_75t_L g4975 ( 
.A1(n_4872),
.A2(n_595),
.B1(n_593),
.B2(n_594),
.C(n_597),
.Y(n_4975)
);

INVx3_ASAP7_75t_SL g4976 ( 
.A(n_4918),
.Y(n_4976)
);

AND2x2_ASAP7_75t_L g4977 ( 
.A(n_4899),
.B(n_597),
.Y(n_4977)
);

OR2x2_ASAP7_75t_L g4978 ( 
.A(n_4887),
.B(n_598),
.Y(n_4978)
);

XOR2x2_ASAP7_75t_L g4979 ( 
.A(n_4972),
.B(n_599),
.Y(n_4979)
);

NAND4xp75_ASAP7_75t_L g4980 ( 
.A(n_4955),
.B(n_602),
.C(n_599),
.D(n_601),
.Y(n_4980)
);

NOR2x1_ASAP7_75t_L g4981 ( 
.A(n_4916),
.B(n_4906),
.Y(n_4981)
);

AOI211x1_ASAP7_75t_SL g4982 ( 
.A1(n_4936),
.A2(n_603),
.B(n_601),
.C(n_602),
.Y(n_4982)
);

NAND2x1p5_ASAP7_75t_L g4983 ( 
.A(n_4885),
.B(n_4933),
.Y(n_4983)
);

OR2x2_ASAP7_75t_L g4984 ( 
.A(n_4939),
.B(n_603),
.Y(n_4984)
);

NAND2xp5_ASAP7_75t_L g4985 ( 
.A(n_4889),
.B(n_605),
.Y(n_4985)
);

O2A1O1Ixp33_ASAP7_75t_SL g4986 ( 
.A1(n_4940),
.A2(n_4920),
.B(n_4913),
.C(n_4934),
.Y(n_4986)
);

OAI32xp33_ASAP7_75t_L g4987 ( 
.A1(n_4960),
.A2(n_625),
.A3(n_634),
.B1(n_617),
.B2(n_606),
.Y(n_4987)
);

OAI21xp5_ASAP7_75t_L g4988 ( 
.A1(n_4890),
.A2(n_606),
.B(n_607),
.Y(n_4988)
);

OR2x2_ASAP7_75t_L g4989 ( 
.A(n_4893),
.B(n_608),
.Y(n_4989)
);

OR2x2_ASAP7_75t_L g4990 ( 
.A(n_4935),
.B(n_608),
.Y(n_4990)
);

NAND2x1_ASAP7_75t_L g4991 ( 
.A(n_4937),
.B(n_609),
.Y(n_4991)
);

AOI221xp5_ASAP7_75t_SL g4992 ( 
.A1(n_4888),
.A2(n_611),
.B1(n_609),
.B2(n_610),
.C(n_614),
.Y(n_4992)
);

OR2x2_ASAP7_75t_L g4993 ( 
.A(n_4942),
.B(n_610),
.Y(n_4993)
);

NAND2xp5_ASAP7_75t_SL g4994 ( 
.A(n_4951),
.B(n_616),
.Y(n_4994)
);

OAI21xp5_ASAP7_75t_SL g4995 ( 
.A1(n_4938),
.A2(n_4970),
.B(n_4967),
.Y(n_4995)
);

AOI211xp5_ASAP7_75t_L g4996 ( 
.A1(n_4894),
.A2(n_619),
.B(n_617),
.C(n_618),
.Y(n_4996)
);

NAND2xp33_ASAP7_75t_L g4997 ( 
.A(n_4952),
.B(n_619),
.Y(n_4997)
);

INVx1_ASAP7_75t_L g4998 ( 
.A(n_4963),
.Y(n_4998)
);

INVx1_ASAP7_75t_SL g4999 ( 
.A(n_4971),
.Y(n_4999)
);

INVx2_ASAP7_75t_SL g5000 ( 
.A(n_4948),
.Y(n_5000)
);

INVx1_ASAP7_75t_L g5001 ( 
.A(n_4944),
.Y(n_5001)
);

INVx2_ASAP7_75t_SL g5002 ( 
.A(n_4961),
.Y(n_5002)
);

INVx1_ASAP7_75t_L g5003 ( 
.A(n_4945),
.Y(n_5003)
);

NAND2xp5_ASAP7_75t_L g5004 ( 
.A(n_4959),
.B(n_620),
.Y(n_5004)
);

OAI22xp5_ASAP7_75t_L g5005 ( 
.A1(n_4973),
.A2(n_622),
.B1(n_620),
.B2(n_621),
.Y(n_5005)
);

AND2x2_ASAP7_75t_L g5006 ( 
.A(n_4968),
.B(n_621),
.Y(n_5006)
);

OR2x2_ASAP7_75t_L g5007 ( 
.A(n_4962),
.B(n_623),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4957),
.Y(n_5008)
);

INVx1_ASAP7_75t_SL g5009 ( 
.A(n_4922),
.Y(n_5009)
);

AOI21xp33_ASAP7_75t_SL g5010 ( 
.A1(n_4901),
.A2(n_623),
.B(n_624),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_4953),
.Y(n_5011)
);

OA22x2_ASAP7_75t_L g5012 ( 
.A1(n_4928),
.A2(n_627),
.B1(n_625),
.B2(n_626),
.Y(n_5012)
);

NAND2x1p5_ASAP7_75t_L g5013 ( 
.A(n_4905),
.B(n_630),
.Y(n_5013)
);

INVx1_ASAP7_75t_L g5014 ( 
.A(n_4958),
.Y(n_5014)
);

INVxp67_ASAP7_75t_L g5015 ( 
.A(n_4884),
.Y(n_5015)
);

OAI321xp33_ASAP7_75t_L g5016 ( 
.A1(n_4891),
.A2(n_632),
.A3(n_634),
.B1(n_629),
.B2(n_631),
.C(n_633),
.Y(n_5016)
);

NAND2xp5_ASAP7_75t_L g5017 ( 
.A(n_4900),
.B(n_629),
.Y(n_5017)
);

HB1xp67_ASAP7_75t_L g5018 ( 
.A(n_4926),
.Y(n_5018)
);

AND2x2_ASAP7_75t_L g5019 ( 
.A(n_4903),
.B(n_631),
.Y(n_5019)
);

OA211x2_ASAP7_75t_L g5020 ( 
.A1(n_4947),
.A2(n_636),
.B(n_633),
.C(n_635),
.Y(n_5020)
);

AOI32xp33_ASAP7_75t_L g5021 ( 
.A1(n_4924),
.A2(n_638),
.A3(n_640),
.B1(n_637),
.B2(n_639),
.Y(n_5021)
);

OR2x2_ASAP7_75t_L g5022 ( 
.A(n_4965),
.B(n_636),
.Y(n_5022)
);

INVx1_ASAP7_75t_L g5023 ( 
.A(n_4969),
.Y(n_5023)
);

NAND2xp5_ASAP7_75t_L g5024 ( 
.A(n_4932),
.B(n_638),
.Y(n_5024)
);

XOR2x2_ASAP7_75t_L g5025 ( 
.A(n_4886),
.B(n_640),
.Y(n_5025)
);

OAI21xp5_ASAP7_75t_SL g5026 ( 
.A1(n_4956),
.A2(n_641),
.B(n_642),
.Y(n_5026)
);

NOR2xp33_ASAP7_75t_L g5027 ( 
.A(n_4966),
.B(n_4974),
.Y(n_5027)
);

XNOR2xp5_ASAP7_75t_L g5028 ( 
.A(n_4946),
.B(n_641),
.Y(n_5028)
);

BUFx2_ASAP7_75t_L g5029 ( 
.A(n_4917),
.Y(n_5029)
);

INVx1_ASAP7_75t_L g5030 ( 
.A(n_4892),
.Y(n_5030)
);

INVx1_ASAP7_75t_SL g5031 ( 
.A(n_4926),
.Y(n_5031)
);

INVx1_ASAP7_75t_L g5032 ( 
.A(n_4904),
.Y(n_5032)
);

AND2x2_ASAP7_75t_L g5033 ( 
.A(n_4914),
.B(n_642),
.Y(n_5033)
);

NOR2xp33_ASAP7_75t_L g5034 ( 
.A(n_4975),
.B(n_643),
.Y(n_5034)
);

AND2x4_ASAP7_75t_SL g5035 ( 
.A(n_4929),
.B(n_643),
.Y(n_5035)
);

NAND2xp5_ASAP7_75t_SL g5036 ( 
.A(n_4902),
.B(n_644),
.Y(n_5036)
);

INVx2_ASAP7_75t_SL g5037 ( 
.A(n_4908),
.Y(n_5037)
);

INVx1_ASAP7_75t_L g5038 ( 
.A(n_4895),
.Y(n_5038)
);

INVx2_ASAP7_75t_SL g5039 ( 
.A(n_4896),
.Y(n_5039)
);

INVx1_ASAP7_75t_L g5040 ( 
.A(n_4910),
.Y(n_5040)
);

INVx1_ASAP7_75t_L g5041 ( 
.A(n_4911),
.Y(n_5041)
);

NAND4xp25_ASAP7_75t_L g5042 ( 
.A(n_4931),
.B(n_647),
.C(n_644),
.D(n_645),
.Y(n_5042)
);

NAND2xp5_ASAP7_75t_L g5043 ( 
.A(n_4949),
.B(n_645),
.Y(n_5043)
);

NAND2xp5_ASAP7_75t_L g5044 ( 
.A(n_4943),
.B(n_647),
.Y(n_5044)
);

NOR2xp33_ASAP7_75t_L g5045 ( 
.A(n_4907),
.B(n_648),
.Y(n_5045)
);

NOR2xp33_ASAP7_75t_L g5046 ( 
.A(n_4912),
.B(n_649),
.Y(n_5046)
);

INVx2_ASAP7_75t_L g5047 ( 
.A(n_4941),
.Y(n_5047)
);

INVx1_ASAP7_75t_L g5048 ( 
.A(n_4964),
.Y(n_5048)
);

INVx1_ASAP7_75t_L g5049 ( 
.A(n_4950),
.Y(n_5049)
);

INVx1_ASAP7_75t_SL g5050 ( 
.A(n_4930),
.Y(n_5050)
);

AOI32xp33_ASAP7_75t_L g5051 ( 
.A1(n_4925),
.A2(n_651),
.A3(n_653),
.B1(n_650),
.B2(n_652),
.Y(n_5051)
);

INVx2_ASAP7_75t_L g5052 ( 
.A(n_4927),
.Y(n_5052)
);

NAND2xp5_ASAP7_75t_L g5053 ( 
.A(n_4954),
.B(n_649),
.Y(n_5053)
);

INVx1_ASAP7_75t_L g5054 ( 
.A(n_4923),
.Y(n_5054)
);

AOI211xp5_ASAP7_75t_L g5055 ( 
.A1(n_4898),
.A2(n_652),
.B(n_650),
.C(n_651),
.Y(n_5055)
);

INVx1_ASAP7_75t_L g5056 ( 
.A(n_4919),
.Y(n_5056)
);

NOR2xp33_ASAP7_75t_L g5057 ( 
.A(n_4909),
.B(n_653),
.Y(n_5057)
);

NAND2xp5_ASAP7_75t_L g5058 ( 
.A(n_4897),
.B(n_654),
.Y(n_5058)
);

INVx1_ASAP7_75t_L g5059 ( 
.A(n_4915),
.Y(n_5059)
);

NAND2xp5_ASAP7_75t_L g5060 ( 
.A(n_4921),
.B(n_655),
.Y(n_5060)
);

NOR2xp33_ASAP7_75t_L g5061 ( 
.A(n_4889),
.B(n_655),
.Y(n_5061)
);

OAI21xp5_ASAP7_75t_L g5062 ( 
.A1(n_4972),
.A2(n_656),
.B(n_657),
.Y(n_5062)
);

AOI322xp5_ASAP7_75t_L g5063 ( 
.A1(n_5019),
.A2(n_663),
.A3(n_661),
.B1(n_659),
.B2(n_657),
.C1(n_658),
.C2(n_660),
.Y(n_5063)
);

NAND2xp5_ASAP7_75t_L g5064 ( 
.A(n_5008),
.B(n_659),
.Y(n_5064)
);

AOI31xp33_ASAP7_75t_L g5065 ( 
.A1(n_4981),
.A2(n_673),
.A3(n_681),
.B(n_663),
.Y(n_5065)
);

INVx1_ASAP7_75t_SL g5066 ( 
.A(n_4976),
.Y(n_5066)
);

INVx1_ASAP7_75t_SL g5067 ( 
.A(n_5031),
.Y(n_5067)
);

INVxp67_ASAP7_75t_L g5068 ( 
.A(n_5018),
.Y(n_5068)
);

INVx2_ASAP7_75t_L g5069 ( 
.A(n_4983),
.Y(n_5069)
);

INVx1_ASAP7_75t_L g5070 ( 
.A(n_4991),
.Y(n_5070)
);

AOI221xp5_ASAP7_75t_L g5071 ( 
.A1(n_5010),
.A2(n_666),
.B1(n_664),
.B2(n_665),
.C(n_667),
.Y(n_5071)
);

NAND2xp5_ASAP7_75t_L g5072 ( 
.A(n_5009),
.B(n_665),
.Y(n_5072)
);

OAI22x1_ASAP7_75t_L g5073 ( 
.A1(n_5047),
.A2(n_668),
.B1(n_666),
.B2(n_667),
.Y(n_5073)
);

INVx1_ASAP7_75t_L g5074 ( 
.A(n_5012),
.Y(n_5074)
);

NAND2xp5_ASAP7_75t_L g5075 ( 
.A(n_5015),
.B(n_668),
.Y(n_5075)
);

INVx1_ASAP7_75t_L g5076 ( 
.A(n_4978),
.Y(n_5076)
);

INVx1_ASAP7_75t_L g5077 ( 
.A(n_4984),
.Y(n_5077)
);

NOR5xp2_ASAP7_75t_L g5078 ( 
.A(n_4995),
.B(n_673),
.C(n_669),
.D(n_670),
.E(n_674),
.Y(n_5078)
);

INVx2_ASAP7_75t_L g5079 ( 
.A(n_5013),
.Y(n_5079)
);

AOI222xp33_ASAP7_75t_L g5080 ( 
.A1(n_5029),
.A2(n_675),
.B1(n_677),
.B2(n_670),
.C1(n_674),
.C2(n_676),
.Y(n_5080)
);

INVx1_ASAP7_75t_L g5081 ( 
.A(n_5006),
.Y(n_5081)
);

NAND3xp33_ASAP7_75t_L g5082 ( 
.A(n_4996),
.B(n_4997),
.C(n_5055),
.Y(n_5082)
);

INVx1_ASAP7_75t_L g5083 ( 
.A(n_5033),
.Y(n_5083)
);

INVx2_ASAP7_75t_L g5084 ( 
.A(n_4989),
.Y(n_5084)
);

AOI222xp33_ASAP7_75t_L g5085 ( 
.A1(n_5049),
.A2(n_678),
.B1(n_680),
.B2(n_675),
.C1(n_676),
.C2(n_679),
.Y(n_5085)
);

INVx1_ASAP7_75t_L g5086 ( 
.A(n_5025),
.Y(n_5086)
);

INVx1_ASAP7_75t_L g5087 ( 
.A(n_4977),
.Y(n_5087)
);

INVx1_ASAP7_75t_L g5088 ( 
.A(n_5035),
.Y(n_5088)
);

NAND2xp5_ASAP7_75t_L g5089 ( 
.A(n_5000),
.B(n_680),
.Y(n_5089)
);

O2A1O1Ixp33_ASAP7_75t_L g5090 ( 
.A1(n_5053),
.A2(n_684),
.B(n_682),
.C(n_683),
.Y(n_5090)
);

NOR2x1_ASAP7_75t_L g5091 ( 
.A(n_4980),
.B(n_5042),
.Y(n_5091)
);

INVx1_ASAP7_75t_L g5092 ( 
.A(n_4990),
.Y(n_5092)
);

OAI322xp33_ASAP7_75t_L g5093 ( 
.A1(n_5002),
.A2(n_689),
.A3(n_688),
.B1(n_686),
.B2(n_684),
.C1(n_685),
.C2(n_687),
.Y(n_5093)
);

NAND2xp5_ASAP7_75t_L g5094 ( 
.A(n_5061),
.B(n_4992),
.Y(n_5094)
);

NAND2xp5_ASAP7_75t_L g5095 ( 
.A(n_4982),
.B(n_685),
.Y(n_5095)
);

OAI22xp33_ASAP7_75t_L g5096 ( 
.A1(n_5060),
.A2(n_689),
.B1(n_686),
.B2(n_688),
.Y(n_5096)
);

OAI321xp33_ASAP7_75t_L g5097 ( 
.A1(n_5027),
.A2(n_692),
.A3(n_694),
.B1(n_690),
.B2(n_691),
.C(n_693),
.Y(n_5097)
);

INVx1_ASAP7_75t_SL g5098 ( 
.A(n_4993),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_5007),
.Y(n_5099)
);

NAND2xp5_ASAP7_75t_L g5100 ( 
.A(n_5001),
.B(n_690),
.Y(n_5100)
);

AND2x2_ASAP7_75t_L g5101 ( 
.A(n_5003),
.B(n_693),
.Y(n_5101)
);

INVx1_ASAP7_75t_L g5102 ( 
.A(n_5004),
.Y(n_5102)
);

INVx1_ASAP7_75t_L g5103 ( 
.A(n_4979),
.Y(n_5103)
);

INVx2_ASAP7_75t_L g5104 ( 
.A(n_5022),
.Y(n_5104)
);

INVx1_ASAP7_75t_L g5105 ( 
.A(n_5024),
.Y(n_5105)
);

NAND2xp5_ASAP7_75t_L g5106 ( 
.A(n_5021),
.B(n_694),
.Y(n_5106)
);

INVx2_ASAP7_75t_SL g5107 ( 
.A(n_4994),
.Y(n_5107)
);

OA21x2_ASAP7_75t_L g5108 ( 
.A1(n_5017),
.A2(n_696),
.B(n_697),
.Y(n_5108)
);

OAI21xp5_ASAP7_75t_SL g5109 ( 
.A1(n_5026),
.A2(n_696),
.B(n_697),
.Y(n_5109)
);

AOI221xp5_ASAP7_75t_L g5110 ( 
.A1(n_4986),
.A2(n_701),
.B1(n_699),
.B2(n_700),
.C(n_702),
.Y(n_5110)
);

INVx1_ASAP7_75t_SL g5111 ( 
.A(n_4999),
.Y(n_5111)
);

AND2x2_ASAP7_75t_L g5112 ( 
.A(n_5062),
.B(n_5037),
.Y(n_5112)
);

INVx1_ASAP7_75t_L g5113 ( 
.A(n_5043),
.Y(n_5113)
);

NAND2xp5_ASAP7_75t_L g5114 ( 
.A(n_5051),
.B(n_699),
.Y(n_5114)
);

OR2x2_ASAP7_75t_L g5115 ( 
.A(n_4985),
.B(n_700),
.Y(n_5115)
);

NOR2xp33_ASAP7_75t_L g5116 ( 
.A(n_4987),
.B(n_703),
.Y(n_5116)
);

AO22x2_ASAP7_75t_L g5117 ( 
.A1(n_5050),
.A2(n_706),
.B1(n_704),
.B2(n_705),
.Y(n_5117)
);

INVx1_ASAP7_75t_L g5118 ( 
.A(n_5020),
.Y(n_5118)
);

INVx1_ASAP7_75t_L g5119 ( 
.A(n_5028),
.Y(n_5119)
);

AND2x2_ASAP7_75t_L g5120 ( 
.A(n_4998),
.B(n_705),
.Y(n_5120)
);

AO22x1_ASAP7_75t_L g5121 ( 
.A1(n_5057),
.A2(n_709),
.B1(n_707),
.B2(n_708),
.Y(n_5121)
);

AOI221x1_ASAP7_75t_L g5122 ( 
.A1(n_4988),
.A2(n_5058),
.B1(n_5059),
.B2(n_5032),
.C(n_5046),
.Y(n_5122)
);

XNOR2xp5_ASAP7_75t_L g5123 ( 
.A(n_5048),
.B(n_707),
.Y(n_5123)
);

OAI21xp33_ASAP7_75t_SL g5124 ( 
.A1(n_5036),
.A2(n_708),
.B(n_709),
.Y(n_5124)
);

INVx1_ASAP7_75t_L g5125 ( 
.A(n_5044),
.Y(n_5125)
);

OR2x2_ASAP7_75t_L g5126 ( 
.A(n_5054),
.B(n_710),
.Y(n_5126)
);

AOI22xp5_ASAP7_75t_L g5127 ( 
.A1(n_5034),
.A2(n_712),
.B1(n_710),
.B2(n_711),
.Y(n_5127)
);

OAI221xp5_ASAP7_75t_L g5128 ( 
.A1(n_5052),
.A2(n_714),
.B1(n_711),
.B2(n_713),
.C(n_715),
.Y(n_5128)
);

AOI22xp33_ASAP7_75t_L g5129 ( 
.A1(n_5039),
.A2(n_717),
.B1(n_714),
.B2(n_716),
.Y(n_5129)
);

INVx1_ASAP7_75t_L g5130 ( 
.A(n_5005),
.Y(n_5130)
);

NOR2x1_ASAP7_75t_L g5131 ( 
.A(n_5030),
.B(n_716),
.Y(n_5131)
);

INVxp67_ASAP7_75t_L g5132 ( 
.A(n_5045),
.Y(n_5132)
);

NAND2xp5_ASAP7_75t_L g5133 ( 
.A(n_5011),
.B(n_717),
.Y(n_5133)
);

O2A1O1Ixp33_ASAP7_75t_L g5134 ( 
.A1(n_5016),
.A2(n_721),
.B(n_719),
.C(n_720),
.Y(n_5134)
);

O2A1O1Ixp33_ASAP7_75t_L g5135 ( 
.A1(n_5056),
.A2(n_724),
.B(n_721),
.C(n_723),
.Y(n_5135)
);

NAND2xp5_ASAP7_75t_SL g5136 ( 
.A(n_5014),
.B(n_724),
.Y(n_5136)
);

OAI22xp33_ASAP7_75t_L g5137 ( 
.A1(n_5023),
.A2(n_727),
.B1(n_725),
.B2(n_726),
.Y(n_5137)
);

INVx1_ASAP7_75t_L g5138 ( 
.A(n_5040),
.Y(n_5138)
);

INVx1_ASAP7_75t_L g5139 ( 
.A(n_5041),
.Y(n_5139)
);

AND2x2_ASAP7_75t_L g5140 ( 
.A(n_5038),
.B(n_725),
.Y(n_5140)
);

INVx1_ASAP7_75t_L g5141 ( 
.A(n_5018),
.Y(n_5141)
);

INVx1_ASAP7_75t_L g5142 ( 
.A(n_5018),
.Y(n_5142)
);

INVx1_ASAP7_75t_L g5143 ( 
.A(n_5018),
.Y(n_5143)
);

INVx2_ASAP7_75t_SL g5144 ( 
.A(n_4981),
.Y(n_5144)
);

INVxp67_ASAP7_75t_SL g5145 ( 
.A(n_4981),
.Y(n_5145)
);

NAND2xp5_ASAP7_75t_L g5146 ( 
.A(n_5008),
.B(n_727),
.Y(n_5146)
);

INVx2_ASAP7_75t_L g5147 ( 
.A(n_4981),
.Y(n_5147)
);

INVx1_ASAP7_75t_L g5148 ( 
.A(n_5018),
.Y(n_5148)
);

NAND2xp5_ASAP7_75t_L g5149 ( 
.A(n_5008),
.B(n_728),
.Y(n_5149)
);

INVxp67_ASAP7_75t_L g5150 ( 
.A(n_5131),
.Y(n_5150)
);

BUFx12f_ASAP7_75t_L g5151 ( 
.A(n_5144),
.Y(n_5151)
);

O2A1O1Ixp33_ASAP7_75t_L g5152 ( 
.A1(n_5068),
.A2(n_732),
.B(n_730),
.C(n_731),
.Y(n_5152)
);

OR2x2_ASAP7_75t_L g5153 ( 
.A(n_5070),
.B(n_730),
.Y(n_5153)
);

AND2x2_ASAP7_75t_L g5154 ( 
.A(n_5069),
.B(n_731),
.Y(n_5154)
);

AOI221xp5_ASAP7_75t_L g5155 ( 
.A1(n_5145),
.A2(n_734),
.B1(n_732),
.B2(n_733),
.C(n_735),
.Y(n_5155)
);

INVxp33_ASAP7_75t_L g5156 ( 
.A(n_5123),
.Y(n_5156)
);

AND2x2_ASAP7_75t_L g5157 ( 
.A(n_5066),
.B(n_733),
.Y(n_5157)
);

INVx1_ASAP7_75t_L g5158 ( 
.A(n_5117),
.Y(n_5158)
);

OAI21xp33_ASAP7_75t_SL g5159 ( 
.A1(n_5141),
.A2(n_735),
.B(n_736),
.Y(n_5159)
);

OAI221xp5_ASAP7_75t_L g5160 ( 
.A1(n_5110),
.A2(n_739),
.B1(n_736),
.B2(n_738),
.C(n_740),
.Y(n_5160)
);

NAND2xp5_ASAP7_75t_L g5161 ( 
.A(n_5121),
.B(n_738),
.Y(n_5161)
);

NOR2xp67_ASAP7_75t_L g5162 ( 
.A(n_5142),
.B(n_739),
.Y(n_5162)
);

NAND2xp5_ASAP7_75t_SL g5163 ( 
.A(n_5065),
.B(n_740),
.Y(n_5163)
);

INVx1_ASAP7_75t_L g5164 ( 
.A(n_5117),
.Y(n_5164)
);

XOR2xp5_ASAP7_75t_L g5165 ( 
.A(n_5082),
.B(n_741),
.Y(n_5165)
);

NOR2xp33_ASAP7_75t_L g5166 ( 
.A(n_5067),
.B(n_5074),
.Y(n_5166)
);

OAI22xp5_ASAP7_75t_L g5167 ( 
.A1(n_5111),
.A2(n_745),
.B1(n_742),
.B2(n_743),
.Y(n_5167)
);

OAI22xp5_ASAP7_75t_L g5168 ( 
.A1(n_5127),
.A2(n_746),
.B1(n_743),
.B2(n_745),
.Y(n_5168)
);

AOI222xp33_ASAP7_75t_L g5169 ( 
.A1(n_5143),
.A2(n_748),
.B1(n_750),
.B2(n_746),
.C1(n_747),
.C2(n_749),
.Y(n_5169)
);

INVx1_ASAP7_75t_L g5170 ( 
.A(n_5148),
.Y(n_5170)
);

NAND2xp5_ASAP7_75t_L g5171 ( 
.A(n_5063),
.B(n_747),
.Y(n_5171)
);

XOR2x2_ASAP7_75t_L g5172 ( 
.A(n_5091),
.B(n_748),
.Y(n_5172)
);

AOI22xp33_ASAP7_75t_L g5173 ( 
.A1(n_5118),
.A2(n_752),
.B1(n_749),
.B2(n_751),
.Y(n_5173)
);

NOR2x1_ASAP7_75t_L g5174 ( 
.A(n_5093),
.B(n_751),
.Y(n_5174)
);

INVxp67_ASAP7_75t_L g5175 ( 
.A(n_5073),
.Y(n_5175)
);

CKINVDCx6p67_ASAP7_75t_R g5176 ( 
.A(n_5072),
.Y(n_5176)
);

NAND2xp5_ASAP7_75t_L g5177 ( 
.A(n_5101),
.B(n_752),
.Y(n_5177)
);

INVxp67_ASAP7_75t_L g5178 ( 
.A(n_5116),
.Y(n_5178)
);

OR2x2_ASAP7_75t_L g5179 ( 
.A(n_5064),
.B(n_753),
.Y(n_5179)
);

NAND2xp5_ASAP7_75t_L g5180 ( 
.A(n_5120),
.B(n_753),
.Y(n_5180)
);

NAND2xp5_ASAP7_75t_L g5181 ( 
.A(n_5085),
.B(n_754),
.Y(n_5181)
);

AOI221xp5_ASAP7_75t_L g5182 ( 
.A1(n_5134),
.A2(n_756),
.B1(n_754),
.B2(n_755),
.C(n_757),
.Y(n_5182)
);

NAND2xp5_ASAP7_75t_SL g5183 ( 
.A(n_5097),
.B(n_756),
.Y(n_5183)
);

BUFx3_ASAP7_75t_L g5184 ( 
.A(n_5079),
.Y(n_5184)
);

NAND2xp5_ASAP7_75t_L g5185 ( 
.A(n_5080),
.B(n_758),
.Y(n_5185)
);

INVxp67_ASAP7_75t_SL g5186 ( 
.A(n_5078),
.Y(n_5186)
);

AOI22xp33_ASAP7_75t_L g5187 ( 
.A1(n_5147),
.A2(n_5107),
.B1(n_5130),
.B2(n_5086),
.Y(n_5187)
);

INVx2_ASAP7_75t_SL g5188 ( 
.A(n_5088),
.Y(n_5188)
);

NAND2xp5_ASAP7_75t_SL g5189 ( 
.A(n_5071),
.B(n_758),
.Y(n_5189)
);

AND2x2_ASAP7_75t_L g5190 ( 
.A(n_5112),
.B(n_759),
.Y(n_5190)
);

NAND3xp33_ASAP7_75t_L g5191 ( 
.A(n_5109),
.B(n_759),
.C(n_760),
.Y(n_5191)
);

INVx1_ASAP7_75t_L g5192 ( 
.A(n_5146),
.Y(n_5192)
);

INVx2_ASAP7_75t_L g5193 ( 
.A(n_5108),
.Y(n_5193)
);

INVxp67_ASAP7_75t_L g5194 ( 
.A(n_5149),
.Y(n_5194)
);

INVx1_ASAP7_75t_L g5195 ( 
.A(n_5126),
.Y(n_5195)
);

AOI22x1_ASAP7_75t_L g5196 ( 
.A1(n_5098),
.A2(n_764),
.B1(n_761),
.B2(n_762),
.Y(n_5196)
);

NAND2xp5_ASAP7_75t_L g5197 ( 
.A(n_5081),
.B(n_764),
.Y(n_5197)
);

INVx2_ASAP7_75t_L g5198 ( 
.A(n_5108),
.Y(n_5198)
);

AOI211x1_ASAP7_75t_L g5199 ( 
.A1(n_5094),
.A2(n_767),
.B(n_765),
.C(n_766),
.Y(n_5199)
);

XOR2x2_ASAP7_75t_L g5200 ( 
.A(n_5075),
.B(n_765),
.Y(n_5200)
);

AND2x2_ASAP7_75t_L g5201 ( 
.A(n_5083),
.B(n_5084),
.Y(n_5201)
);

INVx1_ASAP7_75t_L g5202 ( 
.A(n_5089),
.Y(n_5202)
);

INVx1_ASAP7_75t_L g5203 ( 
.A(n_5140),
.Y(n_5203)
);

INVx2_ASAP7_75t_L g5204 ( 
.A(n_5115),
.Y(n_5204)
);

INVx2_ASAP7_75t_SL g5205 ( 
.A(n_5077),
.Y(n_5205)
);

A2O1A1Ixp33_ASAP7_75t_L g5206 ( 
.A1(n_5135),
.A2(n_768),
.B(n_766),
.C(n_767),
.Y(n_5206)
);

INVx1_ASAP7_75t_L g5207 ( 
.A(n_5100),
.Y(n_5207)
);

INVx1_ASAP7_75t_L g5208 ( 
.A(n_5106),
.Y(n_5208)
);

INVx1_ASAP7_75t_L g5209 ( 
.A(n_5114),
.Y(n_5209)
);

AND2x2_ASAP7_75t_L g5210 ( 
.A(n_5087),
.B(n_768),
.Y(n_5210)
);

NOR3xp33_ASAP7_75t_L g5211 ( 
.A(n_5090),
.B(n_769),
.C(n_770),
.Y(n_5211)
);

A2O1A1Ixp33_ASAP7_75t_L g5212 ( 
.A1(n_5124),
.A2(n_772),
.B(n_770),
.C(n_771),
.Y(n_5212)
);

INVx1_ASAP7_75t_L g5213 ( 
.A(n_5076),
.Y(n_5213)
);

XOR2x2_ASAP7_75t_L g5214 ( 
.A(n_5095),
.B(n_771),
.Y(n_5214)
);

NAND2xp5_ASAP7_75t_SL g5215 ( 
.A(n_5096),
.B(n_5092),
.Y(n_5215)
);

NAND2xp5_ASAP7_75t_L g5216 ( 
.A(n_5137),
.B(n_772),
.Y(n_5216)
);

INVx1_ASAP7_75t_L g5217 ( 
.A(n_5099),
.Y(n_5217)
);

AOI22xp5_ASAP7_75t_L g5218 ( 
.A1(n_5103),
.A2(n_775),
.B1(n_773),
.B2(n_774),
.Y(n_5218)
);

NOR2x1_ASAP7_75t_L g5219 ( 
.A(n_5136),
.B(n_773),
.Y(n_5219)
);

O2A1O1Ixp33_ASAP7_75t_L g5220 ( 
.A1(n_5133),
.A2(n_776),
.B(n_774),
.C(n_775),
.Y(n_5220)
);

INVx2_ASAP7_75t_L g5221 ( 
.A(n_5104),
.Y(n_5221)
);

OAI211xp5_ASAP7_75t_L g5222 ( 
.A1(n_5122),
.A2(n_778),
.B(n_776),
.C(n_777),
.Y(n_5222)
);

INVx2_ASAP7_75t_SL g5223 ( 
.A(n_5138),
.Y(n_5223)
);

A2O1A1Ixp33_ASAP7_75t_L g5224 ( 
.A1(n_5139),
.A2(n_779),
.B(n_777),
.C(n_778),
.Y(n_5224)
);

INVx2_ASAP7_75t_L g5225 ( 
.A(n_5105),
.Y(n_5225)
);

OAI22xp5_ASAP7_75t_SL g5226 ( 
.A1(n_5119),
.A2(n_781),
.B1(n_779),
.B2(n_780),
.Y(n_5226)
);

NAND2xp5_ASAP7_75t_L g5227 ( 
.A(n_5162),
.B(n_5113),
.Y(n_5227)
);

AO21x1_ASAP7_75t_L g5228 ( 
.A1(n_5158),
.A2(n_5125),
.B(n_5102),
.Y(n_5228)
);

NOR3xp33_ASAP7_75t_SL g5229 ( 
.A(n_5222),
.B(n_5128),
.C(n_5132),
.Y(n_5229)
);

NAND2xp5_ASAP7_75t_L g5230 ( 
.A(n_5164),
.B(n_5129),
.Y(n_5230)
);

INVx1_ASAP7_75t_SL g5231 ( 
.A(n_5190),
.Y(n_5231)
);

INVx2_ASAP7_75t_SL g5232 ( 
.A(n_5151),
.Y(n_5232)
);

NOR3xp33_ASAP7_75t_L g5233 ( 
.A(n_5166),
.B(n_788),
.C(n_780),
.Y(n_5233)
);

NOR3xp33_ASAP7_75t_L g5234 ( 
.A(n_5215),
.B(n_789),
.C(n_781),
.Y(n_5234)
);

NAND2x1_ASAP7_75t_SL g5235 ( 
.A(n_5193),
.B(n_782),
.Y(n_5235)
);

HB1xp67_ASAP7_75t_L g5236 ( 
.A(n_5198),
.Y(n_5236)
);

NOR2x1_ASAP7_75t_L g5237 ( 
.A(n_5153),
.B(n_782),
.Y(n_5237)
);

AOI211xp5_ASAP7_75t_L g5238 ( 
.A1(n_5160),
.A2(n_785),
.B(n_783),
.C(n_784),
.Y(n_5238)
);

INVx1_ASAP7_75t_L g5239 ( 
.A(n_5161),
.Y(n_5239)
);

AOI21xp33_ASAP7_75t_SL g5240 ( 
.A1(n_5150),
.A2(n_785),
.B(n_784),
.Y(n_5240)
);

NAND4xp75_ASAP7_75t_L g5241 ( 
.A(n_5219),
.B(n_5159),
.C(n_5199),
.D(n_5174),
.Y(n_5241)
);

AOI221xp5_ASAP7_75t_L g5242 ( 
.A1(n_5175),
.A2(n_787),
.B1(n_783),
.B2(n_786),
.C(n_788),
.Y(n_5242)
);

NOR3xp33_ASAP7_75t_L g5243 ( 
.A(n_5188),
.B(n_797),
.C(n_787),
.Y(n_5243)
);

NOR3xp33_ASAP7_75t_L g5244 ( 
.A(n_5205),
.B(n_798),
.C(n_790),
.Y(n_5244)
);

NAND4xp75_ASAP7_75t_L g5245 ( 
.A(n_5170),
.B(n_793),
.C(n_791),
.D(n_792),
.Y(n_5245)
);

NAND3xp33_ASAP7_75t_L g5246 ( 
.A(n_5182),
.B(n_792),
.C(n_793),
.Y(n_5246)
);

AOI22xp5_ASAP7_75t_L g5247 ( 
.A1(n_5186),
.A2(n_796),
.B1(n_794),
.B2(n_795),
.Y(n_5247)
);

NAND3xp33_ASAP7_75t_L g5248 ( 
.A(n_5187),
.B(n_794),
.C(n_795),
.Y(n_5248)
);

NOR2x1_ASAP7_75t_L g5249 ( 
.A(n_5224),
.B(n_5184),
.Y(n_5249)
);

INVx1_ASAP7_75t_L g5250 ( 
.A(n_5210),
.Y(n_5250)
);

AOI22xp5_ASAP7_75t_L g5251 ( 
.A1(n_5165),
.A2(n_798),
.B1(n_796),
.B2(n_797),
.Y(n_5251)
);

NAND2xp5_ASAP7_75t_L g5252 ( 
.A(n_5157),
.B(n_799),
.Y(n_5252)
);

AND2x4_ASAP7_75t_L g5253 ( 
.A(n_5154),
.B(n_800),
.Y(n_5253)
);

AOI22xp5_ASAP7_75t_SL g5254 ( 
.A1(n_5156),
.A2(n_805),
.B1(n_806),
.B2(n_804),
.Y(n_5254)
);

NOR4xp25_ASAP7_75t_L g5255 ( 
.A(n_5183),
.B(n_807),
.C(n_802),
.D(n_804),
.Y(n_5255)
);

NAND2xp5_ASAP7_75t_L g5256 ( 
.A(n_5173),
.B(n_5218),
.Y(n_5256)
);

NAND3xp33_ASAP7_75t_L g5257 ( 
.A(n_5211),
.B(n_802),
.C(n_808),
.Y(n_5257)
);

NOR3xp33_ASAP7_75t_SL g5258 ( 
.A(n_5163),
.B(n_809),
.C(n_810),
.Y(n_5258)
);

NOR2xp33_ASAP7_75t_L g5259 ( 
.A(n_5177),
.B(n_810),
.Y(n_5259)
);

NOR2x1_ASAP7_75t_L g5260 ( 
.A(n_5167),
.B(n_811),
.Y(n_5260)
);

NOR2xp67_ASAP7_75t_L g5261 ( 
.A(n_5191),
.B(n_812),
.Y(n_5261)
);

AND2x2_ASAP7_75t_L g5262 ( 
.A(n_5201),
.B(n_5221),
.Y(n_5262)
);

OA22x2_ASAP7_75t_L g5263 ( 
.A1(n_5223),
.A2(n_813),
.B1(n_811),
.B2(n_812),
.Y(n_5263)
);

NAND3xp33_ASAP7_75t_L g5264 ( 
.A(n_5196),
.B(n_814),
.C(n_815),
.Y(n_5264)
);

NAND4xp25_ASAP7_75t_L g5265 ( 
.A(n_5178),
.B(n_818),
.C(n_815),
.D(n_817),
.Y(n_5265)
);

NOR2x1_ASAP7_75t_L g5266 ( 
.A(n_5180),
.B(n_819),
.Y(n_5266)
);

NOR2x1_ASAP7_75t_L g5267 ( 
.A(n_5179),
.B(n_819),
.Y(n_5267)
);

INVx1_ASAP7_75t_L g5268 ( 
.A(n_5172),
.Y(n_5268)
);

INVx2_ASAP7_75t_L g5269 ( 
.A(n_5200),
.Y(n_5269)
);

NOR3x1_ASAP7_75t_L g5270 ( 
.A(n_5185),
.B(n_5171),
.C(n_5181),
.Y(n_5270)
);

NOR2x1_ASAP7_75t_L g5271 ( 
.A(n_5197),
.B(n_820),
.Y(n_5271)
);

NAND4xp25_ASAP7_75t_L g5272 ( 
.A(n_5208),
.B(n_823),
.C(n_821),
.D(n_822),
.Y(n_5272)
);

NOR2x1_ASAP7_75t_L g5273 ( 
.A(n_5152),
.B(n_821),
.Y(n_5273)
);

NAND3xp33_ASAP7_75t_L g5274 ( 
.A(n_5206),
.B(n_822),
.C(n_823),
.Y(n_5274)
);

INVx6_ASAP7_75t_L g5275 ( 
.A(n_5176),
.Y(n_5275)
);

INVx1_ASAP7_75t_L g5276 ( 
.A(n_5226),
.Y(n_5276)
);

INVx2_ASAP7_75t_L g5277 ( 
.A(n_5203),
.Y(n_5277)
);

NOR2xp33_ASAP7_75t_L g5278 ( 
.A(n_5213),
.B(n_824),
.Y(n_5278)
);

OAI21xp5_ASAP7_75t_SL g5279 ( 
.A1(n_5217),
.A2(n_824),
.B(n_825),
.Y(n_5279)
);

NAND2xp5_ASAP7_75t_L g5280 ( 
.A(n_5169),
.B(n_825),
.Y(n_5280)
);

AO22x2_ASAP7_75t_L g5281 ( 
.A1(n_5195),
.A2(n_828),
.B1(n_826),
.B2(n_827),
.Y(n_5281)
);

NOR3xp33_ASAP7_75t_SL g5282 ( 
.A(n_5189),
.B(n_826),
.C(n_827),
.Y(n_5282)
);

NOR2xp33_ASAP7_75t_L g5283 ( 
.A(n_5265),
.B(n_5216),
.Y(n_5283)
);

NOR2xp33_ASAP7_75t_L g5284 ( 
.A(n_5232),
.B(n_5212),
.Y(n_5284)
);

INVx2_ASAP7_75t_L g5285 ( 
.A(n_5235),
.Y(n_5285)
);

O2A1O1Ixp33_ASAP7_75t_L g5286 ( 
.A1(n_5236),
.A2(n_5220),
.B(n_5225),
.C(n_5194),
.Y(n_5286)
);

OR2x2_ASAP7_75t_L g5287 ( 
.A(n_5255),
.B(n_5204),
.Y(n_5287)
);

INVx2_ASAP7_75t_L g5288 ( 
.A(n_5281),
.Y(n_5288)
);

AOI22xp5_ASAP7_75t_L g5289 ( 
.A1(n_5275),
.A2(n_5214),
.B1(n_5192),
.B2(n_5209),
.Y(n_5289)
);

OAI221xp5_ASAP7_75t_L g5290 ( 
.A1(n_5234),
.A2(n_5202),
.B1(n_5207),
.B2(n_5155),
.C(n_5168),
.Y(n_5290)
);

AOI21xp5_ASAP7_75t_L g5291 ( 
.A1(n_5227),
.A2(n_829),
.B(n_830),
.Y(n_5291)
);

AOI22xp33_ASAP7_75t_L g5292 ( 
.A1(n_5275),
.A2(n_831),
.B1(n_832),
.B2(n_830),
.Y(n_5292)
);

INVx1_ASAP7_75t_L g5293 ( 
.A(n_5263),
.Y(n_5293)
);

INVxp33_ASAP7_75t_SL g5294 ( 
.A(n_5270),
.Y(n_5294)
);

NAND2xp5_ASAP7_75t_L g5295 ( 
.A(n_5253),
.B(n_831),
.Y(n_5295)
);

AOI211xp5_ASAP7_75t_L g5296 ( 
.A1(n_5228),
.A2(n_836),
.B(n_829),
.C(n_835),
.Y(n_5296)
);

OAI211xp5_ASAP7_75t_L g5297 ( 
.A1(n_5238),
.A2(n_838),
.B(n_835),
.C(n_837),
.Y(n_5297)
);

OAI21xp5_ASAP7_75t_SL g5298 ( 
.A1(n_5262),
.A2(n_837),
.B(n_838),
.Y(n_5298)
);

NAND3xp33_ASAP7_75t_L g5299 ( 
.A(n_5233),
.B(n_839),
.C(n_840),
.Y(n_5299)
);

AOI22xp33_ASAP7_75t_SL g5300 ( 
.A1(n_5276),
.A2(n_5231),
.B1(n_5277),
.B2(n_5248),
.Y(n_5300)
);

OAI221xp5_ASAP7_75t_L g5301 ( 
.A1(n_5230),
.A2(n_843),
.B1(n_841),
.B2(n_842),
.C(n_844),
.Y(n_5301)
);

AOI22xp5_ASAP7_75t_L g5302 ( 
.A1(n_5243),
.A2(n_843),
.B1(n_841),
.B2(n_842),
.Y(n_5302)
);

NOR2x1_ASAP7_75t_L g5303 ( 
.A(n_5245),
.B(n_844),
.Y(n_5303)
);

NAND2xp5_ASAP7_75t_L g5304 ( 
.A(n_5253),
.B(n_846),
.Y(n_5304)
);

INVxp67_ASAP7_75t_L g5305 ( 
.A(n_5237),
.Y(n_5305)
);

INVx1_ASAP7_75t_L g5306 ( 
.A(n_5252),
.Y(n_5306)
);

INVx1_ASAP7_75t_L g5307 ( 
.A(n_5267),
.Y(n_5307)
);

NOR2xp33_ASAP7_75t_SL g5308 ( 
.A(n_5241),
.B(n_845),
.Y(n_5308)
);

NAND2xp5_ASAP7_75t_L g5309 ( 
.A(n_5254),
.B(n_848),
.Y(n_5309)
);

XNOR2xp5_ASAP7_75t_L g5310 ( 
.A(n_5229),
.B(n_847),
.Y(n_5310)
);

OAI222xp33_ASAP7_75t_L g5311 ( 
.A1(n_5249),
.A2(n_873),
.B1(n_855),
.B2(n_881),
.C1(n_865),
.C2(n_847),
.Y(n_5311)
);

NOR4xp25_ASAP7_75t_L g5312 ( 
.A(n_5268),
.B(n_850),
.C(n_848),
.D(n_849),
.Y(n_5312)
);

NAND2x1_ASAP7_75t_SL g5313 ( 
.A(n_5266),
.B(n_851),
.Y(n_5313)
);

XNOR2xp5_ASAP7_75t_L g5314 ( 
.A(n_5251),
.B(n_849),
.Y(n_5314)
);

O2A1O1Ixp33_ASAP7_75t_L g5315 ( 
.A1(n_5240),
.A2(n_853),
.B(n_851),
.C(n_852),
.Y(n_5315)
);

NOR2x1p5_ASAP7_75t_L g5316 ( 
.A(n_5264),
.B(n_852),
.Y(n_5316)
);

AOI22xp5_ASAP7_75t_L g5317 ( 
.A1(n_5244),
.A2(n_855),
.B1(n_853),
.B2(n_854),
.Y(n_5317)
);

NOR3x1_ASAP7_75t_L g5318 ( 
.A(n_5298),
.B(n_5257),
.C(n_5297),
.Y(n_5318)
);

NOR4xp25_ASAP7_75t_L g5319 ( 
.A(n_5286),
.B(n_5239),
.C(n_5250),
.D(n_5269),
.Y(n_5319)
);

NOR3xp33_ASAP7_75t_L g5320 ( 
.A(n_5290),
.B(n_5259),
.C(n_5280),
.Y(n_5320)
);

AOI221x1_ASAP7_75t_L g5321 ( 
.A1(n_5307),
.A2(n_5274),
.B1(n_5246),
.B2(n_5278),
.C(n_5256),
.Y(n_5321)
);

AOI21xp5_ASAP7_75t_L g5322 ( 
.A1(n_5305),
.A2(n_5273),
.B(n_5271),
.Y(n_5322)
);

NAND4xp75_ASAP7_75t_L g5323 ( 
.A(n_5303),
.B(n_5260),
.C(n_5261),
.D(n_5258),
.Y(n_5323)
);

NAND2xp5_ASAP7_75t_L g5324 ( 
.A(n_5296),
.B(n_5247),
.Y(n_5324)
);

INVxp67_ASAP7_75t_L g5325 ( 
.A(n_5308),
.Y(n_5325)
);

NOR2xp67_ASAP7_75t_L g5326 ( 
.A(n_5288),
.B(n_5272),
.Y(n_5326)
);

NAND2xp5_ASAP7_75t_L g5327 ( 
.A(n_5312),
.B(n_5279),
.Y(n_5327)
);

INVx1_ASAP7_75t_L g5328 ( 
.A(n_5313),
.Y(n_5328)
);

INVxp67_ASAP7_75t_L g5329 ( 
.A(n_5295),
.Y(n_5329)
);

AND2x4_ASAP7_75t_L g5330 ( 
.A(n_5285),
.B(n_5282),
.Y(n_5330)
);

NOR2x1_ASAP7_75t_L g5331 ( 
.A(n_5311),
.B(n_5281),
.Y(n_5331)
);

NOR3xp33_ASAP7_75t_L g5332 ( 
.A(n_5300),
.B(n_5242),
.C(n_857),
.Y(n_5332)
);

NAND2x1_ASAP7_75t_L g5333 ( 
.A(n_5293),
.B(n_854),
.Y(n_5333)
);

OAI211xp5_ASAP7_75t_SL g5334 ( 
.A1(n_5289),
.A2(n_859),
.B(n_856),
.C(n_857),
.Y(n_5334)
);

NOR3xp33_ASAP7_75t_L g5335 ( 
.A(n_5284),
.B(n_5283),
.C(n_5304),
.Y(n_5335)
);

OAI21xp5_ASAP7_75t_L g5336 ( 
.A1(n_5331),
.A2(n_5310),
.B(n_5294),
.Y(n_5336)
);

NOR3xp33_ASAP7_75t_L g5337 ( 
.A(n_5325),
.B(n_5287),
.C(n_5306),
.Y(n_5337)
);

INVxp67_ASAP7_75t_SL g5338 ( 
.A(n_5333),
.Y(n_5338)
);

OAI21x1_ASAP7_75t_L g5339 ( 
.A1(n_5322),
.A2(n_5291),
.B(n_5315),
.Y(n_5339)
);

AOI22xp5_ASAP7_75t_L g5340 ( 
.A1(n_5326),
.A2(n_5316),
.B1(n_5299),
.B2(n_5302),
.Y(n_5340)
);

HB1xp67_ASAP7_75t_L g5341 ( 
.A(n_5328),
.Y(n_5341)
);

NAND4xp25_ASAP7_75t_L g5342 ( 
.A(n_5321),
.B(n_5309),
.C(n_5317),
.D(n_5301),
.Y(n_5342)
);

OAI22xp33_ASAP7_75t_L g5343 ( 
.A1(n_5327),
.A2(n_5314),
.B1(n_5292),
.B2(n_863),
.Y(n_5343)
);

AOI22x1_ASAP7_75t_L g5344 ( 
.A1(n_5330),
.A2(n_863),
.B1(n_860),
.B2(n_861),
.Y(n_5344)
);

AOI221xp5_ASAP7_75t_L g5345 ( 
.A1(n_5319),
.A2(n_864),
.B1(n_860),
.B2(n_861),
.C(n_865),
.Y(n_5345)
);

OAI22xp5_ASAP7_75t_L g5346 ( 
.A1(n_5324),
.A2(n_867),
.B1(n_864),
.B2(n_866),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_5338),
.Y(n_5347)
);

OR2x2_ASAP7_75t_L g5348 ( 
.A(n_5342),
.B(n_5330),
.Y(n_5348)
);

NAND5xp2_ASAP7_75t_L g5349 ( 
.A(n_5336),
.B(n_5337),
.C(n_5335),
.D(n_5320),
.E(n_5332),
.Y(n_5349)
);

CKINVDCx5p33_ASAP7_75t_R g5350 ( 
.A(n_5341),
.Y(n_5350)
);

INVx1_ASAP7_75t_L g5351 ( 
.A(n_5339),
.Y(n_5351)
);

NOR4xp75_ASAP7_75t_SL g5352 ( 
.A(n_5346),
.B(n_5323),
.C(n_5318),
.D(n_5329),
.Y(n_5352)
);

NOR2xp67_ASAP7_75t_L g5353 ( 
.A(n_5340),
.B(n_5334),
.Y(n_5353)
);

AOI21xp33_ASAP7_75t_SL g5354 ( 
.A1(n_5347),
.A2(n_5343),
.B(n_5344),
.Y(n_5354)
);

OAI22x1_ASAP7_75t_L g5355 ( 
.A1(n_5350),
.A2(n_5345),
.B1(n_868),
.B2(n_866),
.Y(n_5355)
);

AOI21xp5_ASAP7_75t_L g5356 ( 
.A1(n_5351),
.A2(n_867),
.B(n_868),
.Y(n_5356)
);

NOR3xp33_ASAP7_75t_L g5357 ( 
.A(n_5349),
.B(n_869),
.C(n_870),
.Y(n_5357)
);

NOR3xp33_ASAP7_75t_L g5358 ( 
.A(n_5348),
.B(n_870),
.C(n_871),
.Y(n_5358)
);

AND4x1_ASAP7_75t_L g5359 ( 
.A(n_5357),
.B(n_5352),
.C(n_5353),
.D(n_874),
.Y(n_5359)
);

NOR2xp33_ASAP7_75t_L g5360 ( 
.A(n_5354),
.B(n_871),
.Y(n_5360)
);

OAI222xp33_ASAP7_75t_L g5361 ( 
.A1(n_5360),
.A2(n_5356),
.B1(n_5355),
.B2(n_5358),
.C1(n_876),
.C2(n_878),
.Y(n_5361)
);

INVx3_ASAP7_75t_SL g5362 ( 
.A(n_5361),
.Y(n_5362)
);

INVx2_ASAP7_75t_L g5363 ( 
.A(n_5362),
.Y(n_5363)
);

INVx1_ASAP7_75t_SL g5364 ( 
.A(n_5363),
.Y(n_5364)
);

NOR3xp33_ASAP7_75t_SL g5365 ( 
.A(n_5364),
.B(n_5359),
.C(n_872),
.Y(n_5365)
);

OAI222xp33_ASAP7_75t_L g5366 ( 
.A1(n_5365),
.A2(n_879),
.B1(n_881),
.B2(n_875),
.C1(n_877),
.C2(n_880),
.Y(n_5366)
);

AOI21xp5_ASAP7_75t_L g5367 ( 
.A1(n_5366),
.A2(n_875),
.B(n_877),
.Y(n_5367)
);

AOI22xp5_ASAP7_75t_SL g5368 ( 
.A1(n_5367),
.A2(n_883),
.B1(n_880),
.B2(n_882),
.Y(n_5368)
);

HB1xp67_ASAP7_75t_L g5369 ( 
.A(n_5368),
.Y(n_5369)
);

OR2x6_ASAP7_75t_L g5370 ( 
.A(n_5369),
.B(n_882),
.Y(n_5370)
);

AOI21xp5_ASAP7_75t_L g5371 ( 
.A1(n_5370),
.A2(n_883),
.B(n_884),
.Y(n_5371)
);

AOI211xp5_ASAP7_75t_L g5372 ( 
.A1(n_5371),
.A2(n_887),
.B(n_885),
.C(n_886),
.Y(n_5372)
);


endmodule