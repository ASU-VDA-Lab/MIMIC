module fake_jpeg_7928_n_52 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_52);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_52;

wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_32;

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_5),
.Y(n_22)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_15),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_30),
.B(n_32),
.Y(n_36)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_14),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_3),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_3),
.C(n_4),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_4),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_42),
.B(n_43),
.Y(n_47)
);

OA21x2_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_24),
.B(n_25),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_17),
.B(n_18),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_39),
.B1(n_19),
.B2(n_20),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_30),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_41),
.Y(n_44)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_46),
.B(n_35),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_35),
.C(n_36),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_49),
.Y(n_50)
);

MAJx2_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_44),
.C(n_45),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_51),
.B(n_37),
.Y(n_52)
);


endmodule