module fake_jpeg_12442_n_139 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_8),
.B(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_30),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

AOI21xp33_ASAP7_75t_SL g32 ( 
.A1(n_20),
.A2(n_1),
.B(n_2),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_12),
.C(n_13),
.Y(n_58)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_41),
.Y(n_63)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_11),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_37),
.B(n_38),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_14),
.B(n_7),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_3),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_15),
.A2(n_4),
.B(n_7),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_43),
.A2(n_49),
.B(n_28),
.C(n_44),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx2_ASAP7_75t_R g65 ( 
.A(n_44),
.Y(n_65)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_60)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_23),
.B(n_4),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_32),
.B1(n_14),
.B2(n_37),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_24),
.B(n_10),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

CKINVDCx12_ASAP7_75t_R g66 ( 
.A(n_50),
.Y(n_66)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_22),
.B1(n_15),
.B2(n_13),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_59),
.B1(n_62),
.B2(n_69),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_58),
.B(n_75),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_17),
.B1(n_26),
.B2(n_39),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_17),
.B1(n_26),
.B2(n_52),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_35),
.A2(n_34),
.B(n_51),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_40),
.A2(n_29),
.B1(n_31),
.B2(n_36),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_33),
.B1(n_47),
.B2(n_42),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_59),
.B1(n_64),
.B2(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_65),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_91),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_83),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_76),
.A2(n_56),
.B1(n_71),
.B2(n_53),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_82),
.B1(n_92),
.B2(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_63),
.Y(n_83)
);

XOR2x2_ASAP7_75t_SL g101 ( 
.A(n_86),
.B(n_87),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_68),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_92),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_88),
.B(n_90),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_85),
.B1(n_97),
.B2(n_84),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_53),
.Y(n_90)
);

BUFx24_ASAP7_75t_SL g91 ( 
.A(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_55),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_73),
.B(n_70),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_57),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_94),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_77),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_96),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_60),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_108),
.B1(n_109),
.B2(n_107),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_89),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_106),
.B(n_107),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_85),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_84),
.B1(n_79),
.B2(n_78),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_82),
.C(n_87),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_101),
.C(n_104),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_103),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_112),
.B(n_113),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_111),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_116),
.A2(n_108),
.B1(n_109),
.B2(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_102),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_117),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_104),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_118),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_112),
.B1(n_105),
.B2(n_116),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_115),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_129),
.A2(n_131),
.B1(n_121),
.B2(n_105),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_114),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_128),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_133),
.B(n_126),
.Y(n_134)
);

NOR2xp67_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_135),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_136),
.B(n_133),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_121),
.C(n_127),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_138),
.A2(n_135),
.B(n_124),
.Y(n_139)
);


endmodule