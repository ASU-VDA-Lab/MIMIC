module fake_ariane_1585_n_879 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_879);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_879;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_695;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_586;
wire n_443;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_349;
wire n_391;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_857;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_761;
wire n_733;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_495;
wire n_267;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_600;
wire n_481;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_218;
wire n_839;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_369;
wire n_240;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_644;
wire n_536;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_654;
wire n_455;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_612;
wire n_449;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_371;
wire n_845;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_519;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_184;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g181 ( 
.A(n_132),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_99),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_151),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_105),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_74),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_10),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_145),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_1),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_75),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_169),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_129),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_33),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_94),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_139),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_68),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_140),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_34),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_89),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_31),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_109),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_51),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_64),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_13),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_159),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_113),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_131),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_97),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_162),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_170),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_50),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_134),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_146),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_9),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_82),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_32),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_174),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_125),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_156),
.Y(n_219)
);

BUFx10_ASAP7_75t_L g220 ( 
.A(n_13),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_59),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_39),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_158),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_76),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_22),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_103),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_18),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_61),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_101),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_19),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_44),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_52),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_22),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_23),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_37),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_149),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_21),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_25),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_36),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_65),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_171),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_26),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_47),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_130),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_175),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_168),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_3),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_80),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_56),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_91),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_135),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_58),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_178),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_0),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_208),
.Y(n_255)
);

BUFx8_ASAP7_75t_SL g256 ( 
.A(n_224),
.Y(n_256)
);

AND2x6_ASAP7_75t_L g257 ( 
.A(n_193),
.B(n_27),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_181),
.B(n_0),
.Y(n_258)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_208),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_188),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_201),
.Y(n_261)
);

AND2x4_ASAP7_75t_L g262 ( 
.A(n_201),
.B(n_1),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_218),
.B(n_2),
.Y(n_263)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_208),
.Y(n_264)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_208),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_218),
.B(n_2),
.Y(n_266)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_235),
.Y(n_267)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_235),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_193),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_184),
.B(n_3),
.Y(n_270)
);

AND2x4_ASAP7_75t_L g271 ( 
.A(n_211),
.B(n_4),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_204),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_195),
.B(n_4),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_211),
.Y(n_274)
);

AND2x4_ASAP7_75t_L g275 ( 
.A(n_186),
.B(n_5),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_214),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_196),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_199),
.Y(n_278)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_213),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_227),
.Y(n_280)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_236),
.Y(n_281)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_236),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_185),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_220),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_225),
.Y(n_285)
);

BUFx8_ASAP7_75t_L g286 ( 
.A(n_200),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_220),
.Y(n_287)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_220),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_203),
.B(n_212),
.Y(n_289)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_182),
.Y(n_290)
);

BUFx12f_ASAP7_75t_L g291 ( 
.A(n_185),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_230),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_237),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_233),
.Y(n_294)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_252),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_234),
.B(n_5),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_215),
.B(n_223),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_229),
.B(n_6),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_231),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_239),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_245),
.B(n_6),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_251),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_238),
.B(n_247),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_252),
.B(n_7),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_183),
.B(n_7),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_187),
.B(n_8),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_254),
.A2(n_202),
.B1(n_207),
.B2(n_240),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_L g308 ( 
.A1(n_287),
.A2(n_224),
.B1(n_243),
.B2(n_249),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_269),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_263),
.A2(n_243),
.B1(n_250),
.B2(n_248),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_189),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_283),
.B(n_190),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_284),
.B(n_191),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_269),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_285),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_263),
.A2(n_253),
.B1(n_246),
.B2(n_242),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_285),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_266),
.A2(n_241),
.B1(n_232),
.B2(n_228),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_269),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_284),
.B(n_192),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_284),
.B(n_194),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_294),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_266),
.A2(n_226),
.B1(n_222),
.B2(n_221),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_287),
.A2(n_219),
.B1(n_217),
.B2(n_216),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_284),
.B(n_197),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_280),
.B(n_8),
.Y(n_326)
);

OA22x2_ASAP7_75t_L g327 ( 
.A1(n_260),
.A2(n_210),
.B1(n_209),
.B2(n_206),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_271),
.A2(n_205),
.B1(n_198),
.B2(n_11),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_280),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_271),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_288),
.A2(n_293),
.B1(n_292),
.B2(n_272),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_L g332 ( 
.A1(n_288),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_271),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_333)
);

NAND3x1_ASAP7_75t_L g334 ( 
.A(n_273),
.B(n_16),
.C(n_17),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_269),
.Y(n_335)
);

AO22x2_ASAP7_75t_L g336 ( 
.A1(n_262),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_336)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_281),
.Y(n_337)
);

CKINVDCx6p67_ASAP7_75t_R g338 ( 
.A(n_291),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_288),
.B(n_19),
.Y(n_339)
);

OR2x6_ASAP7_75t_L g340 ( 
.A(n_291),
.B(n_20),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_262),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_288),
.B(n_24),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_262),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_288),
.B(n_180),
.Y(n_344)
);

NAND2xp33_ASAP7_75t_SL g345 ( 
.A(n_304),
.B(n_29),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_304),
.A2(n_30),
.B1(n_35),
.B2(n_38),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_L g347 ( 
.A1(n_279),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_289),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_294),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_261),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_303),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_L g352 ( 
.A1(n_279),
.A2(n_48),
.B1(n_49),
.B2(n_53),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_L g353 ( 
.A1(n_279),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_269),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_274),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_256),
.B(n_60),
.Y(n_356)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_281),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_256),
.Y(n_358)
);

OAI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_301),
.A2(n_298),
.B1(n_258),
.B2(n_270),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_309),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_315),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_351),
.B(n_278),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_314),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_329),
.B(n_303),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_317),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_322),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_359),
.A2(n_306),
.B(n_305),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_319),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_349),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_335),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_350),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_354),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_358),
.B(n_261),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_308),
.B(n_356),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_355),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_338),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_339),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_310),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_337),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_337),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_342),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_357),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_326),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_331),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_311),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_313),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_318),
.B(n_278),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_318),
.B(n_299),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_320),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_312),
.B(n_279),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_321),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_325),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_341),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_357),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_316),
.B(n_279),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_344),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_343),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_343),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_328),
.B(n_299),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_323),
.B(n_281),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_328),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_345),
.A2(n_297),
.B(n_290),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_327),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_340),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_340),
.B(n_283),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_330),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_330),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_307),
.B(n_281),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_340),
.B(n_283),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_333),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_348),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_333),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_336),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_336),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_346),
.B(n_295),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_346),
.Y(n_416)
);

INVxp33_ASAP7_75t_L g417 ( 
.A(n_324),
.Y(n_417)
);

BUFx6f_ASAP7_75t_SL g418 ( 
.A(n_334),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_332),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_348),
.Y(n_420)
);

INVx2_ASAP7_75t_SL g421 ( 
.A(n_347),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_352),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_353),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_338),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_312),
.B(n_295),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_315),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_309),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_315),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_315),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_312),
.B(n_295),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_315),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_416),
.B(n_286),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_363),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_363),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_401),
.B(n_406),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_425),
.B(n_275),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_427),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_362),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_427),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_387),
.B(n_275),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_362),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_364),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_372),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_430),
.Y(n_444)
);

NAND2x1p5_ASAP7_75t_L g445 ( 
.A(n_411),
.B(n_275),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_424),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_375),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_361),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_413),
.B(n_296),
.Y(n_449)
);

BUFx4_ASAP7_75t_SL g450 ( 
.A(n_424),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_373),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_387),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_388),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_388),
.B(n_296),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_376),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_365),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_399),
.B(n_415),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_396),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_396),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_399),
.B(n_277),
.Y(n_460)
);

INVxp33_ASAP7_75t_L g461 ( 
.A(n_405),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_421),
.B(n_281),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_396),
.Y(n_463)
);

INVx3_ASAP7_75t_SL g464 ( 
.A(n_378),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_430),
.B(n_286),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_367),
.A2(n_257),
.B(n_300),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_366),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_369),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_396),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_385),
.A2(n_257),
.B(n_300),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_411),
.B(n_277),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_407),
.B(n_276),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_426),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_360),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_386),
.B(n_286),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_410),
.B(n_276),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_360),
.Y(n_477)
);

AND2x2_ASAP7_75t_SL g478 ( 
.A(n_420),
.B(n_268),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_360),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_389),
.B(n_268),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_360),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_391),
.B(n_268),
.Y(n_482)
);

CKINVDCx6p67_ASAP7_75t_R g483 ( 
.A(n_378),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_368),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_409),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_392),
.B(n_282),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_428),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_412),
.B(n_276),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_397),
.B(n_398),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_414),
.B(n_300),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_402),
.A2(n_302),
.B(n_257),
.Y(n_491)
);

AND2x2_ASAP7_75t_SL g492 ( 
.A(n_422),
.B(n_302),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_429),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_383),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_368),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_408),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_379),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_421),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_395),
.B(n_282),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_431),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_371),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_368),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_368),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_370),
.Y(n_504)
);

AND2x6_ASAP7_75t_L g505 ( 
.A(n_489),
.B(n_440),
.Y(n_505)
);

INVx6_ASAP7_75t_L g506 ( 
.A(n_458),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_446),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_444),
.B(n_498),
.Y(n_508)
);

OR2x6_ASAP7_75t_L g509 ( 
.A(n_435),
.B(n_404),
.Y(n_509)
);

INVxp67_ASAP7_75t_SL g510 ( 
.A(n_457),
.Y(n_510)
);

BUFx6f_ASAP7_75t_SL g511 ( 
.A(n_450),
.Y(n_511)
);

INVx5_ASAP7_75t_L g512 ( 
.A(n_458),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_457),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_458),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_441),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_478),
.B(n_423),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_434),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_500),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_479),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_478),
.B(n_377),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_471),
.B(n_381),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_479),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_446),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_434),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_500),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_454),
.B(n_460),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_461),
.B(n_485),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_454),
.B(n_374),
.Y(n_528)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_464),
.B(n_419),
.Y(n_529)
);

OR2x6_ASAP7_75t_L g530 ( 
.A(n_435),
.B(n_393),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_489),
.B(n_403),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_448),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_479),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_487),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_464),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_439),
.Y(n_536)
);

INVx5_ASAP7_75t_L g537 ( 
.A(n_479),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_460),
.B(n_384),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_471),
.B(n_492),
.Y(n_539)
);

INVx8_ASAP7_75t_L g540 ( 
.A(n_490),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_492),
.B(n_395),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_432),
.B(n_418),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_438),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_440),
.B(n_417),
.Y(n_544)
);

AO21x2_ASAP7_75t_L g545 ( 
.A1(n_466),
.A2(n_400),
.B(n_390),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_439),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_479),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_483),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_495),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_452),
.B(n_417),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_495),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_453),
.Y(n_552)
);

OR2x2_ASAP7_75t_L g553 ( 
.A(n_442),
.B(n_302),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_495),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_442),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_501),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_483),
.B(n_384),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_433),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_494),
.B(n_267),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_436),
.B(n_390),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_SL g561 ( 
.A(n_465),
.B(n_418),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_445),
.B(n_379),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_445),
.B(n_380),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_510),
.B(n_472),
.Y(n_564)
);

INVx6_ASAP7_75t_SL g565 ( 
.A(n_509),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_540),
.Y(n_566)
);

BUFx12f_ASAP7_75t_L g567 ( 
.A(n_507),
.Y(n_567)
);

BUFx2_ASAP7_75t_R g568 ( 
.A(n_535),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_528),
.B(n_461),
.Y(n_569)
);

INVxp67_ASAP7_75t_SL g570 ( 
.A(n_510),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_558),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_544),
.B(n_472),
.Y(n_572)
);

INVx3_ASAP7_75t_SL g573 ( 
.A(n_523),
.Y(n_573)
);

BUFx2_ASAP7_75t_SL g574 ( 
.A(n_511),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_548),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_518),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_525),
.Y(n_577)
);

INVxp67_ASAP7_75t_SL g578 ( 
.A(n_522),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_509),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_540),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_515),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_509),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_532),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_515),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_543),
.Y(n_585)
);

BUFx2_ASAP7_75t_R g586 ( 
.A(n_541),
.Y(n_586)
);

INVx6_ASAP7_75t_SL g587 ( 
.A(n_530),
.Y(n_587)
);

BUFx5_ASAP7_75t_L g588 ( 
.A(n_505),
.Y(n_588)
);

BUFx8_ASAP7_75t_SL g589 ( 
.A(n_511),
.Y(n_589)
);

BUFx2_ASAP7_75t_R g590 ( 
.A(n_541),
.Y(n_590)
);

INVx5_ASAP7_75t_L g591 ( 
.A(n_540),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_530),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_534),
.Y(n_593)
);

INVx5_ASAP7_75t_L g594 ( 
.A(n_530),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_531),
.Y(n_595)
);

NAND2x1p5_ASAP7_75t_L g596 ( 
.A(n_512),
.B(n_459),
.Y(n_596)
);

INVx5_ASAP7_75t_L g597 ( 
.A(n_505),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_556),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_531),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_521),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_521),
.Y(n_601)
);

OAI22xp33_ASAP7_75t_L g602 ( 
.A1(n_508),
.A2(n_445),
.B1(n_456),
.B2(n_467),
.Y(n_602)
);

BUFx5_ASAP7_75t_L g603 ( 
.A(n_505),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_522),
.Y(n_604)
);

NAND2x1p5_ASAP7_75t_L g605 ( 
.A(n_512),
.B(n_459),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_526),
.Y(n_606)
);

INVx5_ASAP7_75t_L g607 ( 
.A(n_505),
.Y(n_607)
);

CKINVDCx11_ASAP7_75t_R g608 ( 
.A(n_552),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_517),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_529),
.Y(n_610)
);

NAND2x1p5_ASAP7_75t_L g611 ( 
.A(n_512),
.B(n_469),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_552),
.Y(n_612)
);

NAND2x1p5_ASAP7_75t_L g613 ( 
.A(n_512),
.B(n_469),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_506),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_583),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_593),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_600),
.B(n_601),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_598),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_576),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_572),
.B(n_513),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_577),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_597),
.Y(n_622)
);

BUFx4f_ASAP7_75t_SL g623 ( 
.A(n_567),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_569),
.A2(n_538),
.B1(n_550),
.B2(n_505),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_610),
.A2(n_538),
.B1(n_557),
.B2(n_542),
.Y(n_625)
);

BUFx4f_ASAP7_75t_SL g626 ( 
.A(n_565),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_609),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_570),
.A2(n_508),
.B1(n_513),
.B2(n_520),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_608),
.B(n_418),
.Y(n_629)
);

INVx4_ASAP7_75t_L g630 ( 
.A(n_597),
.Y(n_630)
);

BUFx12f_ASAP7_75t_L g631 ( 
.A(n_579),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_571),
.Y(n_632)
);

BUFx8_ASAP7_75t_L g633 ( 
.A(n_566),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_606),
.Y(n_634)
);

BUFx12f_ASAP7_75t_L g635 ( 
.A(n_582),
.Y(n_635)
);

BUFx4_ASAP7_75t_R g636 ( 
.A(n_588),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_599),
.Y(n_637)
);

CKINVDCx11_ASAP7_75t_R g638 ( 
.A(n_573),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_570),
.A2(n_520),
.B1(n_560),
.B2(n_516),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_589),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_564),
.A2(n_542),
.B1(n_516),
.B2(n_539),
.Y(n_641)
);

CKINVDCx14_ASAP7_75t_R g642 ( 
.A(n_575),
.Y(n_642)
);

CKINVDCx11_ASAP7_75t_R g643 ( 
.A(n_585),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_564),
.Y(n_644)
);

BUFx12f_ASAP7_75t_L g645 ( 
.A(n_566),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_566),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_SL g647 ( 
.A1(n_594),
.A2(n_561),
.B1(n_527),
.B2(n_539),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_597),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_588),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_SL g650 ( 
.A1(n_594),
.A2(n_561),
.B1(n_475),
.B2(n_468),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_587),
.A2(n_451),
.B1(n_493),
.B2(n_473),
.Y(n_651)
);

OAI22xp33_ASAP7_75t_L g652 ( 
.A1(n_607),
.A2(n_612),
.B1(n_595),
.B2(n_467),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_565),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_612),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_587),
.A2(n_468),
.B1(n_473),
.B2(n_493),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_584),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_584),
.A2(n_456),
.B1(n_496),
.B2(n_555),
.Y(n_657)
);

INVx6_ASAP7_75t_L g658 ( 
.A(n_591),
.Y(n_658)
);

OAI21xp33_ASAP7_75t_L g659 ( 
.A1(n_628),
.A2(n_617),
.B(n_620),
.Y(n_659)
);

INVx5_ASAP7_75t_SL g660 ( 
.A(n_640),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_624),
.A2(n_594),
.B1(n_592),
.B2(n_602),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_615),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_645),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_616),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_625),
.A2(n_602),
.B1(n_462),
.B2(n_607),
.Y(n_665)
);

OAI21xp5_ASAP7_75t_SL g666 ( 
.A1(n_650),
.A2(n_568),
.B(n_586),
.Y(n_666)
);

BUFx6f_ASAP7_75t_SL g667 ( 
.A(n_646),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_SL g668 ( 
.A1(n_639),
.A2(n_607),
.B1(n_588),
.B2(n_603),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_620),
.B(n_581),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_618),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_641),
.A2(n_447),
.B1(n_588),
.B2(n_603),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_632),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_619),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_640),
.Y(n_674)
);

AOI22xp5_ASAP7_75t_L g675 ( 
.A1(n_655),
.A2(n_603),
.B1(n_588),
.B2(n_581),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_621),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_647),
.A2(n_447),
.B1(n_603),
.B2(n_443),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_631),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_SL g679 ( 
.A1(n_644),
.A2(n_603),
.B1(n_586),
.B2(n_590),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_632),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_644),
.A2(n_443),
.B1(n_546),
.B2(n_524),
.Y(n_681)
);

OAI21xp33_ASAP7_75t_L g682 ( 
.A1(n_657),
.A2(n_568),
.B(n_482),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_651),
.A2(n_627),
.B1(n_654),
.B2(n_634),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_656),
.A2(n_488),
.B1(n_476),
.B2(n_574),
.Y(n_684)
);

OAI22xp5_ASAP7_75t_L g685 ( 
.A1(n_642),
.A2(n_590),
.B1(n_560),
.B2(n_553),
.Y(n_685)
);

OAI21xp5_ASAP7_75t_SL g686 ( 
.A1(n_629),
.A2(n_455),
.B(n_476),
.Y(n_686)
);

OAI22xp33_ASAP7_75t_L g687 ( 
.A1(n_626),
.A2(n_591),
.B1(n_580),
.B2(n_614),
.Y(n_687)
);

OAI222xp33_ASAP7_75t_L g688 ( 
.A1(n_637),
.A2(n_536),
.B1(n_562),
.B2(n_563),
.C1(n_433),
.C2(n_437),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_SL g689 ( 
.A1(n_631),
.A2(n_499),
.B1(n_545),
.B2(n_488),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_627),
.A2(n_559),
.B1(n_486),
.B2(n_437),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_622),
.Y(n_691)
);

INVx4_ASAP7_75t_L g692 ( 
.A(n_643),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_646),
.B(n_614),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_649),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_633),
.B(n_591),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_SL g696 ( 
.A1(n_635),
.A2(n_545),
.B1(n_470),
.B2(n_463),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_652),
.Y(n_697)
);

OAI21xp5_ASAP7_75t_SL g698 ( 
.A1(n_642),
.A2(n_480),
.B(n_490),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_635),
.A2(n_449),
.B1(n_506),
.B2(n_563),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_648),
.Y(n_700)
);

AOI222xp33_ASAP7_75t_L g701 ( 
.A1(n_623),
.A2(n_449),
.B1(n_490),
.B2(n_257),
.C1(n_562),
.C2(n_274),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_622),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_SL g703 ( 
.A1(n_622),
.A2(n_449),
.B1(n_578),
.B2(n_506),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_645),
.A2(n_580),
.B1(n_514),
.B2(n_605),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_633),
.B(n_578),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_643),
.A2(n_504),
.B1(n_503),
.B2(n_257),
.Y(n_706)
);

OAI21xp33_ASAP7_75t_SL g707 ( 
.A1(n_630),
.A2(n_519),
.B(n_533),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_653),
.A2(n_504),
.B1(n_503),
.B2(n_257),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_649),
.A2(n_484),
.B1(n_477),
.B2(n_514),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_630),
.A2(n_613),
.B1(n_611),
.B2(n_605),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_648),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_630),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_682),
.A2(n_274),
.B1(n_477),
.B2(n_484),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_697),
.A2(n_274),
.B1(n_648),
.B2(n_638),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_665),
.A2(n_274),
.B1(n_638),
.B2(n_502),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_679),
.A2(n_502),
.B1(n_474),
.B2(n_658),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_685),
.A2(n_474),
.B1(n_658),
.B2(n_481),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_689),
.A2(n_474),
.B1(n_658),
.B2(n_481),
.Y(n_718)
);

OAI221xp5_ASAP7_75t_SL g719 ( 
.A1(n_686),
.A2(n_633),
.B1(n_636),
.B2(n_497),
.C(n_491),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_694),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_684),
.A2(n_554),
.B1(n_533),
.B2(n_519),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_659),
.A2(n_481),
.B1(n_370),
.B2(n_495),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_669),
.B(n_662),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_690),
.A2(n_370),
.B1(n_495),
.B2(n_554),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_684),
.A2(n_596),
.B1(n_613),
.B2(n_611),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_664),
.B(n_670),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_683),
.A2(n_370),
.B1(n_549),
.B2(n_551),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_661),
.A2(n_547),
.B1(n_522),
.B2(n_549),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_698),
.A2(n_596),
.B1(n_537),
.B2(n_604),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_SL g730 ( 
.A1(n_666),
.A2(n_636),
.B1(n_604),
.B2(n_267),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_677),
.A2(n_537),
.B1(n_604),
.B2(n_549),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_673),
.B(n_547),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_SL g733 ( 
.A1(n_667),
.A2(n_267),
.B1(n_551),
.B2(n_547),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_701),
.A2(n_551),
.B1(n_267),
.B2(n_537),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_671),
.A2(n_267),
.B1(n_537),
.B2(n_491),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_676),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_680),
.A2(n_282),
.B1(n_255),
.B2(n_290),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_699),
.A2(n_290),
.B1(n_282),
.B2(n_380),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_681),
.A2(n_282),
.B1(n_255),
.B2(n_290),
.Y(n_739)
);

NAND2xp33_ASAP7_75t_SL g740 ( 
.A(n_692),
.B(n_255),
.Y(n_740)
);

AOI222xp33_ASAP7_75t_L g741 ( 
.A1(n_688),
.A2(n_255),
.B1(n_265),
.B2(n_264),
.C1(n_259),
.C2(n_290),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_672),
.A2(n_255),
.B1(n_382),
.B2(n_394),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_693),
.B(n_62),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_696),
.A2(n_394),
.B1(n_382),
.B2(n_265),
.Y(n_744)
);

INVxp67_ASAP7_75t_SL g745 ( 
.A(n_700),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_SL g746 ( 
.A1(n_667),
.A2(n_265),
.B1(n_264),
.B2(n_259),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_668),
.A2(n_265),
.B1(n_264),
.B2(n_259),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_675),
.A2(n_265),
.B1(n_264),
.B2(n_259),
.Y(n_748)
);

OAI221xp5_ASAP7_75t_L g749 ( 
.A1(n_703),
.A2(n_264),
.B1(n_259),
.B2(n_67),
.C(n_69),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_711),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_678),
.A2(n_63),
.B1(n_66),
.B2(n_70),
.Y(n_751)
);

OAI221xp5_ASAP7_75t_L g752 ( 
.A1(n_706),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.C(n_77),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_705),
.B(n_78),
.Y(n_753)
);

NAND3xp33_ASAP7_75t_L g754 ( 
.A(n_719),
.B(n_692),
.C(n_709),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_740),
.B(n_691),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_740),
.B(n_691),
.Y(n_756)
);

OAI221xp5_ASAP7_75t_L g757 ( 
.A1(n_717),
.A2(n_695),
.B1(n_663),
.B2(n_708),
.C(n_704),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_723),
.B(n_702),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_736),
.B(n_745),
.Y(n_759)
);

OAI21xp33_ASAP7_75t_L g760 ( 
.A1(n_750),
.A2(n_712),
.B(n_702),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_720),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_736),
.B(n_712),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_726),
.B(n_660),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_750),
.B(n_660),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_732),
.B(n_663),
.Y(n_765)
);

XNOR2xp5_ASAP7_75t_L g766 ( 
.A(n_730),
.B(n_674),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_720),
.B(n_663),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_753),
.B(n_687),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_721),
.B(n_710),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_721),
.B(n_707),
.Y(n_770)
);

OAI21xp33_ASAP7_75t_L g771 ( 
.A1(n_722),
.A2(n_79),
.B(n_81),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_729),
.B(n_83),
.Y(n_772)
);

OAI21xp5_ASAP7_75t_SL g773 ( 
.A1(n_751),
.A2(n_84),
.B(n_85),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_743),
.B(n_179),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_725),
.B(n_86),
.Y(n_775)
);

AOI21xp33_ASAP7_75t_L g776 ( 
.A1(n_714),
.A2(n_87),
.B(n_88),
.Y(n_776)
);

NAND3xp33_ASAP7_75t_L g777 ( 
.A(n_749),
.B(n_90),
.C(n_92),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_718),
.B(n_177),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_715),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_731),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_728),
.B(n_176),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_SL g782 ( 
.A1(n_716),
.A2(n_98),
.B(n_100),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_727),
.B(n_724),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_744),
.B(n_102),
.Y(n_784)
);

NAND4xp25_ASAP7_75t_L g785 ( 
.A(n_741),
.B(n_173),
.C(n_106),
.D(n_107),
.Y(n_785)
);

NAND3xp33_ASAP7_75t_L g786 ( 
.A(n_752),
.B(n_104),
.C(n_108),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_759),
.B(n_758),
.Y(n_787)
);

OR2x2_ASAP7_75t_L g788 ( 
.A(n_762),
.B(n_748),
.Y(n_788)
);

NAND3xp33_ASAP7_75t_L g789 ( 
.A(n_754),
.B(n_713),
.C(n_747),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_761),
.B(n_735),
.Y(n_790)
);

NAND3xp33_ASAP7_75t_L g791 ( 
.A(n_768),
.B(n_738),
.C(n_734),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_767),
.B(n_764),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_763),
.B(n_733),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_761),
.Y(n_794)
);

AO21x1_ASAP7_75t_SL g795 ( 
.A1(n_770),
.A2(n_737),
.B(n_742),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_785),
.A2(n_746),
.B1(n_739),
.B2(n_112),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_765),
.B(n_110),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_766),
.B(n_111),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_780),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_768),
.B(n_114),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_760),
.B(n_115),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_777),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_802)
);

NAND4xp75_ASAP7_75t_L g803 ( 
.A(n_769),
.B(n_119),
.C(n_120),
.D(n_121),
.Y(n_803)
);

NAND4xp75_ASAP7_75t_L g804 ( 
.A(n_769),
.B(n_122),
.C(n_123),
.D(n_124),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_782),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_805)
);

XOR2x2_ASAP7_75t_L g806 ( 
.A(n_798),
.B(n_772),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_794),
.Y(n_807)
);

NAND4xp75_ASAP7_75t_L g808 ( 
.A(n_800),
.B(n_772),
.C(n_775),
.D(n_774),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_799),
.B(n_755),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_801),
.A2(n_755),
.B(n_756),
.Y(n_810)
);

NOR2x1_ASAP7_75t_R g811 ( 
.A(n_792),
.B(n_756),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_792),
.B(n_783),
.Y(n_812)
);

XOR2xp5_ASAP7_75t_L g813 ( 
.A(n_791),
.B(n_786),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_787),
.B(n_778),
.Y(n_814)
);

NAND4xp75_ASAP7_75t_L g815 ( 
.A(n_805),
.B(n_781),
.C(n_776),
.D(n_784),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_807),
.Y(n_816)
);

XNOR2xp5_ASAP7_75t_L g817 ( 
.A(n_806),
.B(n_787),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_809),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_813),
.B(n_793),
.Y(n_819)
);

XNOR2x2_ASAP7_75t_L g820 ( 
.A(n_808),
.B(n_789),
.Y(n_820)
);

BUFx2_ASAP7_75t_L g821 ( 
.A(n_818),
.Y(n_821)
);

OAI22x1_ASAP7_75t_L g822 ( 
.A1(n_817),
.A2(n_809),
.B1(n_812),
.B2(n_814),
.Y(n_822)
);

OA22x2_ASAP7_75t_L g823 ( 
.A1(n_818),
.A2(n_796),
.B1(n_773),
.B2(n_811),
.Y(n_823)
);

AOI22x1_ASAP7_75t_SL g824 ( 
.A1(n_820),
.A2(n_810),
.B1(n_815),
.B2(n_795),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_821),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_823),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_822),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_824),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_825),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_828),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_830),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_SL g832 ( 
.A1(n_829),
.A2(n_826),
.B1(n_827),
.B2(n_819),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_830),
.Y(n_833)
);

NOR2x1_ASAP7_75t_L g834 ( 
.A(n_833),
.B(n_824),
.Y(n_834)
);

INVxp67_ASAP7_75t_SL g835 ( 
.A(n_832),
.Y(n_835)
);

AOI221xp5_ASAP7_75t_L g836 ( 
.A1(n_831),
.A2(n_810),
.B1(n_802),
.B2(n_816),
.C(n_801),
.Y(n_836)
);

NOR4xp25_ASAP7_75t_L g837 ( 
.A(n_833),
.B(n_802),
.C(n_771),
.D(n_779),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_833),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_833),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_835),
.A2(n_804),
.B1(n_803),
.B2(n_797),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_834),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_838),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_839),
.B(n_788),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_836),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_837),
.B(n_790),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_841),
.Y(n_846)
);

AND3x1_ASAP7_75t_L g847 ( 
.A(n_842),
.B(n_790),
.C(n_757),
.Y(n_847)
);

INVxp67_ASAP7_75t_SL g848 ( 
.A(n_843),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_845),
.Y(n_849)
);

OAI211xp5_ASAP7_75t_SL g850 ( 
.A1(n_844),
.A2(n_133),
.B(n_136),
.C(n_137),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_SL g851 ( 
.A1(n_849),
.A2(n_845),
.B1(n_840),
.B2(n_142),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_848),
.Y(n_852)
);

OAI211xp5_ASAP7_75t_L g853 ( 
.A1(n_846),
.A2(n_138),
.B(n_141),
.C(n_143),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_847),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_850),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_850),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_848),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_849),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_858),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_852),
.B(n_144),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_851),
.A2(n_147),
.B1(n_148),
.B2(n_150),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_854),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_857),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_856),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_855),
.Y(n_865)
);

INVxp67_ASAP7_75t_SL g866 ( 
.A(n_859),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_863),
.Y(n_867)
);

INVxp67_ASAP7_75t_SL g868 ( 
.A(n_860),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_862),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_865),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_870),
.A2(n_864),
.B1(n_866),
.B2(n_868),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_869),
.A2(n_861),
.B1(n_853),
.B2(n_154),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_867),
.A2(n_172),
.B1(n_153),
.B2(n_155),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_871),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_872),
.Y(n_875)
);

OAI22xp33_ASAP7_75t_L g876 ( 
.A1(n_874),
.A2(n_873),
.B1(n_157),
.B2(n_161),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_876),
.Y(n_877)
);

AOI221xp5_ASAP7_75t_L g878 ( 
.A1(n_877),
.A2(n_875),
.B1(n_163),
.B2(n_164),
.C(n_165),
.Y(n_878)
);

AOI211xp5_ASAP7_75t_L g879 ( 
.A1(n_878),
.A2(n_152),
.B(n_166),
.C(n_167),
.Y(n_879)
);


endmodule