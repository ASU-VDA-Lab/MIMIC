module fake_netlist_1_8765_n_921 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_921);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_921;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_911;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_232;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_171;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_769;
wire n_725;
wire n_818;
wire n_844;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_716;
wire n_653;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_522;
wire n_264;
wire n_883;
wire n_200;
wire n_208;
wire n_573;
wire n_898;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_733;
wire n_861;
wire n_899;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_912;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_123;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_223;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_916;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx3_ASAP7_75t_L g111 ( .A(n_67), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_52), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_87), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_45), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_33), .Y(n_115) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_6), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_33), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_98), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_65), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_99), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_95), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_104), .Y(n_122) );
BUFx8_ASAP7_75t_SL g123 ( .A(n_80), .Y(n_123) );
INVx2_ASAP7_75t_SL g124 ( .A(n_27), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_19), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_109), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_36), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_61), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_96), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_85), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_7), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_32), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_23), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_20), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_45), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_90), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_101), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_27), .Y(n_138) );
BUFx3_ASAP7_75t_L g139 ( .A(n_11), .Y(n_139) );
INVx2_ASAP7_75t_SL g140 ( .A(n_110), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_68), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_43), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_7), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_72), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_19), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_0), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_105), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_26), .Y(n_148) );
BUFx10_ASAP7_75t_L g149 ( .A(n_76), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_22), .Y(n_150) );
CKINVDCx14_ASAP7_75t_R g151 ( .A(n_49), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_8), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_16), .Y(n_153) );
BUFx12f_ASAP7_75t_L g154 ( .A(n_149), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_139), .B(n_0), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_111), .Y(n_156) );
BUFx3_ASAP7_75t_L g157 ( .A(n_111), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_124), .B(n_1), .Y(n_158) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_151), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_139), .B(n_1), .Y(n_160) );
INVx2_ASAP7_75t_SL g161 ( .A(n_111), .Y(n_161) );
AND2x2_ASAP7_75t_L g162 ( .A(n_151), .B(n_2), .Y(n_162) );
BUFx2_ASAP7_75t_L g163 ( .A(n_123), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_113), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_139), .Y(n_165) );
BUFx3_ASAP7_75t_L g166 ( .A(n_140), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_124), .B(n_2), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_140), .B(n_3), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_140), .B(n_3), .Y(n_169) );
AND2x6_ASAP7_75t_L g170 ( .A(n_142), .B(n_4), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_116), .B(n_4), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_142), .Y(n_172) );
AND2x6_ASAP7_75t_L g173 ( .A(n_142), .B(n_5), .Y(n_173) );
BUFx12f_ASAP7_75t_L g174 ( .A(n_149), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_124), .B(n_5), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_116), .B(n_6), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_159), .B(n_149), .Y(n_177) );
AND2x2_ASAP7_75t_L g178 ( .A(n_159), .B(n_149), .Y(n_178) );
AO22x2_ASAP7_75t_L g179 ( .A1(n_167), .A2(n_148), .B1(n_150), .B2(n_113), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_159), .B(n_149), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_167), .B(n_150), .Y(n_181) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_171), .A2(n_153), .B1(n_152), .B2(n_114), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_171), .A2(n_153), .B1(n_152), .B2(n_132), .Y(n_183) );
AO22x2_ASAP7_75t_L g184 ( .A1(n_167), .A2(n_148), .B1(n_150), .B2(n_144), .Y(n_184) );
OAI22xp5_ASAP7_75t_SL g185 ( .A1(n_163), .A2(n_131), .B1(n_117), .B2(n_145), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_163), .B(n_119), .Y(n_186) );
OAI22xp33_ASAP7_75t_L g187 ( .A1(n_163), .A2(n_131), .B1(n_117), .B2(n_134), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_171), .A2(n_135), .B1(n_146), .B2(n_127), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_167), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_163), .B(n_119), .Y(n_190) );
NAND3x1_ASAP7_75t_L g191 ( .A(n_171), .B(n_123), .C(n_120), .Y(n_191) );
OAI22xp33_ASAP7_75t_L g192 ( .A1(n_163), .A2(n_115), .B1(n_133), .B2(n_143), .Y(n_192) );
OAI22xp33_ASAP7_75t_SL g193 ( .A1(n_158), .A2(n_125), .B1(n_138), .B2(n_121), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_167), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_171), .A2(n_121), .B1(n_122), .B2(n_118), .Y(n_195) );
AO22x2_ASAP7_75t_L g196 ( .A1(n_167), .A2(n_118), .B1(n_120), .B2(n_136), .Y(n_196) );
OAI22xp33_ASAP7_75t_L g197 ( .A1(n_158), .A2(n_122), .B1(n_144), .B2(n_136), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_176), .A2(n_147), .B1(n_141), .B2(n_137), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_176), .B(n_112), .Y(n_199) );
CKINVDCx6p67_ASAP7_75t_R g200 ( .A(n_154), .Y(n_200) );
BUFx10_ASAP7_75t_L g201 ( .A(n_167), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_165), .Y(n_202) );
NAND3x1_ASAP7_75t_L g203 ( .A(n_176), .B(n_8), .C(n_9), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_165), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_176), .B(n_126), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_176), .A2(n_130), .B1(n_129), .B2(n_128), .Y(n_206) );
OA22x2_ASAP7_75t_L g207 ( .A1(n_167), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_207) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_172), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_154), .B(n_10), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_167), .Y(n_210) );
OAI22xp33_ASAP7_75t_L g211 ( .A1(n_158), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_211) );
INVx2_ASAP7_75t_SL g212 ( .A(n_154), .Y(n_212) );
OAI22xp33_ASAP7_75t_SL g213 ( .A1(n_158), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_213) );
AO22x2_ASAP7_75t_L g214 ( .A1(n_167), .A2(n_15), .B1(n_16), .B2(n_17), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_165), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_155), .Y(n_216) );
OR2x2_ASAP7_75t_L g217 ( .A(n_162), .B(n_15), .Y(n_217) );
OAI22xp33_ASAP7_75t_SL g218 ( .A1(n_175), .A2(n_17), .B1(n_18), .B2(n_20), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_162), .A2(n_18), .B1(n_21), .B2(n_22), .Y(n_219) );
OAI22xp33_ASAP7_75t_L g220 ( .A1(n_164), .A2(n_21), .B1(n_23), .B2(n_24), .Y(n_220) );
OAI22xp33_ASAP7_75t_SL g221 ( .A1(n_175), .A2(n_24), .B1(n_25), .B2(n_26), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_166), .B(n_62), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_216), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_189), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_194), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_210), .Y(n_226) );
OR2x2_ASAP7_75t_SL g227 ( .A(n_217), .B(n_164), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_179), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_179), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_179), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_184), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_184), .Y(n_232) );
INVxp33_ASAP7_75t_L g233 ( .A(n_186), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_184), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_201), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_177), .B(n_154), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_201), .Y(n_237) );
NOR2xp67_ASAP7_75t_L g238 ( .A(n_181), .B(n_154), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_178), .B(n_154), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_201), .Y(n_240) );
INVxp67_ASAP7_75t_SL g241 ( .A(n_181), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_181), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_207), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_207), .Y(n_244) );
BUFx2_ASAP7_75t_L g245 ( .A(n_196), .Y(n_245) );
BUFx3_ASAP7_75t_L g246 ( .A(n_200), .Y(n_246) );
INVxp67_ASAP7_75t_L g247 ( .A(n_180), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_196), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_196), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_197), .B(n_164), .Y(n_250) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_208), .Y(n_251) );
INVx2_ASAP7_75t_SL g252 ( .A(n_200), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_190), .B(n_162), .Y(n_253) );
INVxp67_ASAP7_75t_SL g254 ( .A(n_212), .Y(n_254) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_202), .A2(n_169), .B(n_168), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_214), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_214), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_214), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_202), .Y(n_259) );
BUFx2_ASAP7_75t_L g260 ( .A(n_199), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_208), .Y(n_261) );
XOR2xp5_ASAP7_75t_L g262 ( .A(n_185), .B(n_162), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_208), .Y(n_263) );
INVx3_ASAP7_75t_L g264 ( .A(n_208), .Y(n_264) );
XOR2xp5_ASAP7_75t_L g265 ( .A(n_187), .B(n_162), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_204), .Y(n_266) );
NAND2xp33_ASAP7_75t_SL g267 ( .A(n_212), .B(n_205), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_204), .Y(n_268) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_203), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_215), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_215), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_219), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_209), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_197), .A2(n_161), .B(n_164), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_195), .B(n_174), .Y(n_275) );
CKINVDCx20_ASAP7_75t_R g276 ( .A(n_182), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_183), .B(n_174), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_222), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_211), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_198), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_206), .B(n_174), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_188), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_211), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_218), .Y(n_284) );
AND2x2_ASAP7_75t_SL g285 ( .A(n_245), .B(n_155), .Y(n_285) );
INVx3_ASAP7_75t_L g286 ( .A(n_235), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_241), .B(n_192), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_241), .B(n_192), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_247), .B(n_233), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_265), .B(n_187), .Y(n_290) );
OAI21xp5_ASAP7_75t_L g291 ( .A1(n_274), .A2(n_222), .B(n_193), .Y(n_291) );
OAI21xp5_ASAP7_75t_L g292 ( .A1(n_274), .A2(n_169), .B(n_168), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_253), .B(n_221), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_245), .B(n_174), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_253), .B(n_191), .Y(n_295) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_248), .B(n_174), .Y(n_296) );
INVx1_ASAP7_75t_SL g297 ( .A(n_246), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_247), .B(n_174), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_253), .B(n_155), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_277), .B(n_155), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_251), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_259), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_224), .Y(n_303) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_251), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_277), .B(n_155), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_259), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_277), .B(n_155), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_265), .B(n_220), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_275), .B(n_155), .Y(n_309) );
OR2x2_ASAP7_75t_L g310 ( .A(n_262), .B(n_220), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_224), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_250), .B(n_191), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_275), .B(n_155), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_225), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_238), .B(n_155), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g316 ( .A(n_248), .B(n_213), .Y(n_316) );
BUFx3_ASAP7_75t_L g317 ( .A(n_246), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_259), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_250), .B(n_155), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_275), .B(n_160), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_246), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_225), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_236), .B(n_239), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_284), .B(n_160), .Y(n_324) );
OAI21xp5_ASAP7_75t_L g325 ( .A1(n_278), .A2(n_168), .B(n_169), .Y(n_325) );
AND2x6_ASAP7_75t_L g326 ( .A(n_249), .B(n_160), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_235), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_284), .B(n_160), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_233), .B(n_175), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_279), .B(n_160), .Y(n_330) );
BUFx3_ASAP7_75t_L g331 ( .A(n_228), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_279), .B(n_160), .Y(n_332) );
OAI21xp5_ASAP7_75t_L g333 ( .A1(n_278), .A2(n_160), .B(n_161), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_226), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_283), .B(n_160), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_326), .Y(n_336) );
OR2x6_ASAP7_75t_L g337 ( .A(n_331), .B(n_249), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_286), .B(n_252), .Y(n_338) );
OR2x6_ASAP7_75t_L g339 ( .A(n_331), .B(n_256), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_303), .B(n_272), .Y(n_340) );
OR2x6_ASAP7_75t_L g341 ( .A(n_331), .B(n_256), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_303), .B(n_272), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_326), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_290), .B(n_260), .Y(n_344) );
NAND2x1p5_ASAP7_75t_L g345 ( .A(n_286), .B(n_228), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_331), .B(n_238), .Y(n_346) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_301), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_309), .B(n_229), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_331), .Y(n_349) );
OR2x6_ASAP7_75t_L g350 ( .A(n_309), .B(n_313), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_303), .Y(n_351) );
BUFx6f_ASAP7_75t_SL g352 ( .A(n_285), .Y(n_352) );
AND2x4_ASAP7_75t_L g353 ( .A(n_286), .B(n_327), .Y(n_353) );
INVx3_ASAP7_75t_L g354 ( .A(n_286), .Y(n_354) );
OR2x6_ASAP7_75t_L g355 ( .A(n_309), .B(n_257), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_309), .B(n_229), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_286), .B(n_237), .Y(n_357) );
AND2x4_ASAP7_75t_L g358 ( .A(n_286), .B(n_237), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_311), .Y(n_359) );
AND2x6_ASAP7_75t_L g360 ( .A(n_294), .B(n_257), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_311), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_311), .B(n_283), .Y(n_362) );
CKINVDCx11_ASAP7_75t_R g363 ( .A(n_297), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_302), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_314), .B(n_243), .Y(n_365) );
AND2x2_ASAP7_75t_SL g366 ( .A(n_285), .B(n_258), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_314), .B(n_243), .Y(n_367) );
INVx1_ASAP7_75t_SL g368 ( .A(n_363), .Y(n_368) );
BUFx2_ASAP7_75t_SL g369 ( .A(n_349), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_364), .Y(n_370) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_352), .A2(n_308), .B1(n_290), .B2(n_310), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_353), .Y(n_372) );
INVx5_ASAP7_75t_L g373 ( .A(n_337), .Y(n_373) );
BUFx2_ASAP7_75t_SL g374 ( .A(n_349), .Y(n_374) );
CKINVDCx20_ASAP7_75t_R g375 ( .A(n_336), .Y(n_375) );
INVx1_ASAP7_75t_SL g376 ( .A(n_364), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_353), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_364), .Y(n_378) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_347), .Y(n_379) );
BUFx2_ASAP7_75t_SL g380 ( .A(n_352), .Y(n_380) );
BUFx8_ASAP7_75t_L g381 ( .A(n_352), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_340), .B(n_314), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_353), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_347), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_351), .Y(n_385) );
BUFx3_ASAP7_75t_L g386 ( .A(n_353), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_353), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_347), .Y(n_388) );
INVx1_ASAP7_75t_SL g389 ( .A(n_357), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_352), .Y(n_390) );
BUFx3_ASAP7_75t_L g391 ( .A(n_336), .Y(n_391) );
INVx4_ASAP7_75t_L g392 ( .A(n_337), .Y(n_392) );
INVx5_ASAP7_75t_L g393 ( .A(n_337), .Y(n_393) );
BUFx8_ASAP7_75t_L g394 ( .A(n_343), .Y(n_394) );
BUFx5_ASAP7_75t_L g395 ( .A(n_360), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_344), .B(n_290), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_370), .Y(n_397) );
OAI21xp5_ASAP7_75t_SL g398 ( .A1(n_371), .A2(n_290), .B(n_308), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_385), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_396), .A2(n_308), .B1(n_310), .B2(n_269), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_373), .A2(n_308), .B1(n_337), .B2(n_323), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_392), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_368), .Y(n_403) );
AOI22xp33_ASAP7_75t_SL g404 ( .A1(n_380), .A2(n_269), .B1(n_366), .B2(n_360), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_385), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_385), .Y(n_406) );
INVx3_ASAP7_75t_L g407 ( .A(n_373), .Y(n_407) );
BUFx3_ASAP7_75t_L g408 ( .A(n_373), .Y(n_408) );
INVx8_ASAP7_75t_L g409 ( .A(n_373), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_370), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_396), .A2(n_310), .B1(n_323), .B2(n_350), .Y(n_411) );
INVx6_ASAP7_75t_L g412 ( .A(n_381), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_371), .A2(n_310), .B1(n_366), .B2(n_360), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_370), .Y(n_414) );
BUFx12f_ASAP7_75t_L g415 ( .A(n_381), .Y(n_415) );
BUFx4f_ASAP7_75t_SL g416 ( .A(n_368), .Y(n_416) );
BUFx3_ASAP7_75t_L g417 ( .A(n_373), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_378), .Y(n_418) );
OAI21xp5_ASAP7_75t_L g419 ( .A1(n_382), .A2(n_291), .B(n_329), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_378), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_371), .B(n_293), .Y(n_421) );
INVx6_ASAP7_75t_L g422 ( .A(n_381), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_380), .A2(n_366), .B1(n_360), .B2(n_344), .Y(n_423) );
OAI22xp33_ASAP7_75t_L g424 ( .A1(n_373), .A2(n_350), .B1(n_287), .B2(n_288), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_378), .Y(n_425) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_379), .Y(n_426) );
BUFx6f_ASAP7_75t_SL g427 ( .A(n_392), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_376), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_376), .Y(n_429) );
OAI22xp33_ASAP7_75t_L g430 ( .A1(n_373), .A2(n_350), .B1(n_287), .B2(n_288), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_382), .Y(n_431) );
BUFx3_ASAP7_75t_L g432 ( .A(n_373), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_380), .A2(n_360), .B1(n_350), .B2(n_285), .Y(n_433) );
BUFx4f_ASAP7_75t_L g434 ( .A(n_381), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_375), .B(n_293), .Y(n_435) );
BUFx6f_ASAP7_75t_SL g436 ( .A(n_392), .Y(n_436) );
INVx1_ASAP7_75t_SL g437 ( .A(n_369), .Y(n_437) );
INVx6_ASAP7_75t_L g438 ( .A(n_381), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_373), .A2(n_337), .B1(n_341), .B2(n_339), .Y(n_439) );
INVx4_ASAP7_75t_L g440 ( .A(n_373), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_413), .A2(n_401), .B1(n_421), .B2(n_424), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_433), .A2(n_393), .B1(n_392), .B2(n_390), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_398), .B(n_340), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_397), .Y(n_444) );
AOI22xp33_ASAP7_75t_SL g445 ( .A1(n_412), .A2(n_393), .B1(n_392), .B2(n_381), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_430), .A2(n_360), .B1(n_391), .B2(n_350), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_434), .B(n_393), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_399), .Y(n_448) );
AOI22xp33_ASAP7_75t_SL g449 ( .A1(n_412), .A2(n_393), .B1(n_392), .B2(n_395), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_411), .A2(n_360), .B1(n_391), .B2(n_350), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_411), .A2(n_423), .B1(n_400), .B2(n_404), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_434), .A2(n_393), .B1(n_390), .B2(n_375), .Y(n_452) );
INVx2_ASAP7_75t_SL g453 ( .A(n_409), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_410), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_415), .A2(n_360), .B1(n_391), .B2(n_395), .Y(n_455) );
AOI22xp33_ASAP7_75t_SL g456 ( .A1(n_412), .A2(n_393), .B1(n_395), .B2(n_394), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_399), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_405), .Y(n_458) );
INVx4_ASAP7_75t_L g459 ( .A(n_409), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_415), .A2(n_360), .B1(n_391), .B2(n_395), .Y(n_460) );
AOI22xp33_ASAP7_75t_SL g461 ( .A1(n_412), .A2(n_438), .B1(n_422), .B2(n_409), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_398), .B(n_342), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_427), .A2(n_395), .B1(n_343), .B2(n_394), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_397), .B(n_393), .Y(n_464) );
AOI22xp33_ASAP7_75t_SL g465 ( .A1(n_422), .A2(n_393), .B1(n_395), .B2(n_394), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_427), .A2(n_395), .B1(n_394), .B2(n_386), .Y(n_466) );
BUFx3_ASAP7_75t_L g467 ( .A(n_409), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_434), .A2(n_393), .B1(n_337), .B2(n_389), .Y(n_468) );
INVx3_ASAP7_75t_L g469 ( .A(n_426), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_405), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_427), .A2(n_395), .B1(n_394), .B2(n_372), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_397), .B(n_369), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_406), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_406), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_431), .B(n_342), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_414), .Y(n_476) );
AOI22xp33_ASAP7_75t_SL g477 ( .A1(n_422), .A2(n_393), .B1(n_395), .B2(n_394), .Y(n_477) );
AOI22xp33_ASAP7_75t_SL g478 ( .A1(n_422), .A2(n_395), .B1(n_369), .B2(n_374), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_414), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_418), .B(n_374), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_416), .B(n_282), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_436), .A2(n_419), .B1(n_431), .B2(n_438), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_435), .B(n_312), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_418), .B(n_374), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_426), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_420), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_420), .Y(n_487) );
OAI22xp33_ASAP7_75t_L g488 ( .A1(n_438), .A2(n_389), .B1(n_288), .B2(n_287), .Y(n_488) );
AOI22xp33_ASAP7_75t_SL g489 ( .A1(n_438), .A2(n_395), .B1(n_372), .B2(n_387), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_425), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_439), .A2(n_341), .B1(n_339), .B2(n_262), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_425), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_436), .A2(n_395), .B1(n_377), .B2(n_387), .Y(n_493) );
OAI21xp5_ASAP7_75t_SL g494 ( .A1(n_407), .A2(n_305), .B(n_300), .Y(n_494) );
NOR2x1_ASAP7_75t_SL g495 ( .A(n_440), .B(n_339), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_426), .Y(n_496) );
AOI22xp33_ASAP7_75t_SL g497 ( .A1(n_409), .A2(n_395), .B1(n_372), .B2(n_387), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_407), .B(n_312), .Y(n_498) );
AOI222xp33_ASAP7_75t_L g499 ( .A1(n_403), .A2(n_312), .B1(n_295), .B2(n_293), .C1(n_258), .C2(n_307), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_428), .B(n_384), .Y(n_500) );
AOI222xp33_ASAP7_75t_L g501 ( .A1(n_436), .A2(n_295), .B1(n_305), .B2(n_307), .C1(n_300), .C2(n_316), .Y(n_501) );
BUFx12f_ASAP7_75t_L g502 ( .A(n_440), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_440), .A2(n_341), .B1(n_339), .B2(n_203), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_402), .A2(n_395), .B1(n_372), .B2(n_387), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_437), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_402), .A2(n_386), .B1(n_383), .B2(n_377), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_428), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_408), .A2(n_386), .B1(n_383), .B2(n_377), .Y(n_508) );
BUFx6f_ASAP7_75t_SL g509 ( .A(n_408), .Y(n_509) );
OAI22xp33_ASAP7_75t_L g510 ( .A1(n_440), .A2(n_339), .B1(n_341), .B2(n_355), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_408), .A2(n_386), .B1(n_383), .B2(n_377), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_432), .A2(n_383), .B1(n_355), .B2(n_285), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_407), .B(n_321), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_451), .A2(n_432), .B1(n_417), .B2(n_407), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_503), .A2(n_432), .B1(n_417), .B2(n_355), .Y(n_515) );
NOR3xp33_ASAP7_75t_SL g516 ( .A(n_481), .B(n_280), .C(n_295), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_494), .A2(n_417), .B1(n_227), .B2(n_339), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_448), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_443), .A2(n_355), .B1(n_170), .B2(n_173), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_462), .A2(n_355), .B1(n_170), .B2(n_173), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_441), .A2(n_355), .B1(n_170), .B2(n_173), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_501), .A2(n_173), .B1(n_170), .B2(n_291), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_500), .B(n_429), .Y(n_523) );
AOI221xp5_ASAP7_75t_L g524 ( .A1(n_483), .A2(n_289), .B1(n_329), .B2(n_160), .C(n_316), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_501), .A2(n_173), .B1(n_170), .B2(n_291), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_491), .A2(n_173), .B1(n_170), .B2(n_356), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_494), .A2(n_227), .B1(n_341), .B2(n_276), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_450), .A2(n_173), .B1(n_170), .B2(n_356), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_476), .B(n_429), .Y(n_529) );
OAI221xp5_ASAP7_75t_L g530 ( .A1(n_482), .A2(n_289), .B1(n_244), .B2(n_260), .C(n_292), .Y(n_530) );
NAND3xp33_ASAP7_75t_L g531 ( .A(n_454), .B(n_172), .C(n_244), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_476), .B(n_170), .Y(n_532) );
OAI221xp5_ASAP7_75t_L g533 ( .A1(n_499), .A2(n_292), .B1(n_267), .B2(n_307), .C(n_300), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_461), .A2(n_227), .B1(n_341), .B2(n_362), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_445), .A2(n_362), .B1(n_359), .B2(n_361), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_500), .B(n_426), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_456), .A2(n_359), .B1(n_351), .B2(n_361), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_446), .A2(n_173), .B1(n_170), .B2(n_356), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_465), .A2(n_285), .B1(n_346), .B2(n_321), .Y(n_539) );
AOI221xp5_ASAP7_75t_L g540 ( .A1(n_488), .A2(n_160), .B1(n_307), .B2(n_300), .C(n_305), .Y(n_540) );
AOI22xp33_ASAP7_75t_SL g541 ( .A1(n_495), .A2(n_426), .B1(n_305), .B2(n_320), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_512), .A2(n_170), .B1(n_173), .B2(n_348), .Y(n_542) );
OAI221xp5_ASAP7_75t_L g543 ( .A1(n_499), .A2(n_292), .B1(n_267), .B2(n_325), .C(n_313), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_510), .A2(n_170), .B1(n_173), .B2(n_348), .Y(n_544) );
AOI222xp33_ASAP7_75t_L g545 ( .A1(n_502), .A2(n_170), .B1(n_173), .B2(n_324), .C1(n_328), .C2(n_313), .Y(n_545) );
NAND2xp33_ASAP7_75t_SL g546 ( .A(n_459), .B(n_379), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_459), .A2(n_348), .B1(n_320), .B2(n_313), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_479), .B(n_170), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_479), .B(n_170), .Y(n_549) );
OAI22xp5_ASAP7_75t_SL g550 ( .A1(n_502), .A2(n_346), .B1(n_297), .B2(n_384), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_459), .A2(n_170), .B1(n_173), .B2(n_346), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_486), .B(n_170), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_459), .A2(n_170), .B1(n_173), .B2(n_346), .Y(n_553) );
NAND2xp33_ASAP7_75t_SL g554 ( .A(n_509), .B(n_379), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_477), .B(n_379), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_448), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_457), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_509), .A2(n_170), .B1(n_173), .B2(n_346), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_509), .A2(n_170), .B1(n_173), .B2(n_320), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_457), .Y(n_560) );
AOI22xp33_ASAP7_75t_SL g561 ( .A1(n_495), .A2(n_320), .B1(n_388), .B2(n_379), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_455), .A2(n_345), .B1(n_384), .B2(n_297), .Y(n_562) );
OA21x2_ASAP7_75t_L g563 ( .A1(n_485), .A2(n_384), .B(n_333), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_460), .A2(n_345), .B1(n_334), .B2(n_322), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_442), .A2(n_173), .B1(n_315), .B2(n_328), .Y(n_565) );
OAI222xp33_ASAP7_75t_L g566 ( .A1(n_454), .A2(n_345), .B1(n_161), .B2(n_299), .C1(n_281), .C2(n_294), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_466), .A2(n_345), .B1(n_334), .B2(n_322), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_467), .A2(n_464), .B1(n_489), .B2(n_463), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_467), .A2(n_173), .B1(n_315), .B2(n_324), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_467), .A2(n_173), .B1(n_315), .B2(n_324), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_471), .A2(n_322), .B1(n_334), .B2(n_298), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_458), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_497), .A2(n_298), .B1(n_365), .B2(n_367), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_486), .B(n_173), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_464), .A2(n_468), .B1(n_452), .B2(n_449), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_447), .A2(n_388), .B(n_379), .Y(n_576) );
AND2x4_ASAP7_75t_L g577 ( .A(n_444), .B(n_379), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_464), .A2(n_315), .B1(n_324), .B2(n_328), .Y(n_578) );
AOI22xp33_ASAP7_75t_SL g579 ( .A1(n_453), .A2(n_388), .B1(n_379), .B2(n_281), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_478), .B(n_379), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_464), .A2(n_315), .B1(n_328), .B2(n_299), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_487), .B(n_172), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_487), .B(n_172), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_453), .A2(n_315), .B1(n_299), .B2(n_325), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_506), .A2(n_315), .B1(n_299), .B2(n_325), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_475), .A2(n_294), .B1(n_281), .B2(n_365), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_458), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_507), .B(n_156), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_490), .B(n_172), .Y(n_589) );
AOI222xp33_ASAP7_75t_L g590 ( .A1(n_470), .A2(n_367), .B1(n_335), .B2(n_332), .C1(n_330), .C2(n_231), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_490), .B(n_172), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_498), .A2(n_326), .B1(n_172), .B2(n_232), .Y(n_592) );
AOI22xp33_ASAP7_75t_SL g593 ( .A1(n_480), .A2(n_388), .B1(n_317), .B2(n_294), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_508), .A2(n_326), .B1(n_172), .B2(n_232), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_511), .A2(n_326), .B1(n_172), .B2(n_230), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_480), .A2(n_326), .B1(n_172), .B2(n_230), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_484), .A2(n_326), .B1(n_172), .B2(n_231), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_484), .A2(n_326), .B1(n_172), .B2(n_234), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_504), .A2(n_492), .B1(n_473), .B2(n_474), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_513), .A2(n_234), .B1(n_239), .B2(n_236), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_492), .A2(n_326), .B1(n_172), .B2(n_330), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_470), .B(n_172), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_473), .A2(n_326), .B1(n_330), .B2(n_335), .Y(n_603) );
OAI211xp5_ASAP7_75t_SL g604 ( .A1(n_493), .A2(n_332), .B(n_335), .C(n_156), .Y(n_604) );
AOI222xp33_ASAP7_75t_L g605 ( .A1(n_474), .A2(n_332), .B1(n_319), .B2(n_333), .C1(n_161), .C2(n_156), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_505), .A2(n_326), .B1(n_319), .B2(n_388), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_472), .A2(n_388), .B1(n_354), .B2(n_317), .Y(n_607) );
AOI222xp33_ASAP7_75t_L g608 ( .A1(n_507), .A2(n_161), .B1(n_166), .B2(n_319), .C1(n_156), .C2(n_333), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_472), .B(n_25), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_444), .A2(n_326), .B1(n_388), .B2(n_296), .Y(n_610) );
AOI22xp33_ASAP7_75t_SL g611 ( .A1(n_444), .A2(n_388), .B1(n_317), .B2(n_347), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_496), .B(n_388), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_485), .Y(n_613) );
NAND3xp33_ASAP7_75t_L g614 ( .A(n_485), .B(n_156), .C(n_165), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_536), .B(n_496), .Y(n_615) );
AOI22xp5_ASAP7_75t_SL g616 ( .A1(n_527), .A2(n_469), .B1(n_496), .B2(n_317), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_523), .B(n_469), .Y(n_617) );
AOI21xp33_ASAP7_75t_L g618 ( .A1(n_609), .A2(n_534), .B(n_535), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_546), .B(n_469), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_517), .A2(n_469), .B1(n_326), .B2(n_357), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_530), .A2(n_165), .B1(n_161), .B2(n_156), .C(n_166), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_536), .B(n_165), .Y(n_622) );
AOI211xp5_ASAP7_75t_L g623 ( .A1(n_539), .A2(n_165), .B(n_166), .C(n_157), .Y(n_623) );
NOR2xp33_ASAP7_75t_SL g624 ( .A(n_566), .B(n_317), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_523), .B(n_28), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_518), .B(n_165), .Y(n_626) );
NAND4xp25_ASAP7_75t_L g627 ( .A(n_514), .B(n_166), .C(n_157), .D(n_255), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_518), .B(n_165), .Y(n_628) );
NAND3xp33_ASAP7_75t_L g629 ( .A(n_545), .B(n_165), .C(n_166), .Y(n_629) );
OAI221xp5_ASAP7_75t_SL g630 ( .A1(n_568), .A2(n_166), .B1(n_157), .B2(n_242), .C(n_223), .Y(n_630) );
NAND3xp33_ASAP7_75t_L g631 ( .A(n_545), .B(n_165), .C(n_157), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_556), .B(n_28), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_556), .B(n_165), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_557), .B(n_29), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_557), .B(n_29), .Y(n_635) );
NAND3xp33_ASAP7_75t_L g636 ( .A(n_516), .B(n_165), .C(n_157), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_560), .B(n_30), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_522), .A2(n_326), .B1(n_165), .B2(n_296), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_560), .B(n_30), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_572), .B(n_31), .Y(n_640) );
AOI21x1_ASAP7_75t_L g641 ( .A1(n_580), .A2(n_278), .B(n_255), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_572), .B(n_31), .Y(n_642) );
OAI221xp5_ASAP7_75t_L g643 ( .A1(n_541), .A2(n_157), .B1(n_223), .B2(n_242), .C(n_226), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_587), .B(n_32), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_587), .B(n_34), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_613), .B(n_34), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_599), .B(n_35), .Y(n_647) );
OAI221xp5_ASAP7_75t_SL g648 ( .A1(n_525), .A2(n_354), .B1(n_273), .B2(n_306), .C(n_318), .Y(n_648) );
AOI22xp33_ASAP7_75t_SL g649 ( .A1(n_550), .A2(n_347), .B1(n_354), .B2(n_273), .Y(n_649) );
OAI21xp5_ASAP7_75t_L g650 ( .A1(n_531), .A2(n_358), .B(n_357), .Y(n_650) );
OAI21xp5_ASAP7_75t_SL g651 ( .A1(n_561), .A2(n_252), .B(n_357), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_529), .B(n_35), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_613), .B(n_36), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_533), .A2(n_515), .B1(n_543), .B2(n_579), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_582), .B(n_37), .Y(n_655) );
NAND3xp33_ASAP7_75t_L g656 ( .A(n_531), .B(n_347), .C(n_302), .Y(n_656) );
NAND3xp33_ASAP7_75t_L g657 ( .A(n_519), .B(n_347), .C(n_302), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_583), .B(n_37), .Y(n_658) );
NAND2x1_ASAP7_75t_L g659 ( .A(n_575), .B(n_354), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_612), .B(n_38), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_612), .B(n_38), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_589), .B(n_39), .Y(n_662) );
NAND3xp33_ASAP7_75t_L g663 ( .A(n_520), .B(n_306), .C(n_302), .Y(n_663) );
NAND3xp33_ASAP7_75t_L g664 ( .A(n_558), .B(n_306), .C(n_302), .Y(n_664) );
NAND3xp33_ASAP7_75t_L g665 ( .A(n_546), .B(n_306), .C(n_318), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_591), .B(n_39), .Y(n_666) );
OAI21xp5_ASAP7_75t_SL g667 ( .A1(n_537), .A2(n_252), .B(n_358), .Y(n_667) );
NAND4xp25_ASAP7_75t_L g668 ( .A(n_551), .B(n_40), .C(n_41), .D(n_42), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_602), .B(n_40), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_577), .B(n_41), .Y(n_670) );
OAI211xp5_ASAP7_75t_SL g671 ( .A1(n_526), .A2(n_338), .B(n_43), .C(n_44), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g672 ( .A1(n_521), .A2(n_42), .B1(n_44), .B2(n_46), .C(n_47), .Y(n_672) );
NAND3xp33_ASAP7_75t_L g673 ( .A(n_555), .B(n_306), .C(n_318), .Y(n_673) );
NAND4xp25_ASAP7_75t_L g674 ( .A(n_553), .B(n_46), .C(n_47), .D(n_48), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_577), .B(n_48), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_577), .B(n_49), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_577), .B(n_50), .Y(n_677) );
OA21x2_ASAP7_75t_L g678 ( .A1(n_576), .A2(n_318), .B(n_261), .Y(n_678) );
OA211x2_ASAP7_75t_L g679 ( .A1(n_554), .A2(n_50), .B(n_51), .C(n_53), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_532), .B(n_318), .Y(n_680) );
OAI21xp5_ASAP7_75t_SL g681 ( .A1(n_593), .A2(n_358), .B(n_357), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_563), .B(n_54), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g683 ( .A(n_544), .B(n_273), .C(n_358), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_548), .B(n_358), .Y(n_684) );
OAI21xp5_ASAP7_75t_SL g685 ( .A1(n_606), .A2(n_327), .B(n_286), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_550), .A2(n_327), .B1(n_304), .B2(n_301), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_549), .B(n_55), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_552), .B(n_56), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_574), .B(n_57), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_565), .A2(n_327), .B1(n_304), .B2(n_301), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_588), .B(n_58), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g692 ( .A(n_559), .B(n_304), .C(n_301), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_588), .B(n_59), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_563), .B(n_60), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_590), .B(n_63), .Y(n_695) );
NAND3xp33_ASAP7_75t_L g696 ( .A(n_569), .B(n_304), .C(n_301), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_563), .Y(n_697) );
NAND2xp33_ASAP7_75t_SL g698 ( .A(n_562), .B(n_327), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_586), .B(n_64), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_590), .B(n_66), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_547), .A2(n_327), .B1(n_304), .B2(n_301), .Y(n_701) );
OAI22xp33_ASAP7_75t_L g702 ( .A1(n_547), .A2(n_327), .B1(n_304), .B2(n_301), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_563), .B(n_69), .Y(n_703) );
OAI221xp5_ASAP7_75t_L g704 ( .A1(n_528), .A2(n_254), .B1(n_240), .B2(n_271), .C(n_270), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_573), .B(n_70), .Y(n_705) );
OAI221xp5_ASAP7_75t_SL g706 ( .A1(n_538), .A2(n_254), .B1(n_73), .B2(n_74), .C(n_75), .Y(n_706) );
NAND3xp33_ASAP7_75t_L g707 ( .A(n_570), .B(n_304), .C(n_301), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_607), .B(n_71), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_567), .B(n_77), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_585), .B(n_78), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_605), .B(n_79), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_540), .A2(n_604), .B1(n_564), .B2(n_524), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_611), .B(n_81), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_578), .B(n_82), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_605), .B(n_83), .Y(n_715) );
NAND2xp5_ASAP7_75t_SL g716 ( .A(n_554), .B(n_304), .Y(n_716) );
OAI221xp5_ASAP7_75t_L g717 ( .A1(n_542), .A2(n_240), .B1(n_266), .B2(n_271), .C(n_270), .Y(n_717) );
OA21x2_ASAP7_75t_L g718 ( .A1(n_614), .A2(n_263), .B(n_261), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_581), .B(n_84), .Y(n_719) );
AOI211xp5_ASAP7_75t_L g720 ( .A1(n_618), .A2(n_571), .B(n_614), .C(n_600), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_647), .B(n_600), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_622), .Y(n_722) );
AND2x4_ASAP7_75t_L g723 ( .A(n_615), .B(n_610), .Y(n_723) );
NAND3xp33_ASAP7_75t_L g724 ( .A(n_654), .B(n_608), .C(n_603), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_622), .B(n_598), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_615), .B(n_584), .Y(n_726) );
NAND3xp33_ASAP7_75t_L g727 ( .A(n_673), .B(n_601), .C(n_597), .Y(n_727) );
OR2x2_ASAP7_75t_L g728 ( .A(n_617), .B(n_596), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_697), .B(n_595), .Y(n_729) );
AND2x4_ASAP7_75t_SL g730 ( .A(n_670), .B(n_675), .Y(n_730) );
NAND3xp33_ASAP7_75t_SL g731 ( .A(n_624), .B(n_586), .C(n_594), .Y(n_731) );
CKINVDCx5p33_ASAP7_75t_R g732 ( .A(n_660), .Y(n_732) );
NOR3xp33_ASAP7_75t_SL g733 ( .A(n_667), .B(n_592), .C(n_88), .Y(n_733) );
NAND3xp33_ASAP7_75t_SL g734 ( .A(n_651), .B(n_86), .C(n_89), .Y(n_734) );
OR2x2_ASAP7_75t_L g735 ( .A(n_660), .B(n_91), .Y(n_735) );
NAND4xp75_ASAP7_75t_L g736 ( .A(n_679), .B(n_92), .C(n_93), .D(n_94), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_697), .B(n_97), .Y(n_737) );
INVxp67_ASAP7_75t_SL g738 ( .A(n_716), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_625), .B(n_100), .Y(n_739) );
AOI221xp5_ASAP7_75t_L g740 ( .A1(n_652), .A2(n_268), .B1(n_266), .B2(n_263), .C(n_304), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_681), .A2(n_304), .B1(n_301), .B2(n_268), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_661), .B(n_102), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_661), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_626), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_646), .B(n_103), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_628), .Y(n_746) );
NOR2x1_ASAP7_75t_L g747 ( .A(n_665), .B(n_301), .Y(n_747) );
AND2x2_ASAP7_75t_L g748 ( .A(n_670), .B(n_106), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_620), .A2(n_264), .B1(n_108), .B2(n_107), .Y(n_749) );
NAND4xp75_ASAP7_75t_L g750 ( .A(n_679), .B(n_251), .C(n_264), .D(n_675), .Y(n_750) );
BUFx2_ASAP7_75t_L g751 ( .A(n_676), .Y(n_751) );
AND2x2_ASAP7_75t_L g752 ( .A(n_676), .B(n_264), .Y(n_752) );
AND2x2_ASAP7_75t_L g753 ( .A(n_677), .B(n_264), .Y(n_753) );
NAND3xp33_ASAP7_75t_L g754 ( .A(n_623), .B(n_251), .C(n_264), .Y(n_754) );
NAND3xp33_ASAP7_75t_L g755 ( .A(n_659), .B(n_251), .C(n_616), .Y(n_755) );
NAND3xp33_ASAP7_75t_L g756 ( .A(n_659), .B(n_251), .C(n_632), .Y(n_756) );
AND2x4_ASAP7_75t_L g757 ( .A(n_619), .B(n_251), .Y(n_757) );
NAND3xp33_ASAP7_75t_L g758 ( .A(n_634), .B(n_637), .C(n_644), .Y(n_758) );
OAI211xp5_ASAP7_75t_SL g759 ( .A1(n_712), .A2(n_672), .B(n_695), .C(n_700), .Y(n_759) );
OAI21xp33_ASAP7_75t_SL g760 ( .A1(n_716), .A2(n_619), .B(n_677), .Y(n_760) );
OR2x2_ASAP7_75t_L g761 ( .A(n_646), .B(n_653), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_653), .B(n_639), .Y(n_762) );
AND2x4_ASAP7_75t_L g763 ( .A(n_641), .B(n_628), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_639), .B(n_642), .Y(n_764) );
NAND3xp33_ASAP7_75t_L g765 ( .A(n_635), .B(n_640), .C(n_698), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g766 ( .A1(n_620), .A2(n_631), .B1(n_629), .B2(n_698), .Y(n_766) );
NAND4xp75_ASAP7_75t_L g767 ( .A(n_642), .B(n_645), .C(n_705), .D(n_699), .Y(n_767) );
AND2x2_ASAP7_75t_L g768 ( .A(n_641), .B(n_682), .Y(n_768) );
OAI221xp5_ASAP7_75t_SL g769 ( .A1(n_685), .A2(n_715), .B1(n_711), .B2(n_643), .C(n_668), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_633), .Y(n_770) );
OAI21xp5_ASAP7_75t_L g771 ( .A1(n_656), .A2(n_649), .B(n_650), .Y(n_771) );
AOI22xp33_ASAP7_75t_SL g772 ( .A1(n_645), .A2(n_686), .B1(n_694), .B2(n_682), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_694), .B(n_633), .Y(n_773) );
NOR2x1_ASAP7_75t_L g774 ( .A(n_713), .B(n_708), .Y(n_774) );
AO21x2_ASAP7_75t_L g775 ( .A1(n_703), .A2(n_709), .B(n_658), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_708), .B(n_678), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_674), .A2(n_683), .B1(n_671), .B2(n_657), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_678), .B(n_713), .Y(n_778) );
OR2x2_ASAP7_75t_L g779 ( .A(n_680), .B(n_678), .Y(n_779) );
INVx2_ASAP7_75t_SL g780 ( .A(n_718), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_630), .B(n_666), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_718), .B(n_684), .Y(n_782) );
CKINVDCx5p33_ASAP7_75t_R g783 ( .A(n_655), .Y(n_783) );
INVx1_ASAP7_75t_SL g784 ( .A(n_662), .Y(n_784) );
NAND4xp75_ASAP7_75t_L g785 ( .A(n_719), .B(n_714), .C(n_710), .D(n_669), .Y(n_785) );
NAND4xp75_ASAP7_75t_L g786 ( .A(n_719), .B(n_714), .C(n_689), .D(n_688), .Y(n_786) );
OR2x6_ASAP7_75t_L g787 ( .A(n_701), .B(n_707), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_718), .B(n_687), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_691), .B(n_693), .Y(n_789) );
AND2x2_ASAP7_75t_L g790 ( .A(n_690), .B(n_696), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_663), .B(n_692), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_621), .B(n_702), .Y(n_792) );
NAND3xp33_ASAP7_75t_L g793 ( .A(n_627), .B(n_664), .C(n_706), .Y(n_793) );
NAND2xp5_ASAP7_75t_SL g794 ( .A(n_636), .B(n_638), .Y(n_794) );
NOR3xp33_ASAP7_75t_L g795 ( .A(n_648), .B(n_704), .C(n_717), .Y(n_795) );
AOI211xp5_ASAP7_75t_L g796 ( .A1(n_618), .A2(n_667), .B(n_681), .C(n_651), .Y(n_796) );
OA211x2_ASAP7_75t_L g797 ( .A1(n_659), .A2(n_624), .B(n_716), .C(n_555), .Y(n_797) );
AND2x2_ASAP7_75t_L g798 ( .A(n_615), .B(n_617), .Y(n_798) );
NAND3xp33_ASAP7_75t_L g799 ( .A(n_654), .B(n_673), .C(n_618), .Y(n_799) );
AND2x2_ASAP7_75t_L g800 ( .A(n_615), .B(n_617), .Y(n_800) );
INVxp67_ASAP7_75t_SL g801 ( .A(n_716), .Y(n_801) );
NAND4xp75_ASAP7_75t_SL g802 ( .A(n_778), .B(n_776), .C(n_781), .D(n_721), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_726), .B(n_743), .Y(n_803) );
NOR4xp25_ASAP7_75t_L g804 ( .A(n_784), .B(n_759), .C(n_799), .D(n_760), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_798), .Y(n_805) );
INVx2_ASAP7_75t_L g806 ( .A(n_780), .Y(n_806) );
BUFx2_ASAP7_75t_L g807 ( .A(n_732), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_800), .Y(n_808) );
NOR3xp33_ASAP7_75t_SL g809 ( .A(n_724), .B(n_734), .C(n_731), .Y(n_809) );
NAND4xp75_ASAP7_75t_L g810 ( .A(n_797), .B(n_774), .C(n_733), .D(n_771), .Y(n_810) );
INVx1_ASAP7_75t_SL g811 ( .A(n_732), .Y(n_811) );
NAND4xp75_ASAP7_75t_L g812 ( .A(n_733), .B(n_721), .C(n_766), .D(n_768), .Y(n_812) );
INVx3_ASAP7_75t_L g813 ( .A(n_780), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_722), .Y(n_814) );
INVx5_ASAP7_75t_L g815 ( .A(n_757), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_796), .A2(n_767), .B1(n_772), .B2(n_781), .Y(n_816) );
BUFx2_ASAP7_75t_L g817 ( .A(n_801), .Y(n_817) );
OAI22x1_ASAP7_75t_L g818 ( .A1(n_751), .A2(n_738), .B1(n_755), .B2(n_783), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_726), .B(n_782), .Y(n_819) );
INVx2_ASAP7_75t_SL g820 ( .A(n_730), .Y(n_820) );
AND2x2_ASAP7_75t_L g821 ( .A(n_768), .B(n_723), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_761), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_723), .B(n_782), .Y(n_823) );
NAND4xp75_ASAP7_75t_L g824 ( .A(n_741), .B(n_747), .C(n_790), .D(n_748), .Y(n_824) );
XOR2xp5_ASAP7_75t_L g825 ( .A(n_783), .B(n_785), .Y(n_825) );
AND2x4_ASAP7_75t_L g826 ( .A(n_763), .B(n_723), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_779), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_762), .B(n_773), .Y(n_828) );
NAND4xp75_ASAP7_75t_SL g829 ( .A(n_791), .B(n_790), .C(n_788), .D(n_739), .Y(n_829) );
XOR2xp5_ASAP7_75t_L g830 ( .A(n_786), .B(n_764), .Y(n_830) );
OR2x2_ASAP7_75t_L g831 ( .A(n_746), .B(n_763), .Y(n_831) );
NOR3xp33_ASAP7_75t_SL g832 ( .A(n_769), .B(n_793), .C(n_794), .Y(n_832) );
INVx1_ASAP7_75t_SL g833 ( .A(n_730), .Y(n_833) );
XNOR2xp5_ASAP7_75t_L g834 ( .A(n_720), .B(n_758), .Y(n_834) );
INVx2_ASAP7_75t_SL g835 ( .A(n_757), .Y(n_835) );
NAND4xp25_ASAP7_75t_SL g836 ( .A(n_777), .B(n_765), .C(n_795), .D(n_756), .Y(n_836) );
NOR4xp25_ASAP7_75t_L g837 ( .A(n_777), .B(n_789), .C(n_725), .D(n_794), .Y(n_837) );
XOR2x2_ASAP7_75t_L g838 ( .A(n_750), .B(n_736), .Y(n_838) );
XNOR2xp5_ASAP7_75t_L g839 ( .A(n_773), .B(n_728), .Y(n_839) );
BUFx2_ASAP7_75t_L g840 ( .A(n_787), .Y(n_840) );
NAND4xp75_ASAP7_75t_SL g841 ( .A(n_791), .B(n_788), .C(n_739), .D(n_737), .Y(n_841) );
OR2x2_ASAP7_75t_L g842 ( .A(n_744), .B(n_770), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_729), .B(n_775), .Y(n_843) );
XNOR2xp5_ASAP7_75t_L g844 ( .A(n_753), .B(n_752), .Y(n_844) );
XOR2xp5_ASAP7_75t_L g845 ( .A(n_735), .B(n_742), .Y(n_845) );
AND2x4_ASAP7_75t_L g846 ( .A(n_729), .B(n_775), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_827), .Y(n_847) );
XNOR2xp5_ASAP7_75t_L g848 ( .A(n_825), .B(n_753), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_827), .Y(n_849) );
INVx2_ASAP7_75t_L g850 ( .A(n_806), .Y(n_850) );
OR2x2_ASAP7_75t_L g851 ( .A(n_819), .B(n_787), .Y(n_851) );
XOR2x2_ASAP7_75t_L g852 ( .A(n_816), .B(n_834), .Y(n_852) );
XOR2x2_ASAP7_75t_L g853 ( .A(n_829), .B(n_754), .Y(n_853) );
XOR2x2_ASAP7_75t_L g854 ( .A(n_802), .B(n_727), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_842), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_842), .Y(n_856) );
XOR2x2_ASAP7_75t_L g857 ( .A(n_810), .B(n_812), .Y(n_857) );
AND2x4_ASAP7_75t_L g858 ( .A(n_820), .B(n_787), .Y(n_858) );
INVxp67_ASAP7_75t_L g859 ( .A(n_836), .Y(n_859) );
XOR2x2_ASAP7_75t_L g860 ( .A(n_830), .B(n_807), .Y(n_860) );
CKINVDCx16_ASAP7_75t_R g861 ( .A(n_811), .Y(n_861) );
INVx2_ASAP7_75t_L g862 ( .A(n_806), .Y(n_862) );
INVxp67_ASAP7_75t_L g863 ( .A(n_840), .Y(n_863) );
OR2x2_ASAP7_75t_L g864 ( .A(n_843), .B(n_745), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_822), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_805), .Y(n_866) );
XOR2x2_ASAP7_75t_L g867 ( .A(n_841), .B(n_792), .Y(n_867) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_839), .B(n_749), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_808), .Y(n_869) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_817), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_814), .Y(n_871) );
XNOR2xp5_ASAP7_75t_L g872 ( .A(n_832), .B(n_740), .Y(n_872) );
OA22x2_ASAP7_75t_L g873 ( .A1(n_818), .A2(n_820), .B1(n_833), .B2(n_826), .Y(n_873) );
XOR2x2_ASAP7_75t_L g874 ( .A(n_838), .B(n_824), .Y(n_874) );
HB1xp67_ASAP7_75t_L g875 ( .A(n_870), .Y(n_875) );
XNOR2x1_ASAP7_75t_L g876 ( .A(n_857), .B(n_818), .Y(n_876) );
OA22x2_ASAP7_75t_L g877 ( .A1(n_859), .A2(n_826), .B1(n_846), .B2(n_804), .Y(n_877) );
AOI22xp5_ASAP7_75t_L g878 ( .A1(n_859), .A2(n_809), .B1(n_832), .B2(n_837), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_870), .Y(n_879) );
INVx1_ASAP7_75t_SL g880 ( .A(n_861), .Y(n_880) );
AOI22xp5_ASAP7_75t_L g881 ( .A1(n_857), .A2(n_852), .B1(n_854), .B2(n_874), .Y(n_881) );
AOI22x1_ASAP7_75t_L g882 ( .A1(n_872), .A2(n_809), .B1(n_813), .B2(n_826), .Y(n_882) );
OA22x2_ASAP7_75t_L g883 ( .A1(n_858), .A2(n_846), .B1(n_821), .B2(n_823), .Y(n_883) );
OA22x2_ASAP7_75t_L g884 ( .A1(n_858), .A2(n_846), .B1(n_821), .B2(n_823), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_871), .Y(n_885) );
OA22x2_ASAP7_75t_L g886 ( .A1(n_863), .A2(n_845), .B1(n_835), .B2(n_813), .Y(n_886) );
AOI22x1_ASAP7_75t_L g887 ( .A1(n_874), .A2(n_813), .B1(n_835), .B2(n_838), .Y(n_887) );
OA22x2_ASAP7_75t_L g888 ( .A1(n_863), .A2(n_844), .B1(n_803), .B2(n_828), .Y(n_888) );
OAI22xp5_ASAP7_75t_L g889 ( .A1(n_873), .A2(n_815), .B1(n_831), .B2(n_828), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_875), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_879), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_885), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_880), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_877), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_886), .Y(n_895) );
CKINVDCx16_ASAP7_75t_R g896 ( .A(n_881), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_878), .Y(n_897) );
AO22x2_ASAP7_75t_L g898 ( .A1(n_894), .A2(n_876), .B1(n_889), .B2(n_852), .Y(n_898) );
AOI22x1_ASAP7_75t_L g899 ( .A1(n_896), .A2(n_887), .B1(n_882), .B2(n_848), .Y(n_899) );
AOI22xp5_ASAP7_75t_L g900 ( .A1(n_893), .A2(n_854), .B1(n_888), .B2(n_867), .Y(n_900) );
OAI322xp33_ASAP7_75t_L g901 ( .A1(n_897), .A2(n_887), .A3(n_882), .B1(n_873), .B2(n_884), .C1(n_883), .C2(n_868), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_890), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g903 ( .A1(n_899), .A2(n_895), .B1(n_890), .B2(n_851), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_902), .Y(n_904) );
INVx2_ASAP7_75t_L g905 ( .A(n_898), .Y(n_905) );
AO22x2_ASAP7_75t_L g906 ( .A1(n_905), .A2(n_891), .B1(n_898), .B2(n_892), .Y(n_906) );
AOI22xp5_ASAP7_75t_L g907 ( .A1(n_903), .A2(n_900), .B1(n_860), .B2(n_891), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_906), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_907), .Y(n_909) );
OR2x2_ASAP7_75t_L g910 ( .A(n_908), .B(n_905), .Y(n_910) );
AND5x1_ASAP7_75t_L g911 ( .A(n_909), .B(n_901), .C(n_868), .D(n_904), .E(n_853), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_910), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_911), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_912), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_914), .Y(n_915) );
NAND4xp25_ASAP7_75t_L g916 ( .A(n_915), .B(n_913), .C(n_864), .D(n_865), .Y(n_916) );
INVxp67_ASAP7_75t_R g917 ( .A(n_916), .Y(n_917) );
AOI22xp5_ASAP7_75t_SL g918 ( .A1(n_917), .A2(n_856), .B1(n_855), .B2(n_869), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_918), .Y(n_919) );
AOI221xp5_ASAP7_75t_L g920 ( .A1(n_919), .A2(n_866), .B1(n_849), .B2(n_847), .C(n_850), .Y(n_920) );
AOI211xp5_ASAP7_75t_L g921 ( .A1(n_920), .A2(n_862), .B(n_850), .C(n_831), .Y(n_921) );
endmodule