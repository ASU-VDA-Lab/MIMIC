module fake_jpeg_23700_n_343 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_17),
.B(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_39),
.Y(n_48)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_8),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NAND3xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_11),
.C(n_15),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_6),
.Y(n_72)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_30),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_67),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_33),
.B1(n_16),
.B2(n_19),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_55),
.A2(n_57),
.B(n_60),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_33),
.B1(n_16),
.B2(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_35),
.A2(n_33),
.B1(n_19),
.B2(n_25),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_66),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_35),
.A2(n_33),
.B1(n_19),
.B2(n_25),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_30),
.Y(n_64)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_16),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_37),
.A2(n_25),
.B1(n_19),
.B2(n_26),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_42),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_25),
.B1(n_20),
.B2(n_24),
.Y(n_69)
);

BUFx24_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_73),
.Y(n_99)
);

OAI22x1_ASAP7_75t_L g106 ( 
.A1(n_72),
.A2(n_61),
.B1(n_59),
.B2(n_48),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_64),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_78),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_22),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_75),
.B(n_88),
.Y(n_118)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_85),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_91),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_27),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_51),
.Y(n_89)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_54),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_67),
.A2(n_38),
.B(n_43),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_92),
.A2(n_57),
.B1(n_55),
.B2(n_65),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_43),
.C(n_38),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_95),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_43),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_97),
.Y(n_119)
);

BUFx4f_ASAP7_75t_SL g97 ( 
.A(n_65),
.Y(n_97)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_102),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_79),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_104),
.A2(n_82),
.B(n_93),
.Y(n_150)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_111),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_70),
.B(n_91),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_47),
.B1(n_68),
.B2(n_25),
.Y(n_107)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_113),
.Y(n_138)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_84),
.A2(n_65),
.B1(n_20),
.B2(n_24),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_84),
.A2(n_38),
.B1(n_43),
.B2(n_60),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_117),
.A2(n_84),
.B1(n_47),
.B2(n_87),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_78),
.B(n_58),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_121),
.B(n_124),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_70),
.B(n_53),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_73),
.Y(n_133)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_125),
.Y(n_160)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_128),
.Y(n_157)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_93),
.B1(n_92),
.B2(n_100),
.Y(n_152)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_137),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_132),
.A2(n_72),
.B(n_81),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_139),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_134),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_110),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_120),
.B(n_75),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_142),
.B(n_144),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_120),
.B(n_106),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_146),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_118),
.B(n_86),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_110),
.B(n_86),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_148),
.Y(n_168)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_103),
.B(n_95),
.Y(n_149)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_150),
.A2(n_104),
.B(n_107),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_151),
.B(n_166),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_152),
.A2(n_53),
.B1(n_47),
.B2(n_50),
.Y(n_195)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_169),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_175),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_149),
.A2(n_103),
.B(n_95),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_159),
.A2(n_165),
.B(n_170),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_126),
.A2(n_77),
.B1(n_117),
.B2(n_94),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_163),
.B1(n_164),
.B2(n_154),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_141),
.A2(n_117),
.B1(n_72),
.B2(n_124),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_126),
.A2(n_117),
.B1(n_83),
.B2(n_71),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_150),
.A2(n_141),
.B(n_133),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_174),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_140),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_43),
.Y(n_175)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_179),
.Y(n_207)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_176),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_180),
.A2(n_185),
.B(n_186),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_174),
.A2(n_127),
.B1(n_148),
.B2(n_144),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_181),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_173),
.B(n_146),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_183),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_165),
.A2(n_171),
.B(n_159),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_184),
.A2(n_194),
.B(n_41),
.Y(n_222)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_128),
.Y(n_188)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_189),
.A2(n_199),
.B1(n_152),
.B2(n_155),
.Y(n_208)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_153),
.A2(n_123),
.B1(n_113),
.B2(n_143),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_195),
.A2(n_116),
.B1(n_163),
.B2(n_167),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_145),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_197),
.C(n_20),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_108),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_142),
.B1(n_96),
.B2(n_143),
.Y(n_199)
);

INVxp33_ASAP7_75t_SL g201 ( 
.A(n_160),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_201),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_137),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_202),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_102),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_203),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_208),
.A2(n_42),
.B1(n_37),
.B2(n_32),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_177),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_210),
.B(n_215),
.C(n_216),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_211),
.A2(n_213),
.B1(n_219),
.B2(n_182),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_185),
.A2(n_155),
.B1(n_162),
.B2(n_168),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_170),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_177),
.B(n_168),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_186),
.A2(n_162),
.B1(n_160),
.B2(n_167),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_217),
.A2(n_220),
.B1(n_224),
.B2(n_225),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_50),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_228),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_184),
.A2(n_116),
.B1(n_111),
.B2(n_112),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_203),
.A2(n_53),
.B1(n_50),
.B2(n_125),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_222),
.A2(n_217),
.B(n_209),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_180),
.A2(n_134),
.B1(n_135),
.B2(n_90),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_80),
.B1(n_21),
.B2(n_22),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_192),
.A2(n_188),
.B1(n_198),
.B2(n_187),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_226),
.A2(n_18),
.B1(n_21),
.B2(n_22),
.Y(n_250)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_230),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_224),
.Y(n_231)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_231),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_232),
.A2(n_243),
.B1(n_247),
.B2(n_248),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_190),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_233),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_236),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_193),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_237),
.B(n_245),
.Y(n_272)
);

AND2x6_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_196),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_219),
.A2(n_179),
.B1(n_200),
.B2(n_178),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_26),
.B(n_24),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_205),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_241),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_221),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_242),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_208),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_204),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_246),
.A2(n_250),
.B1(n_29),
.B2(n_23),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_206),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_18),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_227),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_251),
.A2(n_223),
.B1(n_225),
.B2(n_228),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_0),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_212),
.C(n_240),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_250),
.Y(n_280)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

NOR2xp67_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_216),
.Y(n_259)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_259),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_218),
.C(n_215),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_270),
.C(n_271),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_236),
.A2(n_211),
.B1(n_26),
.B2(n_18),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_262),
.A2(n_265),
.B1(n_267),
.B2(n_12),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_239),
.A2(n_17),
.B1(n_21),
.B2(n_29),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_244),
.A2(n_23),
.B1(n_17),
.B2(n_29),
.Y(n_267)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_234),
.A2(n_23),
.B1(n_37),
.B2(n_42),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_269),
.A2(n_230),
.B1(n_232),
.B2(n_234),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_235),
.C(n_242),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_238),
.B(n_27),
.C(n_28),
.Y(n_271)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_273),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_257),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_279),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_272),
.Y(n_275)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_275),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_247),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_253),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_257),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_283),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_28),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_282),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_28),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_13),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_256),
.C(n_271),
.Y(n_291)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_255),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_287),
.A2(n_266),
.B(n_254),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_14),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_SL g289 ( 
.A1(n_260),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_1),
.B1(n_2),
.B2(n_32),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_291),
.A2(n_294),
.B(n_295),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_264),
.Y(n_292)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_292),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_297),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_270),
.Y(n_297)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_298),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_284),
.A2(n_277),
.B(n_276),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_300),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_269),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_304),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_303),
.A2(n_289),
.B1(n_278),
.B2(n_32),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_32),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_306),
.A2(n_312),
.B(n_12),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_273),
.Y(n_307)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_307),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_286),
.C(n_291),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_308),
.A2(n_314),
.B(n_316),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_31),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_289),
.B(n_32),
.Y(n_312)
);

MAJx2_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_289),
.C(n_14),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_31),
.C(n_27),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_300),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_308),
.C(n_317),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_309),
.B(n_303),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_319),
.A2(n_323),
.B(n_325),
.Y(n_330)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_320),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_322),
.A2(n_3),
.B1(n_4),
.B2(n_14),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_310),
.B(n_9),
.Y(n_323)
);

OAI21xp33_ASAP7_75t_L g324 ( 
.A1(n_315),
.A2(n_12),
.B(n_15),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_324),
.B(n_5),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_28),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_327),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_313),
.C(n_316),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_328),
.A2(n_331),
.B(n_3),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_314),
.C(n_5),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_3),
.Y(n_334)
);

INVxp33_ASAP7_75t_L g336 ( 
.A(n_334),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_333),
.B(n_329),
.Y(n_337)
);

OAI21x1_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_335),
.B(n_330),
.Y(n_338)
);

MAJx2_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_326),
.C(n_4),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_4),
.B1(n_2),
.B2(n_1),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_340),
.A2(n_1),
.B(n_2),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_36),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_342),
.B(n_36),
.Y(n_343)
);


endmodule