module real_aes_6897_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_335;
wire n_177;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g111 ( .A(n_0), .Y(n_111) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_1), .A2(n_153), .B(n_156), .C(n_236), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_2), .A2(n_182), .B(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g482 ( .A(n_3), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_4), .B(n_212), .Y(n_211) );
AOI21xp33_ASAP7_75t_L g465 ( .A1(n_5), .A2(n_182), .B(n_466), .Y(n_465) );
AND2x6_ASAP7_75t_L g153 ( .A(n_6), .B(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g249 ( .A(n_7), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_8), .B(n_42), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_9), .A2(n_181), .B(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_10), .B(n_165), .Y(n_238) );
INVx1_ASAP7_75t_L g470 ( .A(n_11), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_12), .B(n_206), .Y(n_505) );
INVx1_ASAP7_75t_L g145 ( .A(n_13), .Y(n_145) );
INVx1_ASAP7_75t_L g517 ( .A(n_14), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_15), .A2(n_78), .B1(n_125), .B2(n_126), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_15), .Y(n_125) );
A2O1A1Ixp33_ASAP7_75t_L g270 ( .A1(n_16), .A2(n_190), .B(n_271), .C(n_273), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_17), .B(n_212), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_18), .B(n_448), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_19), .B(n_182), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_20), .B(n_196), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_21), .A2(n_206), .B(n_257), .C(n_259), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_22), .B(n_212), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_23), .B(n_165), .Y(n_164) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_24), .A2(n_192), .B(n_273), .C(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_25), .B(n_165), .Y(n_220) );
CKINVDCx16_ASAP7_75t_R g147 ( .A(n_26), .Y(n_147) );
INVx1_ASAP7_75t_L g219 ( .A(n_27), .Y(n_219) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_28), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_29), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_30), .B(n_165), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_31), .A2(n_102), .B1(n_113), .B2(n_737), .Y(n_101) );
INVx1_ASAP7_75t_L g188 ( .A(n_32), .Y(n_188) );
INVx1_ASAP7_75t_L g460 ( .A(n_33), .Y(n_460) );
INVx2_ASAP7_75t_L g151 ( .A(n_34), .Y(n_151) );
AOI222xp33_ASAP7_75t_SL g123 ( .A1(n_35), .A2(n_124), .B1(n_127), .B2(n_721), .C1(n_722), .C2(n_724), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_36), .Y(n_240) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_37), .A2(n_206), .B(n_207), .C(n_209), .Y(n_205) );
INVxp67_ASAP7_75t_L g191 ( .A(n_38), .Y(n_191) );
CKINVDCx14_ASAP7_75t_R g204 ( .A(n_39), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_40), .A2(n_156), .B(n_218), .C(n_222), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_41), .A2(n_153), .B(n_156), .C(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g459 ( .A(n_43), .Y(n_459) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_44), .A2(n_167), .B(n_247), .C(n_248), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_45), .B(n_165), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_46), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_47), .Y(n_184) );
INVx1_ASAP7_75t_L g255 ( .A(n_48), .Y(n_255) );
CKINVDCx16_ASAP7_75t_R g461 ( .A(n_49), .Y(n_461) );
OAI22xp5_ASAP7_75t_SL g732 ( .A1(n_50), .A2(n_60), .B1(n_733), .B2(n_734), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_50), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_51), .B(n_182), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_52), .A2(n_156), .B1(n_259), .B2(n_458), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_53), .Y(n_497) );
CKINVDCx16_ASAP7_75t_R g479 ( .A(n_54), .Y(n_479) );
CKINVDCx14_ASAP7_75t_R g245 ( .A(n_55), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_56), .A2(n_209), .B(n_247), .C(n_469), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_57), .Y(n_122) );
INVx1_ASAP7_75t_L g467 ( .A(n_58), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_59), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_60), .Y(n_734) );
INVx1_ASAP7_75t_L g154 ( .A(n_61), .Y(n_154) );
INVx1_ASAP7_75t_L g144 ( .A(n_62), .Y(n_144) );
INVx1_ASAP7_75t_SL g208 ( .A(n_63), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_64), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_65), .B(n_212), .Y(n_261) );
INVx1_ASAP7_75t_L g160 ( .A(n_66), .Y(n_160) );
A2O1A1Ixp33_ASAP7_75t_SL g447 ( .A1(n_67), .A2(n_209), .B(n_448), .C(n_449), .Y(n_447) );
INVxp67_ASAP7_75t_L g450 ( .A(n_68), .Y(n_450) );
INVx1_ASAP7_75t_L g106 ( .A(n_69), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_70), .A2(n_182), .B(n_244), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_71), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_72), .A2(n_182), .B(n_268), .Y(n_267) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_73), .Y(n_463) );
INVx1_ASAP7_75t_L g523 ( .A(n_74), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_75), .A2(n_181), .B(n_183), .Y(n_180) );
CKINVDCx16_ASAP7_75t_R g216 ( .A(n_76), .Y(n_216) );
INVx1_ASAP7_75t_L g269 ( .A(n_77), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_78), .Y(n_126) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_79), .A2(n_153), .B(n_156), .C(n_525), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_80), .A2(n_182), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g272 ( .A(n_81), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_82), .B(n_189), .Y(n_494) );
INVx2_ASAP7_75t_L g142 ( .A(n_83), .Y(n_142) );
INVx1_ASAP7_75t_L g237 ( .A(n_84), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_85), .B(n_448), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_86), .A2(n_153), .B(n_156), .C(n_481), .Y(n_480) );
OR2x2_ASAP7_75t_L g108 ( .A(n_87), .B(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g435 ( .A(n_87), .B(n_110), .Y(n_435) );
INVx2_ASAP7_75t_L g720 ( .A(n_87), .Y(n_720) );
A2O1A1Ixp33_ASAP7_75t_L g155 ( .A1(n_88), .A2(n_156), .B(n_159), .C(n_169), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_89), .B(n_174), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_90), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_91), .A2(n_153), .B(n_156), .C(n_503), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_92), .Y(n_509) );
INVx1_ASAP7_75t_L g446 ( .A(n_93), .Y(n_446) );
CKINVDCx16_ASAP7_75t_R g514 ( .A(n_94), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_95), .B(n_189), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_96), .B(n_140), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_97), .B(n_140), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_98), .B(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g258 ( .A(n_99), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_100), .A2(n_182), .B(n_445), .Y(n_444) );
CKINVDCx6p67_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g738 ( .A(n_103), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g121 ( .A(n_108), .Y(n_121) );
INVx1_ASAP7_75t_SL g736 ( .A(n_108), .Y(n_736) );
NOR2x2_ASAP7_75t_L g726 ( .A(n_109), .B(n_720), .Y(n_726) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g719 ( .A(n_110), .B(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AOI22xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_123), .B1(n_727), .B2(n_729), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_116), .B(n_119), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g728 ( .A(n_117), .Y(n_728) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_119), .A2(n_730), .B(n_735), .Y(n_729) );
NOR2xp33_ASAP7_75t_SL g119 ( .A(n_120), .B(n_122), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g721 ( .A(n_124), .Y(n_721) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_435), .B1(n_436), .B2(n_717), .Y(n_127) );
OAI22xp5_ASAP7_75t_SL g730 ( .A1(n_128), .A2(n_129), .B1(n_731), .B2(n_732), .Y(n_730) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_SL g722 ( .A1(n_129), .A2(n_435), .B1(n_717), .B2(n_723), .Y(n_722) );
OR2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_369), .Y(n_129) );
NAND5xp2_ASAP7_75t_L g130 ( .A(n_131), .B(n_298), .C(n_328), .D(n_349), .E(n_355), .Y(n_130) );
AOI221xp5_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_228), .B1(n_262), .B2(n_264), .C(n_275), .Y(n_131) );
INVxp67_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_225), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_197), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
A2O1A1Ixp33_ASAP7_75t_SL g349 ( .A1(n_136), .A2(n_213), .B(n_350), .C(n_353), .Y(n_349) );
AND2x2_ASAP7_75t_L g419 ( .A(n_136), .B(n_214), .Y(n_419) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_175), .Y(n_136) );
AND2x2_ASAP7_75t_L g277 ( .A(n_137), .B(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g281 ( .A(n_137), .B(n_278), .Y(n_281) );
OR2x2_ASAP7_75t_L g307 ( .A(n_137), .B(n_214), .Y(n_307) );
AND2x2_ASAP7_75t_L g309 ( .A(n_137), .B(n_200), .Y(n_309) );
AND2x2_ASAP7_75t_L g327 ( .A(n_137), .B(n_199), .Y(n_327) );
INVx1_ASAP7_75t_L g360 ( .A(n_137), .Y(n_360) );
INVx2_ASAP7_75t_SL g137 ( .A(n_138), .Y(n_137) );
BUFx2_ASAP7_75t_L g227 ( .A(n_138), .Y(n_227) );
AND2x2_ASAP7_75t_L g263 ( .A(n_138), .B(n_200), .Y(n_263) );
AND2x2_ASAP7_75t_L g416 ( .A(n_138), .B(n_214), .Y(n_416) );
AO21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_146), .B(n_171), .Y(n_138) );
INVx3_ASAP7_75t_L g212 ( .A(n_139), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_139), .B(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_139), .B(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_SL g496 ( .A(n_139), .B(n_497), .Y(n_496) );
INVx4_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_140), .Y(n_201) );
OA21x2_ASAP7_75t_L g443 ( .A1(n_140), .A2(n_444), .B(n_451), .Y(n_443) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g178 ( .A(n_141), .Y(n_178) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AND2x2_ASAP7_75t_SL g174 ( .A(n_142), .B(n_143), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
OAI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_155), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_L g215 ( .A1(n_148), .A2(n_174), .B(n_216), .C(n_217), .Y(n_215) );
OAI21xp5_ASAP7_75t_L g233 ( .A1(n_148), .A2(n_234), .B(n_235), .Y(n_233) );
OAI22xp33_ASAP7_75t_L g456 ( .A1(n_148), .A2(n_170), .B1(n_457), .B2(n_461), .Y(n_456) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_148), .A2(n_479), .B(n_480), .Y(n_478) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_148), .A2(n_523), .B(n_524), .Y(n_522) );
NAND2x1p5_ASAP7_75t_L g148 ( .A(n_149), .B(n_153), .Y(n_148) );
AND2x4_ASAP7_75t_L g182 ( .A(n_149), .B(n_153), .Y(n_182) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_152), .Y(n_149) );
INVx1_ASAP7_75t_L g193 ( .A(n_150), .Y(n_193) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g157 ( .A(n_151), .Y(n_157) );
INVx1_ASAP7_75t_L g260 ( .A(n_151), .Y(n_260) );
INVx1_ASAP7_75t_L g158 ( .A(n_152), .Y(n_158) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_152), .Y(n_163) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_152), .Y(n_165) );
INVx3_ASAP7_75t_L g190 ( .A(n_152), .Y(n_190) );
INVx1_ASAP7_75t_L g448 ( .A(n_152), .Y(n_448) );
INVx4_ASAP7_75t_SL g170 ( .A(n_153), .Y(n_170) );
BUFx3_ASAP7_75t_L g222 ( .A(n_153), .Y(n_222) );
INVx5_ASAP7_75t_L g185 ( .A(n_156), .Y(n_185) );
AND2x6_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
BUFx3_ASAP7_75t_L g168 ( .A(n_157), .Y(n_168) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_157), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_164), .C(n_166), .Y(n_159) );
O2A1O1Ixp5_ASAP7_75t_L g236 ( .A1(n_161), .A2(n_166), .B(n_237), .C(n_238), .Y(n_236) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
OAI22xp5_ASAP7_75t_SL g458 ( .A1(n_162), .A2(n_163), .B1(n_459), .B2(n_460), .Y(n_458) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx4_ASAP7_75t_L g192 ( .A(n_163), .Y(n_192) );
INVx4_ASAP7_75t_L g206 ( .A(n_165), .Y(n_206) );
INVx2_ASAP7_75t_L g247 ( .A(n_165), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_166), .A2(n_494), .B(n_495), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_166), .A2(n_526), .B(n_527), .Y(n_525) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g273 ( .A(n_168), .Y(n_273) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_SL g183 ( .A1(n_170), .A2(n_184), .B(n_185), .C(n_186), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g203 ( .A1(n_170), .A2(n_185), .B(n_204), .C(n_205), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_SL g244 ( .A1(n_170), .A2(n_185), .B(n_245), .C(n_246), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_SL g254 ( .A1(n_170), .A2(n_185), .B(n_255), .C(n_256), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_SL g268 ( .A1(n_170), .A2(n_185), .B(n_269), .C(n_270), .Y(n_268) );
O2A1O1Ixp33_ASAP7_75t_L g445 ( .A1(n_170), .A2(n_185), .B(n_446), .C(n_447), .Y(n_445) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_170), .A2(n_185), .B(n_467), .C(n_468), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g513 ( .A1(n_170), .A2(n_185), .B(n_514), .C(n_515), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
INVx1_ASAP7_75t_L g196 ( .A(n_173), .Y(n_196) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_173), .A2(n_501), .B(n_508), .Y(n_500) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g232 ( .A(n_174), .Y(n_232) );
OA21x2_ASAP7_75t_L g242 ( .A1(n_174), .A2(n_243), .B(n_250), .Y(n_242) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_174), .A2(n_512), .B(n_518), .Y(n_511) );
AND2x2_ASAP7_75t_L g297 ( .A(n_175), .B(n_198), .Y(n_297) );
OR2x2_ASAP7_75t_L g301 ( .A(n_175), .B(n_214), .Y(n_301) );
AND2x2_ASAP7_75t_L g326 ( .A(n_175), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g373 ( .A(n_175), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_175), .B(n_335), .Y(n_421) );
AO21x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_179), .B(n_194), .Y(n_175) );
INVx1_ASAP7_75t_L g279 ( .A(n_176), .Y(n_279) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_176), .A2(n_522), .B(n_528), .Y(n_521) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AOI21xp5_ASAP7_75t_SL g490 ( .A1(n_177), .A2(n_491), .B(n_492), .Y(n_490) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AO21x2_ASAP7_75t_L g455 ( .A1(n_178), .A2(n_456), .B(n_462), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_178), .B(n_463), .Y(n_462) );
AO21x2_ASAP7_75t_L g477 ( .A1(n_178), .A2(n_478), .B(n_485), .Y(n_477) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
OA21x2_ASAP7_75t_L g278 ( .A1(n_180), .A2(n_195), .B(n_279), .Y(n_278) );
BUFx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_187), .B(n_193), .Y(n_186) );
OAI22xp33_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B1(n_191), .B2(n_192), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g218 ( .A1(n_189), .A2(n_219), .B(n_220), .C(n_221), .Y(n_218) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_189), .A2(n_482), .B(n_483), .C(n_484), .Y(n_481) );
INVx5_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_190), .B(n_249), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_190), .B(n_450), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_190), .B(n_470), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_192), .B(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_192), .B(n_272), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_192), .B(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g221 ( .A(n_193), .Y(n_221) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
OAI322xp33_ASAP7_75t_L g422 ( .A1(n_197), .A2(n_358), .A3(n_381), .B1(n_402), .B2(n_423), .C1(n_425), .C2(n_426), .Y(n_422) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_198), .B(n_278), .Y(n_425) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_213), .Y(n_198) );
AND2x2_ASAP7_75t_L g226 ( .A(n_199), .B(n_227), .Y(n_226) );
AND2x4_ASAP7_75t_L g294 ( .A(n_199), .B(n_214), .Y(n_294) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g335 ( .A(n_200), .B(n_214), .Y(n_335) );
AND2x2_ASAP7_75t_L g379 ( .A(n_200), .B(n_213), .Y(n_379) );
OA21x2_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_211), .Y(n_200) );
OA21x2_ASAP7_75t_L g252 ( .A1(n_201), .A2(n_253), .B(n_261), .Y(n_252) );
OA21x2_ASAP7_75t_L g266 ( .A1(n_201), .A2(n_267), .B(n_274), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_206), .B(n_208), .Y(n_207) );
INVx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_210), .Y(n_506) );
OA21x2_ASAP7_75t_L g464 ( .A1(n_212), .A2(n_465), .B(n_471), .Y(n_464) );
AND2x2_ASAP7_75t_L g262 ( .A(n_213), .B(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g280 ( .A(n_213), .B(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_213), .B(n_309), .Y(n_433) );
INVx3_ASAP7_75t_SL g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g225 ( .A(n_214), .B(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_214), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g347 ( .A(n_214), .B(n_278), .Y(n_347) );
AND2x2_ASAP7_75t_L g374 ( .A(n_214), .B(n_309), .Y(n_374) );
OR2x2_ASAP7_75t_L g430 ( .A(n_214), .B(n_281), .Y(n_430) );
OR2x6_ASAP7_75t_L g214 ( .A(n_215), .B(n_223), .Y(n_214) );
INVx1_ASAP7_75t_SL g316 ( .A(n_225), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_226), .B(n_347), .Y(n_348) );
AND2x2_ASAP7_75t_L g382 ( .A(n_226), .B(n_372), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_226), .B(n_305), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_226), .B(n_427), .Y(n_426) );
OAI31xp33_ASAP7_75t_L g400 ( .A1(n_228), .A2(n_262), .A3(n_401), .B(n_403), .Y(n_400) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_241), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g367 ( .A(n_229), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g383 ( .A(n_229), .B(n_318), .Y(n_383) );
OR2x2_ASAP7_75t_L g390 ( .A(n_229), .B(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g402 ( .A(n_229), .B(n_291), .Y(n_402) );
CKINVDCx16_ASAP7_75t_R g229 ( .A(n_230), .Y(n_229) );
OR2x2_ASAP7_75t_L g336 ( .A(n_230), .B(n_337), .Y(n_336) );
BUFx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g264 ( .A(n_231), .B(n_265), .Y(n_264) );
INVx4_ASAP7_75t_L g285 ( .A(n_231), .Y(n_285) );
AND2x2_ASAP7_75t_L g322 ( .A(n_231), .B(n_266), .Y(n_322) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_239), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_232), .B(n_486), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_232), .B(n_509), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_232), .B(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g321 ( .A(n_241), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_SL g391 ( .A(n_241), .Y(n_391) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_251), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_242), .B(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g291 ( .A(n_242), .B(n_252), .Y(n_291) );
INVx2_ASAP7_75t_L g311 ( .A(n_242), .Y(n_311) );
AND2x2_ASAP7_75t_L g325 ( .A(n_242), .B(n_252), .Y(n_325) );
AND2x2_ASAP7_75t_L g332 ( .A(n_242), .B(n_288), .Y(n_332) );
BUFx3_ASAP7_75t_L g342 ( .A(n_242), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_242), .B(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g287 ( .A(n_251), .Y(n_287) );
AND2x2_ASAP7_75t_L g295 ( .A(n_251), .B(n_285), .Y(n_295) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g265 ( .A(n_252), .B(n_266), .Y(n_265) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_252), .Y(n_319) );
INVx2_ASAP7_75t_L g484 ( .A(n_259), .Y(n_484) );
INVx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx2_ASAP7_75t_SL g302 ( .A(n_263), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_263), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_263), .B(n_372), .Y(n_393) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_264), .B(n_342), .Y(n_395) );
INVx1_ASAP7_75t_SL g429 ( .A(n_264), .Y(n_429) );
INVx1_ASAP7_75t_SL g337 ( .A(n_265), .Y(n_337) );
INVx1_ASAP7_75t_SL g288 ( .A(n_266), .Y(n_288) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_266), .Y(n_299) );
OR2x2_ASAP7_75t_L g310 ( .A(n_266), .B(n_285), .Y(n_310) );
AND2x2_ASAP7_75t_L g324 ( .A(n_266), .B(n_285), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_266), .B(n_314), .Y(n_376) );
A2O1A1Ixp33_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_280), .B(n_282), .C(n_293), .Y(n_275) );
AOI31xp33_ASAP7_75t_L g392 ( .A1(n_276), .A2(n_393), .A3(n_394), .B(n_395), .Y(n_392) );
AND2x2_ASAP7_75t_L g365 ( .A(n_277), .B(n_294), .Y(n_365) );
BUFx3_ASAP7_75t_L g305 ( .A(n_278), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_278), .B(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g341 ( .A(n_278), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_278), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g296 ( .A(n_281), .Y(n_296) );
OAI222xp33_ASAP7_75t_L g405 ( .A1(n_281), .A2(n_406), .B1(n_409), .B2(n_410), .C1(n_411), .C2(n_412), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_283), .B(n_289), .Y(n_282) );
INVx1_ASAP7_75t_L g411 ( .A(n_283), .Y(n_411) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_285), .B(n_288), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_285), .B(n_311), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_285), .B(n_286), .Y(n_381) );
INVx1_ASAP7_75t_L g432 ( .A(n_285), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g362 ( .A(n_286), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g434 ( .A(n_286), .Y(n_434) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx2_ASAP7_75t_L g314 ( .A(n_287), .Y(n_314) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_288), .Y(n_357) );
AOI32xp33_ASAP7_75t_L g293 ( .A1(n_289), .A2(n_294), .A3(n_295), .B1(n_296), .B2(n_297), .Y(n_293) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_291), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g368 ( .A(n_291), .Y(n_368) );
OR2x2_ASAP7_75t_L g409 ( .A(n_291), .B(n_310), .Y(n_409) );
INVx1_ASAP7_75t_L g345 ( .A(n_292), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_294), .B(n_305), .Y(n_330) );
INVx3_ASAP7_75t_L g339 ( .A(n_294), .Y(n_339) );
AOI322xp5_ASAP7_75t_L g355 ( .A1(n_294), .A2(n_339), .A3(n_356), .B1(n_358), .B2(n_361), .C1(n_365), .C2(n_366), .Y(n_355) );
AND2x2_ASAP7_75t_L g331 ( .A(n_295), .B(n_332), .Y(n_331) );
INVxp67_ASAP7_75t_L g408 ( .A(n_295), .Y(n_408) );
A2O1A1O1Ixp25_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B(n_303), .C(n_311), .D(n_312), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_299), .B(n_342), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
OAI221xp5_ASAP7_75t_L g312 ( .A1(n_301), .A2(n_313), .B1(n_316), .B2(n_317), .C(n_320), .Y(n_312) );
INVx1_ASAP7_75t_SL g427 ( .A(n_301), .Y(n_427) );
AOI21xp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_308), .B(n_310), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_305), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OAI221xp5_ASAP7_75t_SL g397 ( .A1(n_307), .A2(n_391), .B1(n_398), .B2(n_399), .C(n_400), .Y(n_397) );
OAI222xp33_ASAP7_75t_L g428 ( .A1(n_308), .A2(n_429), .B1(n_430), .B2(n_431), .C1(n_433), .C2(n_434), .Y(n_428) );
AND2x2_ASAP7_75t_L g386 ( .A(n_309), .B(n_372), .Y(n_386) );
AOI21xp5_ASAP7_75t_L g398 ( .A1(n_309), .A2(n_324), .B(n_371), .Y(n_398) );
INVx1_ASAP7_75t_L g412 ( .A(n_309), .Y(n_412) );
INVx2_ASAP7_75t_SL g315 ( .A(n_310), .Y(n_315) );
AND2x2_ASAP7_75t_L g318 ( .A(n_311), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_SL g352 ( .A(n_314), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_314), .B(n_324), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_315), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_315), .B(n_325), .Y(n_354) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OAI21xp5_ASAP7_75t_SL g320 ( .A1(n_321), .A2(n_323), .B(n_326), .Y(n_320) );
INVx1_ASAP7_75t_SL g338 ( .A(n_322), .Y(n_338) );
AND2x2_ASAP7_75t_L g385 ( .A(n_322), .B(n_368), .Y(n_385) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
AND2x2_ASAP7_75t_L g424 ( .A(n_324), .B(n_342), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_325), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_SL g410 ( .A(n_326), .Y(n_410) );
AOI221xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_331), .B1(n_333), .B2(n_340), .C(n_343), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_336), .B1(n_338), .B2(n_339), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OAI22xp33_ASAP7_75t_L g343 ( .A1(n_337), .A2(n_344), .B1(n_346), .B2(n_348), .Y(n_343) );
OR2x2_ASAP7_75t_L g414 ( .A(n_338), .B(n_342), .Y(n_414) );
OR2x2_ASAP7_75t_L g417 ( .A(n_338), .B(n_352), .Y(n_417) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OAI221xp5_ASAP7_75t_L g413 ( .A1(n_359), .A2(n_414), .B1(n_415), .B2(n_417), .C(n_418), .Y(n_413) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVxp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND3xp33_ASAP7_75t_SL g369 ( .A(n_370), .B(n_384), .C(n_396), .Y(n_369) );
AOI222xp33_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_375), .B1(n_377), .B2(n_380), .C1(n_382), .C2(n_383), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_372), .B(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g394 ( .A(n_374), .Y(n_394) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVxp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AOI221xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B1(n_387), .B2(n_389), .C(n_392), .Y(n_384) );
INVx1_ASAP7_75t_L g399 ( .A(n_385), .Y(n_399) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI21xp33_ASAP7_75t_L g418 ( .A1(n_389), .A2(n_419), .B(n_420), .Y(n_418) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
NOR5xp2_ASAP7_75t_L g396 ( .A(n_397), .B(n_405), .C(n_413), .D(n_422), .E(n_428), .Y(n_396) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
INVxp67_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g723 ( .A(n_436), .Y(n_723) );
AND2x2_ASAP7_75t_SL g436 ( .A(n_437), .B(n_654), .Y(n_436) );
NOR4xp25_ASAP7_75t_L g437 ( .A(n_438), .B(n_584), .C(n_615), .D(n_634), .Y(n_437) );
NAND4xp25_ASAP7_75t_L g438 ( .A(n_439), .B(n_542), .C(n_557), .D(n_575), .Y(n_438) );
AOI222xp33_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_487), .B1(n_519), .B2(n_530), .C1(n_535), .C2(n_537), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_472), .Y(n_440) );
INVx1_ASAP7_75t_L g598 ( .A(n_441), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_452), .Y(n_441) );
AND2x2_ASAP7_75t_L g473 ( .A(n_442), .B(n_464), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_442), .B(n_476), .Y(n_627) );
INVx3_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g534 ( .A(n_443), .B(n_454), .Y(n_534) );
AND2x2_ASAP7_75t_L g543 ( .A(n_443), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g569 ( .A(n_443), .Y(n_569) );
AND2x2_ASAP7_75t_L g590 ( .A(n_443), .B(n_454), .Y(n_590) );
BUFx2_ASAP7_75t_L g613 ( .A(n_443), .Y(n_613) );
AND2x2_ASAP7_75t_L g637 ( .A(n_443), .B(n_455), .Y(n_637) );
AND2x2_ASAP7_75t_L g701 ( .A(n_443), .B(n_464), .Y(n_701) );
AND2x2_ASAP7_75t_L g602 ( .A(n_452), .B(n_533), .Y(n_602) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_453), .B(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_464), .Y(n_453) );
OR2x2_ASAP7_75t_L g562 ( .A(n_454), .B(n_477), .Y(n_562) );
AND2x2_ASAP7_75t_L g574 ( .A(n_454), .B(n_533), .Y(n_574) );
BUFx2_ASAP7_75t_L g706 ( .A(n_454), .Y(n_706) );
INVx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g475 ( .A(n_455), .B(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g556 ( .A(n_455), .B(n_477), .Y(n_556) );
AND2x2_ASAP7_75t_L g609 ( .A(n_455), .B(n_464), .Y(n_609) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_455), .Y(n_645) );
AND2x2_ASAP7_75t_L g532 ( .A(n_464), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_SL g544 ( .A(n_464), .Y(n_544) );
INVx2_ASAP7_75t_L g555 ( .A(n_464), .Y(n_555) );
BUFx2_ASAP7_75t_L g579 ( .A(n_464), .Y(n_579) );
AND2x2_ASAP7_75t_SL g636 ( .A(n_464), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
AOI332xp33_ASAP7_75t_L g557 ( .A1(n_473), .A2(n_558), .A3(n_562), .B1(n_563), .B2(n_567), .B3(n_570), .C1(n_571), .C2(n_573), .Y(n_557) );
NAND2x1_ASAP7_75t_L g642 ( .A(n_473), .B(n_533), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_473), .B(n_547), .Y(n_693) );
A2O1A1Ixp33_ASAP7_75t_SL g575 ( .A1(n_474), .A2(n_576), .B(n_579), .C(n_580), .Y(n_575) );
AND2x2_ASAP7_75t_L g714 ( .A(n_474), .B(n_555), .Y(n_714) );
INVx3_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
OR2x2_ASAP7_75t_L g611 ( .A(n_475), .B(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g616 ( .A(n_475), .B(n_613), .Y(n_616) );
INVx1_ASAP7_75t_L g547 ( .A(n_476), .Y(n_547) );
AND2x2_ASAP7_75t_L g650 ( .A(n_476), .B(n_609), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_476), .B(n_590), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_476), .B(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_476), .B(n_568), .Y(n_676) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx3_ASAP7_75t_L g533 ( .A(n_477), .Y(n_533) );
OAI31xp33_ASAP7_75t_L g715 ( .A1(n_487), .A2(n_636), .A3(n_643), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_498), .Y(n_487) );
AND2x2_ASAP7_75t_L g519 ( .A(n_488), .B(n_520), .Y(n_519) );
NAND2x1_ASAP7_75t_SL g538 ( .A(n_488), .B(n_539), .Y(n_538) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_488), .Y(n_625) );
AND2x2_ASAP7_75t_L g630 ( .A(n_488), .B(n_541), .Y(n_630) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_489), .A2(n_543), .B(n_545), .C(n_548), .Y(n_542) );
OR2x2_ASAP7_75t_L g559 ( .A(n_489), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g572 ( .A(n_489), .Y(n_572) );
AND2x2_ASAP7_75t_L g578 ( .A(n_489), .B(n_521), .Y(n_578) );
INVx2_ASAP7_75t_L g596 ( .A(n_489), .Y(n_596) );
AND2x2_ASAP7_75t_L g607 ( .A(n_489), .B(n_561), .Y(n_607) );
AND2x2_ASAP7_75t_L g639 ( .A(n_489), .B(n_597), .Y(n_639) );
AND2x2_ASAP7_75t_L g643 ( .A(n_489), .B(n_566), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_489), .B(n_498), .Y(n_648) );
AND2x2_ASAP7_75t_L g682 ( .A(n_489), .B(n_683), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_489), .B(n_585), .Y(n_716) );
OR2x6_ASAP7_75t_L g489 ( .A(n_490), .B(n_496), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_498), .B(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g624 ( .A(n_498), .Y(n_624) );
AND2x2_ASAP7_75t_L g686 ( .A(n_498), .B(n_607), .Y(n_686) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_510), .Y(n_498) );
OR2x2_ASAP7_75t_L g540 ( .A(n_499), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g550 ( .A(n_499), .B(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_499), .B(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g658 ( .A(n_499), .Y(n_658) );
AND2x2_ASAP7_75t_L g675 ( .A(n_499), .B(n_521), .Y(n_675) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g566 ( .A(n_500), .B(n_510), .Y(n_566) );
AND2x2_ASAP7_75t_L g595 ( .A(n_500), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g606 ( .A(n_500), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_500), .B(n_561), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_507), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_505), .B(n_506), .Y(n_503) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g520 ( .A(n_511), .B(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g541 ( .A(n_511), .Y(n_541) );
AND2x2_ASAP7_75t_L g597 ( .A(n_511), .B(n_561), .Y(n_597) );
INVx1_ASAP7_75t_L g699 ( .A(n_519), .Y(n_699) );
INVx1_ASAP7_75t_L g703 ( .A(n_520), .Y(n_703) );
INVx2_ASAP7_75t_L g561 ( .A(n_521), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_531), .B(n_534), .Y(n_530) );
INVx1_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_532), .B(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_532), .B(n_637), .Y(n_695) );
OR2x2_ASAP7_75t_L g536 ( .A(n_533), .B(n_534), .Y(n_536) );
INVx1_ASAP7_75t_SL g588 ( .A(n_533), .Y(n_588) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AOI221xp5_ASAP7_75t_L g591 ( .A1(n_539), .A2(n_592), .B1(n_594), .B2(n_598), .C(n_599), .Y(n_591) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g619 ( .A(n_540), .B(n_583), .Y(n_619) );
INVx2_ASAP7_75t_L g551 ( .A(n_541), .Y(n_551) );
INVx1_ASAP7_75t_L g577 ( .A(n_541), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_541), .B(n_561), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_541), .B(n_564), .Y(n_671) );
INVx1_ASAP7_75t_L g679 ( .A(n_541), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_543), .B(n_547), .Y(n_593) );
AND2x4_ASAP7_75t_L g568 ( .A(n_544), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g681 ( .A(n_547), .B(n_637), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_552), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_550), .B(n_582), .Y(n_581) );
INVxp67_ASAP7_75t_L g689 ( .A(n_551), .Y(n_689) );
INVxp67_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
INVx1_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g589 ( .A(n_555), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g661 ( .A(n_555), .B(n_637), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_555), .B(n_574), .Y(n_667) );
AOI322xp5_ASAP7_75t_L g621 ( .A1(n_556), .A2(n_590), .A3(n_597), .B1(n_622), .B2(n_625), .C1(n_626), .C2(n_628), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_556), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OR2x2_ASAP7_75t_L g687 ( .A(n_559), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g633 ( .A(n_560), .Y(n_633) );
INVx2_ASAP7_75t_L g564 ( .A(n_561), .Y(n_564) );
INVx1_ASAP7_75t_L g623 ( .A(n_561), .Y(n_623) );
CKINVDCx16_ASAP7_75t_R g570 ( .A(n_562), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
AND2x2_ASAP7_75t_L g659 ( .A(n_564), .B(n_572), .Y(n_659) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g571 ( .A(n_566), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g614 ( .A(n_566), .B(n_607), .Y(n_614) );
AND2x2_ASAP7_75t_L g618 ( .A(n_566), .B(n_578), .Y(n_618) );
OAI21xp33_ASAP7_75t_SL g628 ( .A1(n_567), .A2(n_629), .B(n_631), .Y(n_628) );
OAI22xp33_ASAP7_75t_L g698 ( .A1(n_567), .A2(n_699), .B1(n_700), .B2(n_702), .Y(n_698) );
INVx3_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g573 ( .A(n_568), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_568), .B(n_588), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_570), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
INVx1_ASAP7_75t_L g710 ( .A(n_577), .Y(n_710) );
INVx4_ASAP7_75t_L g583 ( .A(n_578), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_578), .B(n_605), .Y(n_653) );
INVx1_ASAP7_75t_SL g665 ( .A(n_579), .Y(n_665) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NOR2xp67_ASAP7_75t_L g678 ( .A(n_583), .B(n_679), .Y(n_678) );
OAI211xp5_ASAP7_75t_SL g584 ( .A1(n_585), .A2(n_586), .B(n_591), .C(n_608), .Y(n_584) );
OAI221xp5_ASAP7_75t_SL g704 ( .A1(n_586), .A2(n_624), .B1(n_703), .B2(n_705), .C(n_707), .Y(n_704) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_588), .B(n_701), .Y(n_700) );
OAI31xp33_ASAP7_75t_L g680 ( .A1(n_589), .A2(n_666), .A3(n_681), .B(n_682), .Y(n_680) );
INVx1_ASAP7_75t_L g620 ( .A(n_590), .Y(n_620) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
INVx1_ASAP7_75t_L g670 ( .A(n_595), .Y(n_670) );
AND2x2_ASAP7_75t_L g683 ( .A(n_597), .B(n_606), .Y(n_683) );
AOI21xp33_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_601), .B(n_603), .Y(n_599) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
INVxp67_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_607), .B(n_710), .Y(n_709) );
OAI21xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B(n_614), .Y(n_608) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OAI221xp5_ASAP7_75t_SL g615 ( .A1(n_616), .A2(n_617), .B1(n_619), .B2(n_620), .C(n_621), .Y(n_615) );
A2O1A1Ixp33_ASAP7_75t_L g684 ( .A1(n_616), .A2(n_685), .B(n_687), .C(n_690), .Y(n_684) );
CKINVDCx16_ASAP7_75t_R g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_619), .B(n_669), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx1_ASAP7_75t_L g646 ( .A(n_627), .Y(n_646) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g632 ( .A(n_630), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g674 ( .A(n_630), .B(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OAI211xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_638), .B(n_640), .C(n_649), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g711 ( .A1(n_638), .A2(n_648), .B1(n_712), .B2(n_713), .C(n_715), .Y(n_711) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_643), .B1(n_644), .B2(n_647), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OAI21xp5_ASAP7_75t_SL g649 ( .A1(n_650), .A2(n_651), .B(n_652), .Y(n_649) );
INVx1_ASAP7_75t_SL g712 ( .A(n_651), .Y(n_712) );
INVxp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NOR4xp25_ASAP7_75t_L g654 ( .A(n_655), .B(n_684), .C(n_704), .D(n_711), .Y(n_654) );
OAI211xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_660), .B(n_662), .C(n_680), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
INVxp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
O2A1O1Ixp33_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_666), .B(n_668), .C(n_672), .Y(n_662) );
INVx1_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g691 ( .A(n_669), .Y(n_691) );
OR2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
OR2x2_ASAP7_75t_L g702 ( .A(n_670), .B(n_703), .Y(n_702) );
OAI21xp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_676), .B(n_677), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_692), .B1(n_694), .B2(n_696), .C(n_698), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVxp67_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_701), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
endmodule