module fake_jpeg_31111_n_47 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_47);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_47;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_0),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_20),
.Y(n_28)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_18),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_25),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_30),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_24),
.A2(n_20),
.B1(n_21),
.B2(n_17),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_19),
.C(n_21),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_SL g37 ( 
.A(n_31),
.B(n_32),
.Y(n_37)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_35),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_4),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_SL g39 ( 
.A(n_31),
.B(n_2),
.C(n_3),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_3),
.B(n_4),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_33),
.B1(n_30),
.B2(n_5),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_41),
.B(n_5),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_6),
.B1(n_36),
.B2(n_17),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_44),
.C(n_6),
.Y(n_45)
);

A2O1A1O1Ixp25_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_7),
.B(n_9),
.C(n_12),
.D(n_13),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_16),
.Y(n_47)
);


endmodule