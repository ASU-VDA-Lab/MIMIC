module fake_ibex_1352_n_1203 (n_151, n_147, n_85, n_167, n_128, n_208, n_234, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_8, n_118, n_224, n_183, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_61, n_201, n_14, n_0, n_239, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_80, n_172, n_215, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_92, n_144, n_170, n_213, n_101, n_190, n_113, n_138, n_230, n_96, n_185, n_68, n_117, n_214, n_238, n_79, n_81, n_35, n_159, n_202, n_231, n_158, n_211, n_218, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_19, n_228, n_1203);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_208;
input n_234;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_8;
input n_118;
input n_224;
input n_183;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_61;
input n_201;
input n_14;
input n_0;
input n_239;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_80;
input n_172;
input n_215;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_213;
input n_101;
input n_190;
input n_113;
input n_138;
input n_230;
input n_96;
input n_185;
input n_68;
input n_117;
input n_214;
input n_238;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_218;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_19;
input n_228;

output n_1203;

wire n_1084;
wire n_599;
wire n_778;
wire n_822;
wire n_1042;
wire n_507;
wire n_743;
wire n_1148;
wire n_540;
wire n_754;
wire n_395;
wire n_1104;
wire n_1011;
wire n_992;
wire n_1060;
wire n_756;
wire n_529;
wire n_389;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_1090;
wire n_1110;
wire n_946;
wire n_1196;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_1182;
wire n_926;
wire n_1097;
wire n_1079;
wire n_1031;
wire n_1143;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_510;
wire n_845;
wire n_947;
wire n_972;
wire n_1100;
wire n_446;
wire n_350;
wire n_981;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_1067;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_1080;
wire n_1162;
wire n_1199;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_1125;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_432;
wire n_1034;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_457;
wire n_412;
wire n_357;
wire n_494;
wire n_959;
wire n_336;
wire n_930;
wire n_258;
wire n_861;
wire n_1018;
wire n_1044;
wire n_1106;
wire n_1129;
wire n_449;
wire n_1138;
wire n_547;
wire n_1134;
wire n_727;
wire n_1131;
wire n_1077;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_1174;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_1147;
wire n_542;
wire n_900;
wire n_376;
wire n_1098;
wire n_377;
wire n_584;
wire n_1189;
wire n_531;
wire n_647;
wire n_1187;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_708;
wire n_375;
wire n_317;
wire n_280;
wire n_340;
wire n_698;
wire n_901;
wire n_1096;
wire n_667;
wire n_884;
wire n_1061;
wire n_682;
wire n_850;
wire n_1166;
wire n_1181;
wire n_1140;
wire n_326;
wire n_327;
wire n_879;
wire n_1056;
wire n_723;
wire n_270;
wire n_1144;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_470;
wire n_276;
wire n_339;
wire n_770;
wire n_965;
wire n_348;
wire n_1109;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_671;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_1051;
wire n_854;
wire n_1008;
wire n_1193;
wire n_458;
wire n_244;
wire n_1053;
wire n_1112;
wire n_343;
wire n_310;
wire n_714;
wire n_1076;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_1172;
wire n_1099;
wire n_598;
wire n_825;
wire n_740;
wire n_1169;
wire n_386;
wire n_549;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_1201;
wire n_400;
wire n_306;
wire n_550;
wire n_736;
wire n_1055;
wire n_673;
wire n_732;
wire n_832;
wire n_798;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_1103;
wire n_1161;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_1177;
wire n_1068;
wire n_1057;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_1184;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_1195;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_1141;
wire n_523;
wire n_694;
wire n_787;
wire n_1075;
wire n_1136;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_1197;
wire n_574;
wire n_1168;
wire n_289;
wire n_716;
wire n_865;
wire n_1130;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_1179;
wire n_1192;
wire n_933;
wire n_1081;
wire n_1153;
wire n_279;
wire n_1037;
wire n_374;
wire n_464;
wire n_669;
wire n_538;
wire n_838;
wire n_987;
wire n_1155;
wire n_750;
wire n_1021;
wire n_746;
wire n_1188;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_1117;
wire n_1191;
wire n_1101;
wire n_518;
wire n_367;
wire n_1052;
wire n_852;
wire n_789;
wire n_1133;
wire n_880;
wire n_654;
wire n_1083;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_1178;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_281;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_490;
wire n_407;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_1116;
wire n_623;
wire n_585;
wire n_1030;
wire n_1094;
wire n_1020;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_769;
wire n_487;
wire n_1082;
wire n_1137;
wire n_660;
wire n_524;
wire n_349;
wire n_849;
wire n_765;
wire n_857;
wire n_980;
wire n_454;
wire n_1070;
wire n_1074;
wire n_777;
wire n_1200;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_1120;
wire n_576;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_1180;
wire n_619;
wire n_1089;
wire n_536;
wire n_1124;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_246;
wire n_442;
wire n_858;
wire n_1064;
wire n_922;
wire n_1071;
wire n_1171;
wire n_438;
wire n_851;
wire n_1028;
wire n_1012;
wire n_993;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_1183;
wire n_253;
wire n_300;
wire n_1151;
wire n_1135;
wire n_973;
wire n_1146;
wire n_358;
wire n_771;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_999;
wire n_1038;
wire n_1092;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_1066;
wire n_245;
wire n_589;
wire n_571;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_1062;
wire n_847;
wire n_830;
wire n_1142;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_1072;
wire n_263;
wire n_1173;
wire n_1069;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_262;
wire n_433;
wire n_439;
wire n_299;
wire n_704;
wire n_949;
wire n_1007;
wire n_1126;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_837;
wire n_797;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_699;
wire n_1063;
wire n_351;
wire n_456;
wire n_368;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_1115;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_1054;
wire n_672;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_553;
wire n_554;
wire n_1078;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_1170;
wire n_605;
wire n_539;
wire n_354;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_1049;
wire n_1086;
wire n_763;
wire n_1158;
wire n_745;
wire n_329;
wire n_1149;
wire n_447;
wire n_1176;
wire n_940;
wire n_444;
wire n_562;
wire n_564;
wire n_506;
wire n_868;
wire n_546;
wire n_788;
wire n_1202;
wire n_795;
wire n_1065;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_1160;
wire n_615;
wire n_512;
wire n_950;
wire n_685;
wire n_1026;
wire n_397;
wire n_366;
wire n_283;
wire n_803;
wire n_894;
wire n_1118;
wire n_1033;
wire n_692;
wire n_627;
wire n_990;
wire n_1198;
wire n_709;
wire n_322;
wire n_499;
wire n_888;
wire n_1087;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_1114;
wire n_409;
wire n_1093;
wire n_582;
wire n_978;
wire n_818;
wire n_1167;
wire n_653;
wire n_579;
wire n_843;
wire n_899;
wire n_1059;
wire n_1019;
wire n_902;
wire n_332;
wire n_799;
wire n_1190;
wire n_517;
wire n_817;
wire n_744;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_1107;
wire n_381;
wire n_1073;
wire n_1108;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_1111;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_285;
wire n_247;
wire n_320;
wire n_379;
wire n_1128;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_268;
wire n_440;
wire n_955;
wire n_385;
wire n_414;
wire n_342;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_1145;
wire n_977;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_1113;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_1164;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_1175;
wire n_485;
wire n_1139;
wire n_870;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_1159;
wire n_1119;
wire n_903;
wire n_1154;
wire n_519;
wire n_345;
wire n_408;
wire n_1085;
wire n_361;
wire n_1095;
wire n_455;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_1091;
wire n_885;
wire n_588;
wire n_513;
wire n_877;
wire n_1121;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_1088;
wire n_896;
wire n_528;
wire n_1005;
wire n_1102;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_1150;
wire n_462;
wire n_1194;
wire n_450;
wire n_302;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_1165;
wire n_1185;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_1122;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_912;
wire n_921;
wire n_890;
wire n_874;
wire n_1105;
wire n_1058;
wire n_1163;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_1123;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_1000;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_298;
wire n_587;
wire n_1035;
wire n_760;
wire n_1157;
wire n_751;
wire n_806;
wire n_1127;
wire n_932;
wire n_1186;
wire n_657;
wire n_764;
wire n_1156;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_380;
wire n_749;
wire n_866;
wire n_559;
wire n_425;
wire n_1050;

INVx1_ASAP7_75t_L g240 ( 
.A(n_17),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_103),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_16),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_133),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_55),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_114),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_104),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_153),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_192),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_124),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_142),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_202),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_185),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_19),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_101),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_211),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_172),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_227),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_176),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_187),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_175),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_16),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_77),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_146),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_166),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_140),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_205),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_96),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_74),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_134),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_137),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_144),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_182),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_81),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_58),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_191),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_105),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_48),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_179),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_173),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_229),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_148),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_222),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_167),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_207),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_215),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_197),
.B(n_149),
.Y(n_287)
);

INVxp33_ASAP7_75t_SL g288 ( 
.A(n_165),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_95),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_L g290 ( 
.A(n_40),
.B(n_169),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_111),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_138),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_13),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_69),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_107),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_131),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_231),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_214),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_112),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_157),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_0),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_125),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_12),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_35),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_42),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_178),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_75),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_2),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_45),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_27),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_39),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_35),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_200),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_181),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_232),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_19),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_108),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_129),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_230),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_186),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_128),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_71),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_92),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_87),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_59),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_151),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_139),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_109),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_118),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_83),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_52),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_110),
.Y(n_332)
);

INVxp33_ASAP7_75t_SL g333 ( 
.A(n_117),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_189),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_213),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_115),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_180),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_209),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_99),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_237),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_206),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_122),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_60),
.Y(n_343)
);

BUFx2_ASAP7_75t_SL g344 ( 
.A(n_4),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_106),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_3),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_216),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_53),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_84),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_204),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_141),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_210),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_198),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_136),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_162),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_44),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_12),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_65),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_102),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_159),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_226),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_89),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_15),
.B(n_201),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_90),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_194),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_11),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_150),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_79),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_223),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_40),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_127),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_120),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_97),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_123),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_155),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_64),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_2),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_60),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_228),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_195),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_3),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_235),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_170),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_158),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_177),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_184),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_29),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_160),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_220),
.Y(n_389)
);

INVxp33_ASAP7_75t_L g390 ( 
.A(n_21),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g391 ( 
.A(n_217),
.B(n_121),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_11),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_212),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_113),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_41),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_66),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_79),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_27),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_218),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_31),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_233),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_23),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_219),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_196),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_75),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_52),
.Y(n_406)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_168),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_224),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_71),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_143),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_100),
.Y(n_411)
);

NOR2xp67_ASAP7_75t_L g412 ( 
.A(n_20),
.B(n_47),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_308),
.B(n_1),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_341),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_319),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_390),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_251),
.B(n_1),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_319),
.Y(n_418)
);

NAND2xp33_ASAP7_75t_L g419 ( 
.A(n_254),
.B(n_80),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_401),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_319),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_319),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_346),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_346),
.B(n_5),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_358),
.Y(n_425)
);

INVx5_ASAP7_75t_L g426 ( 
.A(n_375),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_358),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_375),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_375),
.Y(n_429)
);

OAI22x1_ASAP7_75t_R g430 ( 
.A1(n_242),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_259),
.B(n_6),
.Y(n_431)
);

INVx5_ASAP7_75t_L g432 ( 
.A(n_375),
.Y(n_432)
);

BUFx8_ASAP7_75t_L g433 ( 
.A(n_298),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_390),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_381),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_240),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_254),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_267),
.B(n_8),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_263),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_254),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_296),
.B(n_10),
.Y(n_441)
);

OAI21x1_ASAP7_75t_L g442 ( 
.A1(n_256),
.A2(n_85),
.B(n_82),
.Y(n_442)
);

INVx5_ASAP7_75t_L g443 ( 
.A(n_247),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_267),
.B(n_10),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_257),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_247),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_254),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_263),
.A2(n_387),
.B1(n_325),
.B2(n_245),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_270),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_325),
.B(n_13),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_247),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_317),
.B(n_14),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_270),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_331),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_282),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_262),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_289),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_280),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_275),
.Y(n_459)
);

INVx6_ASAP7_75t_L g460 ( 
.A(n_277),
.Y(n_460)
);

INVx5_ASAP7_75t_L g461 ( 
.A(n_277),
.Y(n_461)
);

AND2x6_ASAP7_75t_L g462 ( 
.A(n_317),
.B(n_86),
.Y(n_462)
);

AND2x6_ASAP7_75t_L g463 ( 
.A(n_354),
.B(n_88),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_331),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_294),
.Y(n_465)
);

AND2x6_ASAP7_75t_L g466 ( 
.A(n_354),
.B(n_91),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_280),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_303),
.Y(n_468)
);

OA21x2_ASAP7_75t_L g469 ( 
.A1(n_292),
.A2(n_94),
.B(n_93),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_292),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_277),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_331),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_323),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_323),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_347),
.Y(n_475)
);

INVx6_ASAP7_75t_L g476 ( 
.A(n_331),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_400),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_400),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_387),
.B(n_18),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_296),
.B(n_18),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_304),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_400),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_400),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_305),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_360),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_307),
.Y(n_486)
);

OA21x2_ASAP7_75t_L g487 ( 
.A1(n_380),
.A2(n_132),
.B(n_238),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_405),
.Y(n_488)
);

CKINVDCx11_ASAP7_75t_R g489 ( 
.A(n_244),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_380),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_405),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_399),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_388),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_309),
.B(n_24),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_405),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_408),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_405),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_424),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_446),
.B(n_260),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_438),
.B(n_399),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_415),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_446),
.B(n_250),
.Y(n_502)
);

NAND3xp33_ASAP7_75t_L g503 ( 
.A(n_414),
.B(n_322),
.C(n_301),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_438),
.Y(n_504)
);

OR2x6_ASAP7_75t_L g505 ( 
.A(n_416),
.B(n_344),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_415),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_446),
.B(n_310),
.Y(n_507)
);

AO22x2_ASAP7_75t_L g508 ( 
.A1(n_434),
.A2(n_448),
.B1(n_438),
.B2(n_444),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_451),
.B(n_311),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_444),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_444),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_418),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_418),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_452),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_418),
.Y(n_515)
);

NAND2xp33_ASAP7_75t_L g516 ( 
.A(n_466),
.B(n_287),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_418),
.Y(n_517)
);

INVx5_ASAP7_75t_L g518 ( 
.A(n_466),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_421),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_421),
.Y(n_520)
);

INVx4_ASAP7_75t_SL g521 ( 
.A(n_462),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_451),
.B(n_411),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_451),
.B(n_260),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_421),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_471),
.B(n_261),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_445),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_422),
.Y(n_527)
);

NAND2xp33_ASAP7_75t_L g528 ( 
.A(n_466),
.B(n_462),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_471),
.B(n_411),
.Y(n_529)
);

INVxp67_ASAP7_75t_SL g530 ( 
.A(n_441),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_471),
.B(n_261),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_427),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_422),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_445),
.Y(n_534)
);

NAND3x1_ASAP7_75t_L g535 ( 
.A(n_455),
.B(n_269),
.C(n_244),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_449),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_460),
.B(n_241),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_428),
.Y(n_538)
);

BUFx10_ASAP7_75t_L g539 ( 
.A(n_460),
.Y(n_539)
);

INVx1_ASAP7_75t_SL g540 ( 
.A(n_439),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_453),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_453),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_443),
.B(n_264),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g544 ( 
.A(n_420),
.B(n_456),
.Y(n_544)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_462),
.Y(n_545)
);

OAI22xp33_ASAP7_75t_L g546 ( 
.A1(n_485),
.A2(n_269),
.B1(n_293),
.B2(n_312),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_458),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_458),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_428),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_461),
.B(n_243),
.Y(n_550)
);

INVxp33_ASAP7_75t_SL g551 ( 
.A(n_457),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_467),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_470),
.Y(n_553)
);

BUFx10_ASAP7_75t_L g554 ( 
.A(n_496),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_428),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_473),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_473),
.Y(n_557)
);

BUFx4f_ASAP7_75t_L g558 ( 
.A(n_441),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_474),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_461),
.B(n_264),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_475),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_463),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_436),
.B(n_278),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_461),
.B(n_246),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_429),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_429),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_429),
.Y(n_567)
);

OR2x6_ASAP7_75t_L g568 ( 
.A(n_480),
.B(n_412),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_429),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_426),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_426),
.Y(n_571)
);

AO21x2_ASAP7_75t_L g572 ( 
.A1(n_442),
.A2(n_363),
.B(n_249),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_426),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_426),
.Y(n_574)
);

NOR3xp33_ASAP7_75t_L g575 ( 
.A(n_450),
.B(n_402),
.C(n_348),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_459),
.B(n_248),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_465),
.B(n_252),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_468),
.B(n_253),
.Y(n_578)
);

INVx6_ASAP7_75t_L g579 ( 
.A(n_433),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_431),
.B(n_255),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_432),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_490),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_433),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_432),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_466),
.A2(n_316),
.B1(n_357),
.B2(n_356),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_432),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_SL g587 ( 
.A(n_480),
.B(n_268),
.Y(n_587)
);

NAND2xp33_ASAP7_75t_L g588 ( 
.A(n_466),
.B(n_391),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_492),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_433),
.B(n_481),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_492),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_484),
.B(n_486),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_423),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_425),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_432),
.Y(n_595)
);

AND2x2_ASAP7_75t_SL g596 ( 
.A(n_417),
.B(n_258),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_432),
.B(n_265),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_437),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_437),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_435),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_494),
.A2(n_368),
.B1(n_370),
.B2(n_366),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_437),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_413),
.B(n_343),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_476),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_476),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_479),
.Y(n_606)
);

AO22x2_ASAP7_75t_L g607 ( 
.A1(n_430),
.A2(n_395),
.B1(n_396),
.B2(n_377),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_472),
.Y(n_608)
);

AO22x2_ASAP7_75t_L g609 ( 
.A1(n_472),
.A2(n_409),
.B1(n_271),
.B2(n_272),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_440),
.Y(n_610)
);

BUFx10_ASAP7_75t_L g611 ( 
.A(n_476),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_472),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_469),
.A2(n_333),
.B1(n_288),
.B2(n_266),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_483),
.Y(n_614)
);

NAND3xp33_ASAP7_75t_L g615 ( 
.A(n_419),
.B(n_378),
.C(n_376),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_483),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_469),
.A2(n_333),
.B1(n_288),
.B2(n_273),
.Y(n_617)
);

INVxp67_ASAP7_75t_L g618 ( 
.A(n_442),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_440),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_493),
.A2(n_279),
.B1(n_286),
.B2(n_268),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_440),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_491),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_491),
.B(n_392),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_487),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_590),
.B(n_335),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_575),
.A2(n_279),
.B1(n_306),
.B2(n_286),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_575),
.A2(n_306),
.B1(n_318),
.B2(n_313),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_530),
.B(n_382),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_530),
.B(n_407),
.Y(n_629)
);

OR2x2_ASAP7_75t_L g630 ( 
.A(n_540),
.B(n_397),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_606),
.B(n_487),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_563),
.B(n_398),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_510),
.B(n_487),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_505),
.B(n_313),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_511),
.B(n_274),
.Y(n_635)
);

BUFx12f_ASAP7_75t_L g636 ( 
.A(n_505),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_614),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_514),
.B(n_281),
.Y(n_638)
);

NOR3xp33_ASAP7_75t_L g639 ( 
.A(n_546),
.B(n_489),
.C(n_406),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_539),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_596),
.A2(n_318),
.B1(n_345),
.B2(n_337),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_544),
.B(n_353),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_504),
.B(n_291),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_504),
.B(n_295),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_508),
.A2(n_345),
.B1(n_355),
.B2(n_337),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_507),
.B(n_361),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_502),
.B(n_276),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_603),
.B(n_489),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_553),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_596),
.A2(n_372),
.B1(n_385),
.B2(n_355),
.Y(n_650)
);

NAND3xp33_ASAP7_75t_SL g651 ( 
.A(n_620),
.B(n_385),
.C(n_372),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_499),
.B(n_283),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_523),
.B(n_284),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_SL g654 ( 
.A(n_545),
.B(n_404),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_525),
.B(n_285),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_508),
.A2(n_404),
.B1(n_293),
.B2(n_299),
.Y(n_656)
);

OR2x2_ASAP7_75t_SL g657 ( 
.A(n_607),
.B(n_535),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_531),
.B(n_300),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_508),
.A2(n_290),
.B1(n_302),
.B2(n_297),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_592),
.B(n_314),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_507),
.B(n_509),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_562),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_592),
.B(n_315),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_498),
.B(n_321),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_528),
.A2(n_419),
.B(n_326),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_509),
.A2(n_365),
.B1(n_324),
.B2(n_327),
.Y(n_666)
);

OAI22xp33_ASAP7_75t_L g667 ( 
.A1(n_546),
.A2(n_328),
.B1(n_329),
.B2(n_330),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_500),
.B(n_332),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_558),
.A2(n_601),
.B1(n_607),
.B2(n_585),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_500),
.B(n_336),
.Y(n_670)
);

INVxp67_ASAP7_75t_SL g671 ( 
.A(n_558),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_L g672 ( 
.A1(n_618),
.A2(n_342),
.B(n_338),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_561),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_539),
.B(n_583),
.Y(n_674)
);

AOI22xp5_ASAP7_75t_L g675 ( 
.A1(n_579),
.A2(n_349),
.B1(n_350),
.B2(n_351),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_SL g676 ( 
.A1(n_607),
.A2(n_393),
.B1(n_320),
.B2(n_334),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_522),
.B(n_362),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_568),
.B(n_25),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_537),
.B(n_339),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_580),
.B(n_340),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_580),
.B(n_503),
.Y(n_681)
);

O2A1O1Ixp33_ASAP7_75t_L g682 ( 
.A1(n_593),
.A2(n_410),
.B(n_403),
.C(n_386),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_522),
.B(n_352),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_529),
.B(n_359),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_532),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_529),
.B(n_367),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_551),
.B(n_383),
.Y(n_687)
);

OR2x6_ASAP7_75t_L g688 ( 
.A(n_579),
.B(n_364),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_554),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_594),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_543),
.B(n_560),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_587),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_600),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_518),
.B(n_389),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_518),
.B(n_394),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_576),
.B(n_369),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_576),
.B(n_371),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_609),
.A2(n_373),
.B1(n_374),
.B2(n_379),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_577),
.B(n_384),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_577),
.B(n_497),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_578),
.B(n_497),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_521),
.B(n_25),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_578),
.B(n_98),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_609),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_609),
.B(n_26),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_613),
.B(n_447),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_528),
.A2(n_495),
.B(n_488),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_613),
.B(n_447),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_526),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_534),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_617),
.B(n_454),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_536),
.Y(n_712)
);

NOR2xp67_ASAP7_75t_L g713 ( 
.A(n_623),
.B(n_28),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_516),
.A2(n_482),
.B1(n_478),
.B2(n_477),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_564),
.Y(n_715)
);

NAND2xp33_ASAP7_75t_L g716 ( 
.A(n_617),
.B(n_615),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_624),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_541),
.B(n_542),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_550),
.B(n_116),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_550),
.B(n_119),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_547),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_548),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_552),
.Y(n_723)
);

NAND2xp33_ASAP7_75t_L g724 ( 
.A(n_570),
.B(n_454),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_588),
.B(n_126),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_556),
.Y(n_726)
);

AND2x6_ASAP7_75t_SL g727 ( 
.A(n_557),
.B(n_559),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_588),
.A2(n_582),
.B1(n_591),
.B2(n_589),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_611),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_604),
.Y(n_730)
);

INVx5_ASAP7_75t_L g731 ( 
.A(n_616),
.Y(n_731)
);

OR2x4_ASAP7_75t_L g732 ( 
.A(n_608),
.B(n_612),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_572),
.B(n_464),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_572),
.A2(n_464),
.B1(n_30),
.B2(n_31),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_597),
.B(n_464),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_622),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_571),
.B(n_29),
.Y(n_737)
);

INVx5_ASAP7_75t_L g738 ( 
.A(n_605),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_669),
.A2(n_573),
.B1(n_581),
.B2(n_584),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_628),
.B(n_574),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_628),
.B(n_574),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_629),
.B(n_586),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_718),
.Y(n_743)
);

OAI21xp5_ASAP7_75t_L g744 ( 
.A1(n_631),
.A2(n_595),
.B(n_586),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_634),
.B(n_32),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_631),
.A2(n_595),
.B(n_501),
.Y(n_746)
);

O2A1O1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_667),
.A2(n_619),
.B(n_610),
.C(n_602),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_688),
.B(n_33),
.Y(n_748)
);

XOR2xp5_ASAP7_75t_L g749 ( 
.A(n_689),
.B(n_33),
.Y(n_749)
);

O2A1O1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_659),
.A2(n_602),
.B(n_599),
.C(n_598),
.Y(n_750)
);

OAI21xp33_ASAP7_75t_L g751 ( 
.A1(n_642),
.A2(n_654),
.B(n_661),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_629),
.B(n_34),
.Y(n_752)
);

AND2x4_ASAP7_75t_L g753 ( 
.A(n_688),
.B(n_671),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_726),
.B(n_36),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_681),
.B(n_37),
.Y(n_755)
);

OAI321xp33_ASAP7_75t_L g756 ( 
.A1(n_659),
.A2(n_621),
.A3(n_569),
.B1(n_567),
.B2(n_566),
.C(n_565),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_723),
.B(n_38),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_691),
.A2(n_527),
.B(n_566),
.Y(n_758)
);

NAND2xp33_ASAP7_75t_SL g759 ( 
.A(n_634),
.B(n_38),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_688),
.A2(n_520),
.B1(n_565),
.B2(n_555),
.Y(n_760)
);

A2O1A1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_672),
.A2(n_697),
.B(n_690),
.C(n_703),
.Y(n_761)
);

BUFx8_ASAP7_75t_L g762 ( 
.A(n_636),
.Y(n_762)
);

NOR3xp33_ASAP7_75t_L g763 ( 
.A(n_651),
.B(n_506),
.C(n_512),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_630),
.B(n_41),
.Y(n_764)
);

AND2x2_ASAP7_75t_SL g765 ( 
.A(n_641),
.B(n_42),
.Y(n_765)
);

OA21x2_ASAP7_75t_L g766 ( 
.A1(n_672),
.A2(n_527),
.B(n_515),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_728),
.A2(n_520),
.B1(n_549),
.B2(n_538),
.Y(n_767)
);

A2O1A1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_725),
.A2(n_682),
.B(n_708),
.C(n_706),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_702),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_706),
.A2(n_533),
.B(n_517),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_693),
.B(n_43),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_708),
.A2(n_711),
.B(n_665),
.Y(n_772)
);

OAI21xp5_ASAP7_75t_L g773 ( 
.A1(n_707),
.A2(n_513),
.B(n_517),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_625),
.B(n_666),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_711),
.A2(n_644),
.B(n_643),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_729),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_643),
.A2(n_644),
.B(n_664),
.Y(n_777)
);

NOR2xp67_ASAP7_75t_L g778 ( 
.A(n_648),
.B(n_44),
.Y(n_778)
);

INVx8_ASAP7_75t_L g779 ( 
.A(n_702),
.Y(n_779)
);

A2O1A1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_709),
.A2(n_712),
.B(n_721),
.C(n_710),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_660),
.B(n_46),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_717),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_660),
.B(n_46),
.Y(n_783)
);

NOR3xp33_ASAP7_75t_L g784 ( 
.A(n_639),
.B(n_519),
.C(n_538),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_663),
.B(n_47),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_663),
.B(n_49),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_646),
.B(n_49),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_650),
.B(n_50),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_635),
.B(n_51),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_638),
.B(n_51),
.Y(n_790)
);

OA22x2_ASAP7_75t_L g791 ( 
.A1(n_656),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_685),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_687),
.B(n_56),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_627),
.B(n_57),
.Y(n_794)
);

AO22x1_ASAP7_75t_L g795 ( 
.A1(n_705),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_795)
);

NOR3xp33_ASAP7_75t_L g796 ( 
.A(n_676),
.B(n_61),
.C(n_62),
.Y(n_796)
);

AOI221xp5_ASAP7_75t_L g797 ( 
.A1(n_626),
.A2(n_524),
.B1(n_64),
.B2(n_65),
.C(n_66),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_662),
.B(n_63),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_645),
.B(n_63),
.Y(n_799)
);

OR2x6_ASAP7_75t_L g800 ( 
.A(n_640),
.B(n_67),
.Y(n_800)
);

O2A1O1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_678),
.A2(n_68),
.B(n_69),
.C(n_70),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_668),
.B(n_70),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_670),
.B(n_72),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_674),
.B(n_72),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_698),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_680),
.Y(n_806)
);

O2A1O1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_670),
.A2(n_73),
.B(n_77),
.C(n_78),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_736),
.Y(n_808)
);

A2O1A1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_722),
.A2(n_78),
.B(n_130),
.C(n_135),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_696),
.B(n_239),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_727),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_699),
.B(n_234),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_L g813 ( 
.A1(n_717),
.A2(n_145),
.B1(n_147),
.B2(n_152),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_734),
.A2(n_677),
.B(n_714),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_675),
.B(n_154),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_652),
.B(n_156),
.Y(n_816)
);

A2O1A1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_677),
.A2(n_161),
.B(n_163),
.C(n_164),
.Y(n_817)
);

OR2x6_ASAP7_75t_L g818 ( 
.A(n_715),
.B(n_171),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_647),
.A2(n_174),
.B1(n_183),
.B2(n_188),
.Y(n_819)
);

AO21x1_ASAP7_75t_L g820 ( 
.A1(n_719),
.A2(n_190),
.B(n_193),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_700),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_701),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_731),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_653),
.A2(n_655),
.B(n_658),
.Y(n_824)
);

AOI21x1_ASAP7_75t_L g825 ( 
.A1(n_735),
.A2(n_199),
.B(n_203),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_683),
.B(n_225),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_684),
.B(n_221),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_649),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_686),
.B(n_208),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_679),
.B(n_673),
.Y(n_830)
);

BUFx3_ASAP7_75t_L g831 ( 
.A(n_732),
.Y(n_831)
);

NAND3xp33_ASAP7_75t_L g832 ( 
.A(n_713),
.B(n_737),
.C(n_720),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_657),
.A2(n_637),
.B1(n_731),
.B2(n_730),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_731),
.B(n_694),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_731),
.B(n_695),
.Y(n_835)
);

BUFx2_ASAP7_75t_L g836 ( 
.A(n_738),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_724),
.A2(n_528),
.B(n_631),
.Y(n_837)
);

INVxp67_ASAP7_75t_L g838 ( 
.A(n_738),
.Y(n_838)
);

CKINVDCx10_ASAP7_75t_R g839 ( 
.A(n_738),
.Y(n_839)
);

AOI21xp33_ASAP7_75t_L g840 ( 
.A1(n_692),
.A2(n_642),
.B(n_716),
.Y(n_840)
);

O2A1O1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_667),
.A2(n_659),
.B(n_716),
.C(n_669),
.Y(n_841)
);

OAI22x1_ASAP7_75t_L g842 ( 
.A1(n_641),
.A2(n_650),
.B1(n_634),
.B2(n_656),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_631),
.A2(n_528),
.B(n_633),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_631),
.A2(n_528),
.B(n_633),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_704),
.A2(n_530),
.B1(n_558),
.B2(n_669),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_L g846 ( 
.A1(n_631),
.A2(n_618),
.B(n_633),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_631),
.A2(n_528),
.B(n_633),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_672),
.A2(n_631),
.B(n_681),
.C(n_697),
.Y(n_848)
);

OAI21xp5_ASAP7_75t_L g849 ( 
.A1(n_733),
.A2(n_618),
.B(n_631),
.Y(n_849)
);

AO32x2_ASAP7_75t_L g850 ( 
.A1(n_845),
.A2(n_805),
.A3(n_833),
.B1(n_819),
.B2(n_767),
.Y(n_850)
);

AOI221xp5_ASAP7_75t_SL g851 ( 
.A1(n_841),
.A2(n_848),
.B1(n_775),
.B2(n_761),
.C(n_768),
.Y(n_851)
);

OR2x2_ASAP7_75t_L g852 ( 
.A(n_743),
.B(n_794),
.Y(n_852)
);

CKINVDCx11_ASAP7_75t_R g853 ( 
.A(n_776),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_SL g854 ( 
.A1(n_748),
.A2(n_818),
.B(n_849),
.Y(n_854)
);

A2O1A1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_777),
.A2(n_824),
.B(n_755),
.C(n_793),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_SL g856 ( 
.A1(n_748),
.A2(n_799),
.B(n_796),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_806),
.B(n_764),
.Y(n_857)
);

AO22x2_ASAP7_75t_L g858 ( 
.A1(n_788),
.A2(n_745),
.B1(n_769),
.B2(n_749),
.Y(n_858)
);

INVx4_ASAP7_75t_L g859 ( 
.A(n_779),
.Y(n_859)
);

AO31x2_ASAP7_75t_L g860 ( 
.A1(n_820),
.A2(n_817),
.A3(n_809),
.B(n_837),
.Y(n_860)
);

AO32x2_ASAP7_75t_L g861 ( 
.A1(n_760),
.A2(n_813),
.A3(n_756),
.B1(n_791),
.B2(n_750),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_744),
.A2(n_746),
.B(n_814),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_765),
.B(n_800),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_758),
.A2(n_812),
.B(n_810),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_800),
.Y(n_865)
);

OAI21xp33_ASAP7_75t_L g866 ( 
.A1(n_751),
.A2(n_783),
.B(n_781),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_762),
.Y(n_867)
);

O2A1O1Ixp5_ASAP7_75t_L g868 ( 
.A1(n_840),
.A2(n_816),
.B(n_814),
.C(n_787),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_780),
.A2(n_770),
.B(n_830),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_839),
.Y(n_870)
);

OAI21x1_ASAP7_75t_L g871 ( 
.A1(n_825),
.A2(n_773),
.B(n_766),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_826),
.A2(n_829),
.B(n_827),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_831),
.B(n_753),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_769),
.A2(n_818),
.B1(n_786),
.B2(n_785),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_753),
.B(n_811),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_823),
.B(n_778),
.Y(n_876)
);

CKINVDCx11_ASAP7_75t_R g877 ( 
.A(n_800),
.Y(n_877)
);

INVx1_ASAP7_75t_SL g878 ( 
.A(n_759),
.Y(n_878)
);

OAI21xp5_ASAP7_75t_L g879 ( 
.A1(n_739),
.A2(n_740),
.B(n_741),
.Y(n_879)
);

OR2x2_ASAP7_75t_L g880 ( 
.A(n_752),
.B(n_742),
.Y(n_880)
);

INVx1_ASAP7_75t_SL g881 ( 
.A(n_836),
.Y(n_881)
);

A2O1A1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_789),
.A2(n_790),
.B(n_747),
.C(n_807),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_762),
.Y(n_883)
);

CKINVDCx20_ASAP7_75t_R g884 ( 
.A(n_838),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_804),
.B(n_815),
.Y(n_885)
);

AO21x2_ASAP7_75t_L g886 ( 
.A1(n_832),
.A2(n_771),
.B(n_798),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_802),
.B(n_803),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_821),
.A2(n_822),
.B1(n_754),
.B2(n_757),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_782),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_801),
.B(n_792),
.Y(n_890)
);

OR2x2_ASAP7_75t_L g891 ( 
.A(n_828),
.B(n_795),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_784),
.A2(n_763),
.B(n_834),
.C(n_835),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_L g893 ( 
.A1(n_743),
.A2(n_530),
.B1(n_558),
.B2(n_748),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_743),
.B(n_530),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_743),
.A2(n_530),
.B1(n_558),
.B2(n_748),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_743),
.A2(n_530),
.B1(n_558),
.B2(n_748),
.Y(n_896)
);

AO32x2_ASAP7_75t_L g897 ( 
.A1(n_845),
.A2(n_659),
.A3(n_805),
.B1(n_833),
.B2(n_669),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_846),
.A2(n_528),
.B(n_849),
.Y(n_898)
);

OAI21xp33_ASAP7_75t_L g899 ( 
.A1(n_761),
.A2(n_774),
.B(n_848),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_743),
.B(n_530),
.Y(n_900)
);

OAI22x1_ASAP7_75t_L g901 ( 
.A1(n_748),
.A2(n_641),
.B1(n_650),
.B2(n_656),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_808),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_846),
.A2(n_528),
.B(n_849),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_841),
.A2(n_761),
.B(n_777),
.C(n_824),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_743),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_782),
.Y(n_906)
);

INVx4_ASAP7_75t_L g907 ( 
.A(n_779),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_SL g908 ( 
.A1(n_748),
.A2(n_669),
.B(n_656),
.Y(n_908)
);

O2A1O1Ixp5_ASAP7_75t_SL g909 ( 
.A1(n_840),
.A2(n_659),
.B(n_733),
.C(n_427),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_843),
.A2(n_847),
.B(n_844),
.Y(n_910)
);

INVx1_ASAP7_75t_SL g911 ( 
.A(n_748),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_846),
.A2(n_528),
.B(n_849),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_762),
.Y(n_913)
);

A2O1A1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_841),
.A2(n_761),
.B(n_777),
.C(n_824),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_743),
.B(n_632),
.Y(n_915)
);

NAND3xp33_ASAP7_75t_L g916 ( 
.A(n_761),
.B(n_716),
.C(n_797),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_743),
.Y(n_917)
);

AND3x4_ASAP7_75t_L g918 ( 
.A(n_796),
.B(n_639),
.C(n_634),
.Y(n_918)
);

BUFx4f_ASAP7_75t_L g919 ( 
.A(n_748),
.Y(n_919)
);

NAND2x1p5_ASAP7_75t_L g920 ( 
.A(n_748),
.B(n_776),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_846),
.A2(n_528),
.B(n_849),
.Y(n_921)
);

NAND3xp33_ASAP7_75t_L g922 ( 
.A(n_761),
.B(n_716),
.C(n_797),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_846),
.A2(n_528),
.B(n_849),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_743),
.A2(n_530),
.B1(n_558),
.B2(n_748),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_846),
.A2(n_528),
.B(n_849),
.Y(n_925)
);

A2O1A1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_841),
.A2(n_761),
.B(n_777),
.C(n_824),
.Y(n_926)
);

AO31x2_ASAP7_75t_L g927 ( 
.A1(n_820),
.A2(n_845),
.A3(n_848),
.B(n_772),
.Y(n_927)
);

CKINVDCx6p67_ASAP7_75t_R g928 ( 
.A(n_839),
.Y(n_928)
);

NAND3xp33_ASAP7_75t_L g929 ( 
.A(n_761),
.B(n_716),
.C(n_797),
.Y(n_929)
);

NOR2xp67_ASAP7_75t_L g930 ( 
.A(n_748),
.B(n_704),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_762),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_782),
.Y(n_932)
);

NAND3xp33_ASAP7_75t_L g933 ( 
.A(n_761),
.B(n_716),
.C(n_797),
.Y(n_933)
);

AO32x2_ASAP7_75t_L g934 ( 
.A1(n_845),
.A2(n_659),
.A3(n_805),
.B1(n_833),
.B2(n_669),
.Y(n_934)
);

OA21x2_ASAP7_75t_L g935 ( 
.A1(n_849),
.A2(n_733),
.B(n_846),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_743),
.B(n_632),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_808),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_808),
.Y(n_938)
);

OAI21xp33_ASAP7_75t_L g939 ( 
.A1(n_761),
.A2(n_774),
.B(n_848),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_743),
.B(n_632),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_806),
.B(n_648),
.Y(n_941)
);

AO31x2_ASAP7_75t_L g942 ( 
.A1(n_820),
.A2(n_845),
.A3(n_848),
.B(n_772),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_743),
.B(n_540),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_748),
.B(n_654),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_846),
.A2(n_528),
.B(n_849),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_SL g946 ( 
.A1(n_748),
.A2(n_704),
.B(n_818),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_743),
.B(n_530),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_743),
.B(n_530),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_762),
.Y(n_949)
);

OA22x2_ASAP7_75t_L g950 ( 
.A1(n_842),
.A2(n_650),
.B1(n_641),
.B2(n_656),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_748),
.B(n_654),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_743),
.B(n_632),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_748),
.A2(n_669),
.B1(n_765),
.B2(n_845),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_748),
.A2(n_669),
.B1(n_765),
.B2(n_845),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_843),
.A2(n_847),
.B(n_844),
.Y(n_955)
);

O2A1O1Ixp5_ASAP7_75t_SL g956 ( 
.A1(n_840),
.A2(n_659),
.B(n_733),
.C(n_427),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_748),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_743),
.B(n_632),
.Y(n_958)
);

CKINVDCx20_ASAP7_75t_R g959 ( 
.A(n_762),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_SL g960 ( 
.A1(n_748),
.A2(n_704),
.B(n_818),
.Y(n_960)
);

NAND2x1p5_ASAP7_75t_L g961 ( 
.A(n_748),
.B(n_776),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_806),
.B(n_648),
.Y(n_962)
);

INVx4_ASAP7_75t_L g963 ( 
.A(n_883),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_859),
.B(n_907),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_904),
.A2(n_926),
.B(n_914),
.Y(n_965)
);

AO21x2_ASAP7_75t_L g966 ( 
.A1(n_862),
.A2(n_955),
.B(n_910),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_943),
.B(n_915),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_898),
.A2(n_912),
.B(n_903),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_905),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_921),
.A2(n_925),
.B(n_923),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_911),
.Y(n_971)
);

OR3x4_ASAP7_75t_SL g972 ( 
.A(n_928),
.B(n_877),
.C(n_959),
.Y(n_972)
);

INVxp67_ASAP7_75t_L g973 ( 
.A(n_894),
.Y(n_973)
);

AND2x6_ASAP7_75t_L g974 ( 
.A(n_957),
.B(n_953),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_902),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_919),
.Y(n_976)
);

OR3x4_ASAP7_75t_SL g977 ( 
.A(n_918),
.B(n_913),
.C(n_867),
.Y(n_977)
);

AO21x1_ASAP7_75t_L g978 ( 
.A1(n_908),
.A2(n_954),
.B(n_953),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_917),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_936),
.B(n_940),
.Y(n_980)
);

NOR2xp67_ASAP7_75t_L g981 ( 
.A(n_931),
.B(n_949),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_930),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_852),
.B(n_941),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_880),
.B(n_954),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_881),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_855),
.A2(n_872),
.B(n_864),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_853),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_916),
.A2(n_929),
.B(n_933),
.C(n_922),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_856),
.A2(n_882),
.B(n_885),
.C(n_888),
.Y(n_989)
);

INVxp67_ASAP7_75t_SL g990 ( 
.A(n_935),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_866),
.A2(n_869),
.B(n_945),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_937),
.B(n_938),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_952),
.Y(n_993)
);

OAI21x1_ASAP7_75t_L g994 ( 
.A1(n_909),
.A2(n_956),
.B(n_868),
.Y(n_994)
);

AND2x6_ASAP7_75t_L g995 ( 
.A(n_906),
.B(n_932),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_946),
.A2(n_960),
.B1(n_854),
.B2(n_856),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_958),
.Y(n_997)
);

INVxp67_ASAP7_75t_L g998 ( 
.A(n_900),
.Y(n_998)
);

OAI21x1_ASAP7_75t_L g999 ( 
.A1(n_889),
.A2(n_879),
.B(n_935),
.Y(n_999)
);

INVx5_ASAP7_75t_L g1000 ( 
.A(n_906),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_962),
.B(n_950),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_SL g1002 ( 
.A1(n_879),
.A2(n_893),
.B(n_895),
.Y(n_1002)
);

OA21x2_ASAP7_75t_L g1003 ( 
.A1(n_892),
.A2(n_887),
.B(n_890),
.Y(n_1003)
);

OR2x6_ASAP7_75t_L g1004 ( 
.A(n_920),
.B(n_961),
.Y(n_1004)
);

OA21x2_ASAP7_75t_L g1005 ( 
.A1(n_891),
.A2(n_942),
.B(n_927),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_863),
.A2(n_901),
.B1(n_858),
.B2(n_896),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_857),
.B(n_948),
.Y(n_1007)
);

AO21x2_ASAP7_75t_L g1008 ( 
.A1(n_886),
.A2(n_942),
.B(n_927),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_924),
.A2(n_951),
.B(n_944),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_947),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_858),
.B(n_865),
.Y(n_1011)
);

CKINVDCx6p67_ASAP7_75t_R g1012 ( 
.A(n_884),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_870),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_878),
.A2(n_875),
.B1(n_876),
.B2(n_873),
.Y(n_1014)
);

AO31x2_ASAP7_75t_L g1015 ( 
.A1(n_860),
.A2(n_861),
.A3(n_897),
.B(n_934),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_850),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_943),
.B(n_915),
.Y(n_1017)
);

OR2x6_ASAP7_75t_L g1018 ( 
.A(n_946),
.B(n_779),
.Y(n_1018)
);

BUFx2_ASAP7_75t_L g1019 ( 
.A(n_919),
.Y(n_1019)
);

BUFx2_ASAP7_75t_R g1020 ( 
.A(n_867),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_883),
.Y(n_1021)
);

OA21x2_ASAP7_75t_L g1022 ( 
.A1(n_871),
.A2(n_851),
.B(n_955),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_855),
.A2(n_914),
.B(n_904),
.Y(n_1023)
);

NAND2x1p5_ASAP7_75t_L g1024 ( 
.A(n_919),
.B(n_859),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_SL g1025 ( 
.A1(n_874),
.A2(n_908),
.B(n_953),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_859),
.B(n_907),
.Y(n_1026)
);

OR2x2_ASAP7_75t_L g1027 ( 
.A(n_943),
.B(n_630),
.Y(n_1027)
);

BUFx2_ASAP7_75t_SL g1028 ( 
.A(n_959),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_899),
.B(n_939),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_855),
.A2(n_914),
.B(n_904),
.Y(n_1030)
);

NAND2x1p5_ASAP7_75t_L g1031 ( 
.A(n_919),
.B(n_859),
.Y(n_1031)
);

BUFx3_ASAP7_75t_L g1032 ( 
.A(n_964),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_964),
.Y(n_1033)
);

AO21x2_ASAP7_75t_L g1034 ( 
.A1(n_986),
.A2(n_991),
.B(n_1023),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_1001),
.A2(n_974),
.B1(n_978),
.B2(n_1025),
.Y(n_1035)
);

OR2x6_ASAP7_75t_L g1036 ( 
.A(n_996),
.B(n_1018),
.Y(n_1036)
);

AO21x2_ASAP7_75t_L g1037 ( 
.A1(n_986),
.A2(n_991),
.B(n_1023),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_966),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_966),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_984),
.B(n_975),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_985),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_971),
.Y(n_1042)
);

BUFx4f_ASAP7_75t_L g1043 ( 
.A(n_1018),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_999),
.B(n_1000),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1003),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_SL g1046 ( 
.A1(n_996),
.A2(n_982),
.B(n_973),
.C(n_998),
.Y(n_1046)
);

AO21x2_ASAP7_75t_L g1047 ( 
.A1(n_1030),
.A2(n_965),
.B(n_968),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_989),
.A2(n_988),
.B(n_965),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_1001),
.A2(n_974),
.B1(n_1006),
.B2(n_983),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_1022),
.Y(n_1050)
);

INVx5_ASAP7_75t_L g1051 ( 
.A(n_995),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_992),
.B(n_980),
.Y(n_1052)
);

OA21x2_ASAP7_75t_L g1053 ( 
.A1(n_994),
.A2(n_970),
.B(n_968),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_990),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_990),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_969),
.Y(n_1056)
);

INVxp67_ASAP7_75t_R g1057 ( 
.A(n_972),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_1026),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_967),
.B(n_1017),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_979),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1016),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_1050),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_1051),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1047),
.B(n_1005),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_1054),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_1044),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_1049),
.A2(n_1006),
.B1(n_974),
.B2(n_1002),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_1047),
.B(n_1005),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_SL g1069 ( 
.A1(n_1043),
.A2(n_974),
.B1(n_1011),
.B2(n_1036),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_1055),
.Y(n_1070)
);

OAI221xp5_ASAP7_75t_L g1071 ( 
.A1(n_1048),
.A2(n_973),
.B1(n_998),
.B2(n_983),
.C(n_1007),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_1047),
.B(n_1008),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_1047),
.B(n_1008),
.Y(n_1073)
);

NAND2x1_ASAP7_75t_L g1074 ( 
.A(n_1036),
.B(n_995),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_1042),
.B(n_1015),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1038),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_1036),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_1059),
.A2(n_1007),
.B1(n_1009),
.B2(n_1010),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_1053),
.B(n_1039),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1040),
.B(n_1029),
.Y(n_1080)
);

CKINVDCx14_ASAP7_75t_R g1081 ( 
.A(n_1052),
.Y(n_1081)
);

CKINVDCx14_ASAP7_75t_R g1082 ( 
.A(n_1052),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1045),
.B(n_1034),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_1083),
.B(n_1034),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1062),
.Y(n_1085)
);

INVxp67_ASAP7_75t_SL g1086 ( 
.A(n_1070),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_1083),
.B(n_1034),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1083),
.B(n_1034),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1072),
.B(n_1037),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1072),
.B(n_1037),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1080),
.B(n_1061),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1072),
.B(n_1037),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_1073),
.B(n_1037),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_1066),
.B(n_1036),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1076),
.Y(n_1095)
);

INVx2_ASAP7_75t_SL g1096 ( 
.A(n_1074),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_1081),
.B(n_963),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_1070),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1064),
.B(n_1068),
.Y(n_1099)
);

INVx5_ASAP7_75t_L g1100 ( 
.A(n_1063),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_1065),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_1086),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_1097),
.B(n_1081),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1099),
.B(n_1078),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1085),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1095),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1095),
.Y(n_1107)
);

OR2x2_ASAP7_75t_L g1108 ( 
.A(n_1099),
.B(n_1075),
.Y(n_1108)
);

OR2x2_ASAP7_75t_L g1109 ( 
.A(n_1099),
.B(n_1075),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1084),
.B(n_1068),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1084),
.B(n_1068),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1084),
.B(n_1079),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_1100),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1091),
.B(n_1078),
.Y(n_1114)
);

NOR2x1p5_ASAP7_75t_L g1115 ( 
.A(n_1086),
.B(n_1074),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1106),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_1103),
.Y(n_1117)
);

OR2x2_ASAP7_75t_L g1118 ( 
.A(n_1108),
.B(n_1087),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1105),
.Y(n_1119)
);

OR2x2_ASAP7_75t_L g1120 ( 
.A(n_1108),
.B(n_1087),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1107),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_1115),
.B(n_1096),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1112),
.B(n_1110),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1112),
.B(n_1087),
.Y(n_1124)
);

INVx1_ASAP7_75t_SL g1125 ( 
.A(n_1109),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_1102),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1104),
.B(n_1088),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1110),
.B(n_1088),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1116),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1127),
.B(n_1111),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1124),
.B(n_1111),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1125),
.B(n_1088),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1116),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_1126),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1121),
.Y(n_1135)
);

OAI31xp33_ASAP7_75t_L g1136 ( 
.A1(n_1122),
.A2(n_1082),
.A3(n_1071),
.B(n_1113),
.Y(n_1136)
);

OAI32xp33_ASAP7_75t_L g1137 ( 
.A1(n_1117),
.A2(n_1113),
.A3(n_1109),
.B1(n_1071),
.B2(n_987),
.Y(n_1137)
);

INVxp67_ASAP7_75t_L g1138 ( 
.A(n_1118),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1121),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_1122),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1124),
.B(n_1089),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1123),
.B(n_1089),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1119),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1119),
.Y(n_1144)
);

OAI32xp33_ASAP7_75t_L g1145 ( 
.A1(n_1118),
.A2(n_987),
.A3(n_1101),
.B1(n_1096),
.B2(n_1098),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_1122),
.B(n_1100),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1137),
.A2(n_1046),
.B(n_1082),
.C(n_1021),
.Y(n_1147)
);

AOI32xp33_ASAP7_75t_L g1148 ( 
.A1(n_1140),
.A2(n_1123),
.A3(n_1102),
.B1(n_1120),
.B2(n_1096),
.Y(n_1148)
);

AOI211xp5_ASAP7_75t_L g1149 ( 
.A1(n_1137),
.A2(n_1057),
.B(n_1114),
.C(n_981),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1146),
.A2(n_1057),
.B(n_1074),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1138),
.A2(n_1089),
.B1(n_1092),
.B2(n_1090),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1129),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1140),
.A2(n_1090),
.B1(n_1093),
.B2(n_1092),
.Y(n_1153)
);

INVxp67_ASAP7_75t_L g1154 ( 
.A(n_1134),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1129),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1141),
.A2(n_1090),
.B1(n_1093),
.B2(n_1092),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1154),
.A2(n_1136),
.B1(n_1094),
.B2(n_1077),
.Y(n_1157)
);

AOI21xp33_ASAP7_75t_SL g1158 ( 
.A1(n_1148),
.A2(n_1136),
.B(n_1145),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_1152),
.Y(n_1159)
);

OAI221xp5_ASAP7_75t_SL g1160 ( 
.A1(n_1149),
.A2(n_1067),
.B1(n_1035),
.B2(n_1120),
.C(n_1132),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1155),
.Y(n_1161)
);

NAND4xp75_ASAP7_75t_L g1162 ( 
.A(n_1150),
.B(n_1153),
.C(n_1151),
.D(n_1156),
.Y(n_1162)
);

NOR3xp33_ASAP7_75t_SL g1163 ( 
.A(n_1147),
.B(n_1013),
.C(n_1145),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1147),
.A2(n_1043),
.B(n_1143),
.Y(n_1164)
);

AOI221x1_ASAP7_75t_SL g1165 ( 
.A1(n_1149),
.A2(n_1142),
.B1(n_1130),
.B2(n_1128),
.C(n_1139),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1154),
.B(n_1028),
.Y(n_1166)
);

OAI222xp33_ASAP7_75t_L g1167 ( 
.A1(n_1148),
.A2(n_1131),
.B1(n_1141),
.B2(n_1069),
.C1(n_1077),
.C2(n_1139),
.Y(n_1167)
);

OAI221xp5_ASAP7_75t_SL g1168 ( 
.A1(n_1148),
.A2(n_1067),
.B1(n_1014),
.B2(n_1069),
.C(n_1012),
.Y(n_1168)
);

NAND2xp33_ASAP7_75t_SL g1169 ( 
.A(n_1163),
.B(n_963),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_1158),
.B(n_1100),
.Y(n_1170)
);

INVxp67_ASAP7_75t_L g1171 ( 
.A(n_1166),
.Y(n_1171)
);

AOI211x1_ASAP7_75t_L g1172 ( 
.A1(n_1167),
.A2(n_1131),
.B(n_1135),
.C(n_1133),
.Y(n_1172)
);

NAND4xp75_ASAP7_75t_L g1173 ( 
.A(n_1164),
.B(n_972),
.C(n_1020),
.D(n_1009),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_L g1174 ( 
.A(n_1160),
.B(n_1135),
.C(n_1133),
.Y(n_1174)
);

NAND4xp25_ASAP7_75t_SL g1175 ( 
.A(n_1157),
.B(n_1020),
.C(n_1014),
.D(n_977),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1161),
.Y(n_1176)
);

NAND3xp33_ASAP7_75t_L g1177 ( 
.A(n_1172),
.B(n_1168),
.C(n_1159),
.Y(n_1177)
);

NAND3xp33_ASAP7_75t_L g1178 ( 
.A(n_1170),
.B(n_1168),
.C(n_1159),
.Y(n_1178)
);

NAND4xp25_ASAP7_75t_L g1179 ( 
.A(n_1169),
.B(n_1165),
.C(n_1162),
.D(n_977),
.Y(n_1179)
);

NOR3xp33_ASAP7_75t_L g1180 ( 
.A(n_1175),
.B(n_976),
.C(n_1019),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1171),
.B(n_1143),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1176),
.B(n_1144),
.Y(n_1182)
);

AOI221x1_ASAP7_75t_L g1183 ( 
.A1(n_1174),
.A2(n_997),
.B1(n_993),
.B2(n_1060),
.C(n_1056),
.Y(n_1183)
);

NOR2x1_ASAP7_75t_L g1184 ( 
.A(n_1173),
.B(n_1004),
.Y(n_1184)
);

NAND2xp33_ASAP7_75t_L g1185 ( 
.A(n_1184),
.B(n_1024),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1181),
.Y(n_1186)
);

OR2x6_ASAP7_75t_L g1187 ( 
.A(n_1178),
.B(n_1024),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1182),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_R g1189 ( 
.A(n_1179),
.B(n_976),
.Y(n_1189)
);

NAND4xp25_ASAP7_75t_L g1190 ( 
.A(n_1177),
.B(n_1058),
.C(n_1032),
.D(n_1033),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_1183),
.Y(n_1191)
);

NOR2x1_ASAP7_75t_L g1192 ( 
.A(n_1187),
.B(n_1027),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1186),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1187),
.Y(n_1194)
);

NAND3xp33_ASAP7_75t_SL g1195 ( 
.A(n_1189),
.B(n_1180),
.C(n_1031),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1192),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1194),
.Y(n_1197)
);

XOR2xp5_ASAP7_75t_L g1198 ( 
.A(n_1197),
.B(n_1193),
.Y(n_1198)
);

NAND3xp33_ASAP7_75t_SL g1199 ( 
.A(n_1198),
.B(n_1197),
.C(n_1196),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_SL g1200 ( 
.A1(n_1199),
.A2(n_1195),
.B(n_1191),
.Y(n_1200)
);

OAI21xp33_ASAP7_75t_L g1201 ( 
.A1(n_1200),
.A2(n_1190),
.B(n_1188),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1201),
.B(n_1185),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1202),
.A2(n_1041),
.B1(n_1058),
.B2(n_1032),
.Y(n_1203)
);


endmodule