module fake_ibex_525_n_144 (n_7, n_20, n_17, n_25, n_36, n_18, n_3, n_22, n_28, n_32, n_4, n_33, n_5, n_11, n_30, n_6, n_29, n_13, n_2, n_8, n_26, n_35, n_14, n_0, n_9, n_34, n_12, n_15, n_37, n_24, n_31, n_10, n_23, n_21, n_27, n_19, n_16, n_1, n_144);

input n_7;
input n_20;
input n_17;
input n_25;
input n_36;
input n_18;
input n_3;
input n_22;
input n_28;
input n_32;
input n_4;
input n_33;
input n_5;
input n_11;
input n_30;
input n_6;
input n_29;
input n_13;
input n_2;
input n_8;
input n_26;
input n_35;
input n_14;
input n_0;
input n_9;
input n_34;
input n_12;
input n_15;
input n_37;
input n_24;
input n_31;
input n_10;
input n_23;
input n_21;
input n_27;
input n_19;
input n_16;
input n_1;

output n_144;

wire n_85;
wire n_128;
wire n_84;
wire n_64;
wire n_73;
wire n_65;
wire n_103;
wire n_95;
wire n_139;
wire n_55;
wire n_130;
wire n_63;
wire n_98;
wire n_129;
wire n_143;
wire n_106;
wire n_76;
wire n_118;
wire n_67;
wire n_38;
wire n_124;
wire n_110;
wire n_47;
wire n_108;
wire n_82;
wire n_78;
wire n_60;
wire n_86;
wire n_70;
wire n_87;
wire n_69;
wire n_75;
wire n_109;
wire n_127;
wire n_121;
wire n_137;
wire n_48;
wire n_57;
wire n_59;
wire n_125;
wire n_39;
wire n_62;
wire n_71;
wire n_120;
wire n_93;
wire n_122;
wire n_116;
wire n_61;
wire n_94;
wire n_134;
wire n_42;
wire n_77;
wire n_112;
wire n_88;
wire n_133;
wire n_44;
wire n_142;
wire n_51;
wire n_46;
wire n_80;
wire n_49;
wire n_66;
wire n_40;
wire n_74;
wire n_90;
wire n_58;
wire n_43;
wire n_140;
wire n_136;
wire n_119;
wire n_100;
wire n_72;
wire n_114;
wire n_97;
wire n_102;
wire n_131;
wire n_123;
wire n_52;
wire n_99;
wire n_135;
wire n_105;
wire n_126;
wire n_111;
wire n_104;
wire n_41;
wire n_45;
wire n_141;
wire n_89;
wire n_83;
wire n_53;
wire n_107;
wire n_115;
wire n_50;
wire n_92;
wire n_101;
wire n_113;
wire n_138;
wire n_96;
wire n_68;
wire n_117;
wire n_79;
wire n_81;
wire n_132;
wire n_56;
wire n_91;
wire n_54;

BUFx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx8_ASAP7_75t_SL g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

OAI21x1_ASAP7_75t_L g46 ( 
.A1(n_3),
.A2(n_7),
.B(n_6),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_23),
.B(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

OAI22x1_ASAP7_75t_SL g63 ( 
.A1(n_30),
.A2(n_27),
.B1(n_2),
.B2(n_12),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_5),
.B(n_9),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

AOI22x1_ASAP7_75t_SL g67 ( 
.A1(n_33),
.A2(n_2),
.B1(n_21),
.B2(n_11),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_15),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_44),
.B(n_51),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_53),
.B(n_49),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_70),
.B1(n_41),
.B2(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_71),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

NOR3xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_56),
.C(n_45),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_61),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

BUFx6f_ASAP7_75t_SL g83 ( 
.A(n_38),
.Y(n_83)
);

NOR3xp33_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_65),
.C(n_66),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_54),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

BUFx6f_ASAP7_75t_SL g87 ( 
.A(n_42),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_59),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_42),
.B(n_52),
.Y(n_91)
);

BUFx8_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

NAND2xp33_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_39),
.Y(n_93)
);

NOR3xp33_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_46),
.C(n_39),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_94),
.A2(n_70),
.B(n_85),
.C(n_81),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_95),
.B(n_89),
.C(n_82),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_83),
.Y(n_100)
);

NOR3xp33_ASAP7_75t_SL g101 ( 
.A(n_74),
.B(n_75),
.C(n_78),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_74),
.A2(n_87),
.B1(n_80),
.B2(n_88),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_93),
.B(n_91),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_95),
.B1(n_74),
.B2(n_77),
.Y(n_106)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_79),
.C(n_84),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_72),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_77),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_76),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_72),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_96),
.B(n_79),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_91),
.B(n_89),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_103),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_102),
.Y(n_115)
);

AOI222xp33_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_111),
.B1(n_109),
.B2(n_107),
.C1(n_97),
.C2(n_112),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_99),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_110),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_106),
.B1(n_105),
.B2(n_104),
.Y(n_121)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_123),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_98),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

INVx4_ASAP7_75t_R g128 ( 
.A(n_118),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_122),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_115),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_115),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_132),
.B1(n_117),
.B2(n_131),
.Y(n_137)
);

XOR2x1_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_125),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_117),
.B1(n_131),
.B2(n_133),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_139),
.A2(n_127),
.B1(n_129),
.B2(n_128),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_121),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_141),
.Y(n_144)
);


endmodule