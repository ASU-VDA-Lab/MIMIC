module fake_jpeg_14152_n_393 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_393);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_393;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_16),
.B(n_0),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_46),
.B(n_22),
.C(n_25),
.Y(n_105)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_R g48 ( 
.A(n_28),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_59),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx5_ASAP7_75t_SL g123 ( 
.A(n_50),
.Y(n_123)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_51),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_26),
.B(n_15),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_52),
.B(n_54),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_18),
.B(n_15),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_18),
.B(n_14),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_55),
.B(n_61),
.Y(n_102)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_69),
.Y(n_89)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_28),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_18),
.B(n_14),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_26),
.B(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_30),
.B(n_13),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_30),
.B(n_13),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_66),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_39),
.B(n_13),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_0),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_28),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_77),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_43),
.Y(n_71)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_24),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_80),
.Y(n_120)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_41),
.Y(n_94)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_43),
.B1(n_19),
.B2(n_21),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_84),
.A2(n_99),
.B1(n_111),
.B2(n_113),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_17),
.B1(n_40),
.B2(n_37),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_91),
.A2(n_58),
.B1(n_73),
.B2(n_79),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_46),
.A2(n_40),
.B1(n_37),
.B2(n_35),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_92),
.A2(n_108),
.B1(n_50),
.B2(n_74),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_46),
.A2(n_36),
.B1(n_22),
.B2(n_25),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_93),
.A2(n_109),
.B1(n_114),
.B2(n_118),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_105),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_71),
.A2(n_43),
.B1(n_21),
.B2(n_19),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_23),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_116),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_44),
.A2(n_35),
.B1(n_40),
.B2(n_37),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_44),
.A2(n_36),
.B1(n_23),
.B2(n_17),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_78),
.A2(n_21),
.B1(n_19),
.B2(n_17),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_78),
.A2(n_41),
.B1(n_29),
.B2(n_33),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_64),
.A2(n_41),
.B1(n_29),
.B2(n_33),
.Y(n_114)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx3_ASAP7_75t_SL g165 ( 
.A(n_115),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_54),
.B(n_33),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_53),
.A2(n_81),
.B1(n_76),
.B2(n_56),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_64),
.A2(n_41),
.B1(n_29),
.B2(n_33),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_124),
.A2(n_49),
.B1(n_74),
.B2(n_4),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_55),
.A2(n_12),
.B(n_18),
.C(n_3),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_127),
.B(n_48),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_61),
.B(n_1),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_2),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_63),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_129),
.B(n_141),
.Y(n_202)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_68),
.B1(n_80),
.B2(n_77),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_132),
.A2(n_142),
.B1(n_146),
.B2(n_154),
.Y(n_186)
);

OR2x2_ASAP7_75t_SL g133 ( 
.A(n_127),
.B(n_102),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_133),
.Y(n_191)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_135),
.Y(n_175)
);

BUFx24_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_136),
.Y(n_176)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_88),
.Y(n_138)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_138),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_100),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_151),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_L g141 ( 
.A1(n_98),
.A2(n_66),
.B(n_51),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_106),
.A2(n_45),
.B1(n_60),
.B2(n_76),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_143),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_101),
.B(n_70),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_145),
.B(n_153),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_81),
.B1(n_59),
.B2(n_97),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_150),
.Y(n_196)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_120),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_83),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_155),
.B(n_157),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_87),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_123),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_128),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_158),
.Y(n_199)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_117),
.A2(n_58),
.B1(n_75),
.B2(n_47),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_160),
.A2(n_121),
.B1(n_112),
.B2(n_108),
.Y(n_177)
);

AOI21xp33_ASAP7_75t_L g161 ( 
.A1(n_107),
.A2(n_48),
.B(n_58),
.Y(n_161)
);

MAJx2_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_166),
.C(n_92),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_105),
.B(n_72),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_162),
.Y(n_211)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_104),
.Y(n_163)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_164),
.A2(n_115),
.B1(n_110),
.B2(n_103),
.Y(n_193)
);

OR2x2_ASAP7_75t_SL g166 ( 
.A(n_89),
.B(n_67),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_171),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_94),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_89),
.B(n_12),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_169),
.A2(n_170),
.B1(n_110),
.B2(n_103),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_112),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_95),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_172),
.Y(n_198)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_119),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_82),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_155),
.A2(n_121),
.B1(n_112),
.B2(n_119),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_174),
.A2(n_193),
.B1(n_212),
.B2(n_171),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_177),
.A2(n_168),
.B1(n_172),
.B2(n_163),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_136),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_185),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_136),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_187),
.A2(n_74),
.B(n_3),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_137),
.B(n_95),
.C(n_125),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_197),
.C(n_208),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_137),
.B(n_126),
.C(n_82),
.Y(n_197)
);

INVxp67_ASAP7_75t_SL g219 ( 
.A(n_205),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_136),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_206),
.B(n_209),
.Y(n_217)
);

AND2x6_ASAP7_75t_L g207 ( 
.A(n_133),
.B(n_2),
.Y(n_207)
);

NOR2x1_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_143),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_137),
.B(n_126),
.C(n_96),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_150),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_159),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_213),
.B(n_157),
.Y(n_218)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_210),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_223),
.Y(n_255)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_218),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_220),
.A2(n_228),
.B1(n_232),
.B2(n_244),
.Y(n_252)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_221),
.Y(n_275)
);

OA22x2_ASAP7_75t_L g222 ( 
.A1(n_193),
.A2(n_154),
.B1(n_140),
.B2(n_164),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_222),
.B(n_230),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_210),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_184),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_234),
.Y(n_258)
);

BUFx5_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_225),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_178),
.A2(n_151),
.B1(n_147),
.B2(n_131),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_227),
.A2(n_239),
.B1(n_240),
.B2(n_205),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_211),
.A2(n_166),
.B1(n_131),
.B2(n_153),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_139),
.C(n_130),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_231),
.C(n_233),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_148),
.C(n_134),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_186),
.A2(n_169),
.B1(n_145),
.B2(n_165),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_167),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_184),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_135),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_237),
.Y(n_263)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_236),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_SL g238 ( 
.A1(n_187),
.A2(n_165),
.B(n_152),
.C(n_149),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_238),
.A2(n_243),
.B(n_244),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_212),
.A2(n_87),
.B1(n_165),
.B2(n_156),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_203),
.A2(n_156),
.B1(n_138),
.B2(n_96),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_188),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_241),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_199),
.B(n_173),
.Y(n_242)
);

A2O1A1O1Ixp25_ASAP7_75t_L g267 ( 
.A1(n_242),
.A2(n_204),
.B(n_195),
.C(n_201),
.D(n_176),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_243),
.B(n_6),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_191),
.A2(n_149),
.B1(n_3),
.B2(n_4),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_179),
.B(n_149),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_245),
.B(n_246),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_179),
.B(n_202),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_192),
.B(n_2),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_247),
.Y(n_262)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_188),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_248),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_216),
.A2(n_190),
.B1(n_192),
.B2(n_207),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_249),
.A2(n_253),
.B1(n_271),
.B2(n_240),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_250),
.A2(n_254),
.B(n_256),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_223),
.A2(n_177),
.B1(n_206),
.B2(n_185),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_226),
.A2(n_182),
.B(n_184),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_238),
.A2(n_176),
.B(n_200),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_268),
.Y(n_280)
);

MAJx2_ASAP7_75t_L g260 ( 
.A(n_215),
.B(n_204),
.C(n_195),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_229),
.C(n_231),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_227),
.A2(n_234),
.B(n_224),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_264),
.B(n_265),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_237),
.A2(n_235),
.B(n_217),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_267),
.B(n_221),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_239),
.A2(n_194),
.B1(n_201),
.B2(n_189),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_222),
.A2(n_189),
.B1(n_196),
.B2(n_175),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_10),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_232),
.A2(n_175),
.B1(n_196),
.B2(n_181),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_215),
.B(n_205),
.C(n_181),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_233),
.C(n_238),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_228),
.B(n_2),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_274),
.B(n_277),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_281),
.B(n_272),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_282),
.B(n_288),
.C(n_294),
.Y(n_307)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_275),
.Y(n_283)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_283),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_262),
.B(n_242),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_284),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_255),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_304),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_251),
.B(n_238),
.C(n_219),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_289),
.A2(n_290),
.B1(n_295),
.B2(n_296),
.Y(n_306)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_275),
.Y(n_291)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_291),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_261),
.Y(n_293)
);

INVx11_ASAP7_75t_L g324 ( 
.A(n_293),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_251),
.B(n_238),
.C(n_241),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_270),
.A2(n_222),
.B1(n_248),
.B2(n_214),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_270),
.A2(n_222),
.B1(n_236),
.B2(n_180),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_225),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_297),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_276),
.B(n_180),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_298),
.A2(n_300),
.B1(n_303),
.B2(n_278),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_260),
.B(n_6),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_274),
.C(n_254),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_273),
.B(n_7),
.Y(n_300)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_301),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_253),
.B(n_7),
.Y(n_302)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_302),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_270),
.A2(n_7),
.B1(n_9),
.B2(n_252),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_279),
.B(n_9),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_264),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_305),
.B(n_288),
.C(n_281),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_285),
.Y(n_311)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_311),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_312),
.B(n_277),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_314),
.B(n_317),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_315),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_283),
.B(n_279),
.Y(n_316)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_316),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_299),
.B(n_273),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_303),
.A2(n_263),
.B1(n_269),
.B2(n_256),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_322),
.Y(n_335)
);

FAx1_ASAP7_75t_SL g322 ( 
.A(n_294),
.B(n_258),
.CI(n_263),
.CON(n_322),
.SN(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_280),
.A2(n_265),
.B1(n_249),
.B2(n_250),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_323),
.A2(n_292),
.B1(n_295),
.B2(n_296),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_291),
.B(n_304),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_325),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_326),
.B(n_317),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_327),
.B(n_331),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_328),
.A2(n_306),
.B1(n_305),
.B2(n_319),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_320),
.B(n_293),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_329),
.B(n_339),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_314),
.B(n_286),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_330),
.B(n_307),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_307),
.B(n_258),
.C(n_286),
.Y(n_331)
);

BUFx12_ASAP7_75t_L g333 ( 
.A(n_324),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_333),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_316),
.B(n_302),
.Y(n_336)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_336),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_320),
.B(n_292),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_338),
.B(n_313),
.Y(n_350)
);

INVx2_ASAP7_75t_R g339 ( 
.A(n_322),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_323),
.A2(n_257),
.B(n_280),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_341),
.A2(n_289),
.B(n_308),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_308),
.B(n_275),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_343),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_344),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_347),
.B(n_357),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_348),
.B(n_355),
.Y(n_363)
);

AOI21x1_ASAP7_75t_L g366 ( 
.A1(n_349),
.A2(n_341),
.B(n_340),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_350),
.B(n_352),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_331),
.A2(n_310),
.B(n_322),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_330),
.B(n_310),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_337),
.A2(n_321),
.B1(n_319),
.B2(n_311),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_356),
.B(n_334),
.C(n_340),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_335),
.B(n_312),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_339),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_359),
.B(n_365),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_362),
.B(n_309),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_353),
.B(n_326),
.C(n_335),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_364),
.B(n_367),
.C(n_345),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_351),
.B(n_355),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_366),
.B(n_328),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_357),
.B(n_337),
.C(n_334),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_349),
.A2(n_347),
.B(n_345),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_368),
.A2(n_346),
.B1(n_354),
.B2(n_332),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_369),
.B(n_375),
.Y(n_384)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_370),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_371),
.B(n_376),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_374),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_363),
.B(n_348),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_361),
.B(n_346),
.C(n_342),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_359),
.B(n_342),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_360),
.B(n_309),
.C(n_343),
.Y(n_377)
);

INVxp33_ASAP7_75t_L g381 ( 
.A(n_377),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_377),
.A2(n_361),
.B1(n_358),
.B2(n_336),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_378),
.B(n_380),
.Y(n_385)
);

BUFx24_ASAP7_75t_SL g380 ( 
.A(n_373),
.Y(n_380)
);

OAI221xp5_ASAP7_75t_L g386 ( 
.A1(n_379),
.A2(n_339),
.B1(n_358),
.B2(n_325),
.C(n_360),
.Y(n_386)
);

AOI322xp5_ASAP7_75t_L g390 ( 
.A1(n_386),
.A2(n_387),
.A3(n_333),
.B1(n_259),
.B2(n_267),
.C1(n_266),
.C2(n_301),
.Y(n_390)
);

AOI322xp5_ASAP7_75t_L g387 ( 
.A1(n_384),
.A2(n_333),
.A3(n_324),
.B1(n_372),
.B2(n_259),
.C1(n_321),
.C2(n_376),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_383),
.B(n_374),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_388),
.B(n_381),
.C(n_382),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_389),
.A2(n_390),
.B(n_385),
.Y(n_391)
);

AOI321xp33_ASAP7_75t_L g392 ( 
.A1(n_391),
.A2(n_333),
.A3(n_266),
.B1(n_268),
.B2(n_287),
.C(n_9),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_392),
.B(n_287),
.Y(n_393)
);


endmodule