module real_jpeg_13716_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_336, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_336;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx10_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_3),
.A2(n_36),
.B1(n_61),
.B2(n_63),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_36),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_3),
.A2(n_36),
.B1(n_51),
.B2(n_56),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_4),
.A2(n_61),
.B1(n_63),
.B2(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_4),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_4),
.B(n_56),
.C(n_66),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_4),
.B(n_87),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_4),
.A2(n_122),
.B(n_175),
.Y(n_191)
);

O2A1O1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_4),
.A2(n_23),
.B(n_86),
.C(n_202),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_159),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_4),
.B(n_21),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_4),
.B(n_29),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_5),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_89),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_5),
.A2(n_61),
.B1(n_63),
.B2(n_89),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_5),
.A2(n_51),
.B1(n_56),
.B2(n_89),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_6),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_6),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_60),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_60),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_6),
.A2(n_51),
.B1(n_56),
.B2(n_60),
.Y(n_263)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_8),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_74),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_8),
.A2(n_51),
.B1(n_56),
.B2(n_74),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_8),
.A2(n_61),
.B1(n_63),
.B2(n_74),
.Y(n_252)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_10),
.A2(n_61),
.B1(n_63),
.B2(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_10),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_10),
.A2(n_51),
.B1(n_56),
.B2(n_171),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_171),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_171),
.Y(n_273)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_11),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_12),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_12),
.A2(n_51),
.B1(n_56),
.B2(n_131),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_12),
.A2(n_61),
.B1(n_63),
.B2(n_131),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_12),
.A2(n_23),
.B1(n_24),
.B2(n_131),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_13),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_13),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g259 ( 
.A(n_13),
.B(n_24),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_14),
.A2(n_32),
.B1(n_51),
.B2(n_56),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_14),
.A2(n_32),
.B1(n_61),
.B2(n_63),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_14),
.A2(n_23),
.B1(n_24),
.B2(n_32),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_15),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_15),
.A2(n_61),
.B1(n_63),
.B2(n_78),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_15),
.A2(n_51),
.B1(n_56),
.B2(n_78),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_15),
.A2(n_23),
.B1(n_24),
.B2(n_78),
.Y(n_209)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_39),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_37),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_33),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_26),
.B(n_31),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_21),
.A2(n_26),
.B1(n_31),
.B2(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_21),
.A2(n_26),
.B1(n_35),
.B2(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_22),
.A2(n_73),
.B(n_75),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_22),
.A2(n_27),
.B1(n_73),
.B2(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_22),
.B(n_77),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_22),
.A2(n_27),
.B1(n_98),
.B2(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_22),
.A2(n_75),
.B(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_22),
.A2(n_27),
.B1(n_130),
.B2(n_273),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_23),
.A2(n_24),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

AOI32xp33_ASAP7_75t_L g258 ( 
.A1(n_23),
.A2(n_25),
.A3(n_30),
.B1(n_246),
.B2(n_259),
.Y(n_258)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_26),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_27),
.A2(n_130),
.B(n_132),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_27),
.A2(n_30),
.B(n_159),
.C(n_245),
.Y(n_244)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_33),
.B(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_34),
.B(n_331),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_330),
.B(n_332),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_318),
.B(n_329),
.Y(n_40)
);

AO21x1_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_147),
.B(n_315),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_134),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_109),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_44),
.B(n_109),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_79),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_45),
.B(n_80),
.C(n_95),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B(n_72),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_46),
.A2(n_47),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_57),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_48),
.A2(n_49),
.B1(n_72),
.B2(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_48),
.A2(n_49),
.B1(n_57),
.B2(n_58),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_53),
.B(n_54),
.Y(n_49)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_50),
.A2(n_53),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_50),
.B(n_176),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_50),
.A2(n_53),
.B1(n_121),
.B2(n_263),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

INVx5_ASAP7_75t_SL g56 ( 
.A(n_51),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_56),
.B1(n_66),
.B2(n_67),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_51),
.B(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_53),
.B(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_55),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_64),
.B1(n_69),
.B2(n_71),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_59),
.A2(n_64),
.B1(n_71),
.B2(n_126),
.Y(n_125)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

AO22x1_ASAP7_75t_SL g87 ( 
.A1(n_61),
.A2(n_63),
.B1(n_85),
.B2(n_86),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_61),
.B(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g202 ( 
.A1(n_63),
.A2(n_85),
.B(n_159),
.Y(n_202)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_64),
.A2(n_71),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_64),
.B(n_161),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_64),
.A2(n_71),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_64),
.A2(n_71),
.B1(n_126),
.B2(n_252),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_70),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_68),
.A2(n_170),
.B(n_172),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_68),
.B(n_159),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_68),
.A2(n_172),
.B(n_251),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_71),
.B(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_95),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_80),
.A2(n_81),
.B(n_92),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_92),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_82),
.A2(n_88),
.B1(n_90),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_82),
.A2(n_90),
.B1(n_103),
.B2(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_82),
.A2(n_207),
.B(n_208),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_82),
.A2(n_90),
.B1(n_222),
.B2(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_82),
.A2(n_208),
.B(n_249),
.Y(n_271)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_87),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_83),
.B(n_209),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_83),
.A2(n_87),
.B(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_87),
.B(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_90),
.A2(n_222),
.B(n_223),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_90),
.A2(n_128),
.B(n_223),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_SL g157 ( 
.A1(n_93),
.A2(n_158),
.B(n_160),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_93),
.A2(n_160),
.B(n_234),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_99),
.B2(n_108),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_96),
.A2(n_97),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_SL g145 ( 
.A(n_97),
.B(n_100),
.C(n_105),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_97),
.B(n_138),
.C(n_145),
.Y(n_328)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_100),
.Y(n_107)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_104),
.A2(n_105),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_105),
.B(n_139),
.C(n_143),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_115),
.C(n_116),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_110),
.A2(n_111),
.B1(n_115),
.B2(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_115),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_116),
.B(n_312),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_127),
.C(n_129),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_117),
.A2(n_118),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_124),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_119),
.A2(n_124),
.B1(n_125),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_119),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_122),
.A2(n_174),
.B(n_175),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_122),
.A2(n_123),
.B1(n_204),
.B2(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_122),
.A2(n_123),
.B1(n_229),
.B2(n_262),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_123),
.A2(n_181),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_123),
.B(n_159),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_123),
.A2(n_189),
.B(n_204),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_127),
.B(n_129),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_133),
.B(n_244),
.Y(n_243)
);

OAI21xp33_ASAP7_75t_L g315 ( 
.A1(n_134),
.A2(n_316),
.B(n_317),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_146),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_135),
.B(n_146),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_145),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_140),
.Y(n_324)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_144),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_309),
.B(n_314),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_297),
.B(n_308),
.Y(n_148)
);

OAI321xp33_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_265),
.A3(n_290),
.B1(n_295),
.B2(n_296),
.C(n_336),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_238),
.B(n_264),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_216),
.B(n_237),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_197),
.B(n_215),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_177),
.B(n_196),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_164),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_155),
.B(n_164),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_162),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_156),
.A2(n_157),
.B1(n_162),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_173),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_169),
.C(n_173),
.Y(n_198)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_174),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_185),
.B(n_195),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_179),
.B(n_183),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_190),
.B(n_194),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_187),
.B(n_188),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_198),
.B(n_199),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_205),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_210),
.C(n_214),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_203),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_203),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_210),
.B1(n_213),
.B2(n_214),
.Y(n_205)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_206),
.Y(n_214)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_210),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_217),
.B(n_218),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_230),
.B2(n_231),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_233),
.C(n_235),
.Y(n_239)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_221),
.B(n_225),
.C(n_228),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_235),
.B2(n_236),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_232),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_233),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_239),
.B(n_240),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_254),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_241),
.B(n_255),
.C(n_256),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_247),
.B2(n_253),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_242),
.B(n_248),
.C(n_250),
.Y(n_279)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_247),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_250),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_260),
.B2(n_261),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_261),
.Y(n_275)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_280),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_266),
.B(n_280),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_276),
.C(n_279),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_267),
.A2(n_268),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_275),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_274),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_274),
.C(n_275),
.Y(n_289)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_272),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_276),
.B(n_279),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_278),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_289),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_282),
.B(n_284),
.C(n_289),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_288),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_287),
.C(n_288),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_291),
.B(n_292),
.Y(n_295)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_307),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_307),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_302),
.C(n_303),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_311),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_328),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_328),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_327),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_323),
.B1(n_325),
.B2(n_326),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_321),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_323),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_325),
.C(n_327),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_331),
.Y(n_334)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);


endmodule