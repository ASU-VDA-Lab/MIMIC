module fake_jpeg_11558_n_234 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_234);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_234;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NAND2x1_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_0),
.Y(n_40)
);

AND2x4_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_34),
.Y(n_68)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_12),
.Y(n_45)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_50),
.Y(n_79)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_22),
.B(n_11),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_56),
.Y(n_86)
);

HAxp5_ASAP7_75t_SL g52 ( 
.A(n_19),
.B(n_0),
.CON(n_52),
.SN(n_52)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_57),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_26),
.B(n_31),
.Y(n_54)
);

NAND3xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_31),
.C(n_27),
.Y(n_81)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_59),
.Y(n_89)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_36),
.Y(n_92)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_62),
.Y(n_91)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_60),
.B(n_35),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_64),
.B(n_82),
.Y(n_113)
);

NOR2xp67_ASAP7_75t_SL g119 ( 
.A(n_68),
.B(n_10),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_34),
.B1(n_38),
.B2(n_21),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_69),
.A2(n_72),
.B1(n_83),
.B2(n_53),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_28),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_73),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_21),
.B1(n_38),
.B2(n_18),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_20),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_20),
.Y(n_74)
);

MAJx2_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_75),
.C(n_80),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_28),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_24),
.B1(n_33),
.B2(n_17),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_77),
.A2(n_85),
.B1(n_23),
.B2(n_46),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_27),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_36),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_17),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_53),
.A2(n_18),
.B1(n_36),
.B2(n_25),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_33),
.B1(n_24),
.B2(n_25),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_42),
.B(n_37),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_87),
.B(n_2),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_92),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_41),
.B1(n_58),
.B2(n_25),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_94),
.A2(n_95),
.B1(n_121),
.B2(n_78),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_68),
.A2(n_37),
.B1(n_35),
.B2(n_23),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_90),
.Y(n_96)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_97),
.A2(n_122),
.B1(n_93),
.B2(n_65),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_98),
.B(n_114),
.Y(n_147)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_71),
.Y(n_140)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_66),
.A2(n_43),
.B(n_50),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_108),
.A2(n_119),
.B(n_10),
.Y(n_142)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_89),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_112),
.Y(n_129)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_66),
.A2(n_50),
.B(n_3),
.C(n_4),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_116),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_67),
.B(n_2),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_120),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_68),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_118),
.A2(n_88),
.B1(n_84),
.B2(n_64),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_73),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_75),
.A2(n_74),
.B1(n_70),
.B2(n_82),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_5),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_122),
.B(n_86),
.Y(n_127)
);

A2O1A1O1Ixp25_ASAP7_75t_L g165 ( 
.A1(n_127),
.A2(n_113),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_133),
.Y(n_152)
);

O2A1O1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_78),
.B(n_84),
.C(n_87),
.Y(n_130)
);

AO22x1_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_120),
.B1(n_103),
.B2(n_110),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_136),
.B1(n_96),
.B2(n_101),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_100),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_98),
.A2(n_93),
.B1(n_71),
.B2(n_8),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_102),
.B(n_93),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_144),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_94),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_95),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_105),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_106),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_109),
.C(n_102),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_160),
.C(n_162),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_142),
.A2(n_119),
.B(n_115),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_157),
.B(n_140),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_165),
.C(n_141),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_154),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_111),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_155),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_156),
.Y(n_178)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_109),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_123),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_112),
.C(n_107),
.Y(n_162)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_113),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_164),
.B(n_146),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_166),
.A2(n_136),
.B1(n_132),
.B2(n_145),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_132),
.A2(n_96),
.B1(n_99),
.B2(n_5),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_7),
.C(n_131),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_124),
.C(n_133),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_161),
.A2(n_130),
.B(n_141),
.Y(n_169)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_169),
.A2(n_171),
.B(n_172),
.Y(n_190)
);

AOI221xp5_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_147),
.B1(n_128),
.B2(n_138),
.C(n_144),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_126),
.C(n_145),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_148),
.C(n_149),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_175),
.B(n_181),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_156),
.B(n_143),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_166),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_161),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_162),
.Y(n_196)
);

NAND3xp33_ASAP7_75t_SL g186 ( 
.A(n_180),
.B(n_152),
.C(n_150),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_187),
.Y(n_203)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_189),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_173),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_178),
.A2(n_153),
.B1(n_156),
.B2(n_154),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_192),
.A2(n_199),
.B(n_182),
.Y(n_202)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_193),
.B(n_195),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_176),
.A2(n_153),
.B1(n_168),
.B2(n_140),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_194),
.A2(n_182),
.B1(n_178),
.B2(n_169),
.Y(n_205)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_197),
.C(n_198),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_157),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_198),
.C(n_170),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_207),
.C(n_208),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_209),
.Y(n_210)
);

AO21x1_ASAP7_75t_L g212 ( 
.A1(n_205),
.A2(n_192),
.B(n_199),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_174),
.C(n_183),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_175),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_191),
.B1(n_187),
.B2(n_195),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_206),
.B(n_190),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_211),
.B(n_214),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_212),
.A2(n_215),
.B(n_177),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_204),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_188),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_193),
.C(n_165),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_137),
.Y(n_221)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_135),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_219),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_210),
.A2(n_200),
.B1(n_201),
.B2(n_184),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_135),
.C(n_137),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_221),
.Y(n_226)
);

OAI221xp5_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_184),
.B1(n_210),
.B2(n_215),
.C(n_219),
.Y(n_225)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_225),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_222),
.B(n_220),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_226),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_228),
.Y(n_231)
);

INVxp33_ASAP7_75t_L g229 ( 
.A(n_224),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_229),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_232),
.A2(n_230),
.B(n_231),
.Y(n_233)
);

BUFx24_ASAP7_75t_SL g234 ( 
.A(n_233),
.Y(n_234)
);


endmodule