module fake_jpeg_18078_n_255 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_255);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_255;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_7),
.B(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_41),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_0),
.C(n_1),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_26),
.B1(n_18),
.B2(n_25),
.Y(n_57)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_43),
.Y(n_53)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_44),
.B(n_58),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_31),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_36),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_34),
.B1(n_27),
.B2(n_19),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_30),
.B1(n_29),
.B2(n_33),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_27),
.B1(n_19),
.B2(n_34),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_50),
.A2(n_55),
.B1(n_17),
.B2(n_25),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_27),
.B1(n_19),
.B2(n_26),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_32),
.C(n_29),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_28),
.Y(n_61)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_68),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_65),
.A2(n_76),
.B1(n_81),
.B2(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_73),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_17),
.B1(n_18),
.B2(n_33),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_79),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_31),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_20),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_39),
.C(n_36),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_82),
.Y(n_109)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_46),
.A2(n_30),
.B1(n_32),
.B2(n_22),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_39),
.C(n_35),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_32),
.Y(n_84)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_86),
.Y(n_113)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_56),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_88),
.A2(n_46),
.B1(n_49),
.B2(n_47),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_32),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_89),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_53),
.A2(n_22),
.B1(n_24),
.B2(n_20),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_115),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_64),
.A2(n_58),
.B(n_53),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_95),
.A2(n_96),
.B(n_20),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_48),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_112),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_105),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_77),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_110),
.A2(n_82),
.B1(n_71),
.B2(n_75),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_47),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_55),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_20),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_20),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_112),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g118 ( 
.A1(n_70),
.A2(n_49),
.B1(n_46),
.B2(n_60),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_49),
.B1(n_72),
.B2(n_80),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_123),
.B1(n_134),
.B2(n_96),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_121),
.A2(n_133),
.B1(n_93),
.B2(n_127),
.Y(n_161)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_103),
.A2(n_98),
.B1(n_108),
.B2(n_99),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_76),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_125),
.C(n_129),
.Y(n_169)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_72),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_116),
.Y(n_130)
);

XNOR2x1_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_141),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_133),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_74),
.B1(n_69),
.B2(n_83),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_137),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_79),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_101),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_88),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_138),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_85),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_139),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_140),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_96),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_102),
.A2(n_99),
.B(n_111),
.C(n_117),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_143),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_104),
.B(n_74),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_106),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_144),
.A2(n_100),
.B1(n_93),
.B2(n_4),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_104),
.B(n_21),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_100),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_111),
.B(n_110),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_146),
.A2(n_131),
.B(n_141),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_151),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_163),
.Y(n_174)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_119),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_159),
.B(n_160),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_135),
.Y(n_162)
);

BUFx24_ASAP7_75t_SL g172 ( 
.A(n_162),
.Y(n_172)
);

AO22x2_ASAP7_75t_L g163 ( 
.A1(n_123),
.A2(n_24),
.B1(n_21),
.B2(n_5),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_144),
.A2(n_21),
.B1(n_3),
.B2(n_6),
.Y(n_165)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_0),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_168),
.Y(n_178)
);

NOR2x1_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_7),
.Y(n_167)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

OA22x2_ASAP7_75t_L g168 ( 
.A1(n_120),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_121),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_170)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_147),
.Y(n_173)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_130),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_181),
.C(n_148),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_176),
.A2(n_150),
.B(n_160),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_129),
.B(n_125),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_180),
.A2(n_192),
.B(n_168),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_122),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_11),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_151),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_187),
.A2(n_167),
.B1(n_154),
.B2(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_156),
.Y(n_191)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

NAND3xp33_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_14),
.C(n_15),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_193),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_206),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_195),
.A2(n_204),
.B1(n_208),
.B2(n_183),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_201),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_174),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_209),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_150),
.C(n_146),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_205),
.C(n_178),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_179),
.A2(n_163),
.B1(n_155),
.B2(n_158),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_157),
.C(n_158),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_176),
.A2(n_171),
.B(n_152),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_168),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g210 ( 
.A(n_207),
.B(n_174),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_179),
.A2(n_168),
.B1(n_163),
.B2(n_171),
.Y(n_208)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_216),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_204),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_214),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_172),
.C(n_180),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_195),
.A2(n_188),
.B1(n_178),
.B2(n_191),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_185),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_218),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_182),
.C(n_187),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_196),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_163),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_208),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_232),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_227),
.B(n_215),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_200),
.Y(n_228)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_202),
.C(n_207),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_230),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_221),
.A2(n_193),
.B(n_207),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_186),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_225),
.A2(n_213),
.B(n_215),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_233),
.A2(n_240),
.B(n_210),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_229),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_234),
.A2(n_232),
.B(n_184),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_223),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_198),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_224),
.Y(n_243)
);

AO22x1_ASAP7_75t_L g240 ( 
.A1(n_231),
.A2(n_210),
.B1(n_222),
.B2(n_163),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_242),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_223),
.C(n_217),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_243),
.B(n_244),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_238),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_247),
.B(n_248),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_239),
.B1(n_234),
.B2(n_240),
.Y(n_248)
);

A2O1A1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_249),
.A2(n_246),
.B(n_149),
.C(n_15),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_251),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_249),
.A2(n_16),
.B(n_11),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_253),
.B(n_250),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_252),
.Y(n_255)
);


endmodule