module real_jpeg_6921_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_1),
.A2(n_47),
.B1(n_89),
.B2(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_2),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_3),
.A2(n_146),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_3),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_3),
.A2(n_63),
.B1(n_185),
.B2(n_327),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_3),
.A2(n_185),
.B1(n_312),
.B2(n_347),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g415 ( 
.A1(n_3),
.A2(n_185),
.B1(n_416),
.B2(n_418),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_4),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_4),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_4),
.A2(n_116),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_L g229 ( 
.A1(n_4),
.A2(n_116),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g386 ( 
.A1(n_4),
.A2(n_116),
.B1(n_320),
.B2(n_387),
.Y(n_386)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_5),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_6),
.Y(n_181)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_6),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_6),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_6),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_7),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_7),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_7),
.A2(n_148),
.B1(n_197),
.B2(n_276),
.Y(n_275)
);

OAI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_7),
.A2(n_148),
.B1(n_309),
.B2(n_311),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_7),
.A2(n_148),
.B1(n_300),
.B2(n_373),
.Y(n_372)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_8),
.Y(n_130)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_8),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_8),
.Y(n_137)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_8),
.Y(n_144)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_9),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_10),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_10),
.A2(n_262),
.B1(n_289),
.B2(n_291),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_10),
.B(n_302),
.C(n_304),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_10),
.B(n_108),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_10),
.B(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_10),
.B(n_92),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_10),
.B(n_114),
.Y(n_382)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_11),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_11),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_11),
.Y(n_147)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_11),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_11),
.Y(n_188)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_11),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_11),
.Y(n_233)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_12),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_12),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_13),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_13),
.A2(n_36),
.B1(n_55),
.B2(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_14),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_14),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_14),
.A2(n_38),
.B1(n_49),
.B2(n_88),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_14),
.A2(n_88),
.B1(n_209),
.B2(n_211),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_15),
.A2(n_55),
.B1(n_60),
.B2(n_61),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_15),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_15),
.A2(n_60),
.B1(n_121),
.B2(n_123),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_15),
.A2(n_49),
.B1(n_52),
.B2(n_60),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_16),
.A2(n_152),
.B1(n_153),
.B2(n_155),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_16),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_16),
.A2(n_152),
.B1(n_194),
.B2(n_196),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_16),
.A2(n_56),
.B1(n_76),
.B2(n_152),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_16),
.A2(n_152),
.B1(n_319),
.B2(n_321),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_236),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_235),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_200),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_20),
.B(n_200),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_157),
.C(n_166),
.Y(n_20)
);

FAx1_ASAP7_75t_SL g278 ( 
.A(n_21),
.B(n_157),
.CI(n_166),
.CON(n_278),
.SN(n_278)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_93),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_22),
.B(n_94),
.C(n_124),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_53),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_23),
.B(n_53),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_33),
.B1(n_41),
.B2(n_46),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_24),
.A2(n_43),
.B(n_46),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_24),
.A2(n_268),
.B1(n_270),
.B2(n_272),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_24),
.A2(n_308),
.B(n_315),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_24),
.A2(n_262),
.B(n_315),
.Y(n_343)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_25),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_25),
.B(n_318),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_25),
.A2(n_358),
.B1(n_359),
.B2(n_360),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_25),
.A2(n_42),
.B1(n_269),
.B2(n_386),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_30),
.Y(n_320)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_31),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_31),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_33),
.Y(n_179)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_35),
.Y(n_305)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_38),
.Y(n_310)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_40),
.Y(n_388)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_45),
.Y(n_342)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_45),
.Y(n_361)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g322 ( 
.A(n_50),
.Y(n_322)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_64),
.B1(n_87),
.B2(n_92),
.Y(n_53)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_54),
.Y(n_176)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AO22x2_ASAP7_75t_L g108 ( 
.A1(n_57),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_58),
.Y(n_163)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_58),
.Y(n_294)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_59),
.Y(n_220)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_59),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_59),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_64),
.A2(n_87),
.B1(n_92),
.B2(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_64),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_64),
.A2(n_92),
.B1(n_160),
.B2(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_64),
.B(n_296),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_79),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_69),
.B1(n_72),
.B2(n_76),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_73),
.A2(n_80),
.B1(n_82),
.B2(n_84),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_78),
.Y(n_174)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_79),
.A2(n_326),
.B(n_330),
.Y(n_325)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_86),
.Y(n_303)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_91),
.Y(n_290)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_92),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_92),
.B(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_124),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_113),
.B1(n_119),
.B2(n_120),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_95),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_95),
.A2(n_119),
.B1(n_275),
.B2(n_415),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_108),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_102),
.B1(n_103),
.B2(n_107),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_101),
.Y(n_397)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_101),
.Y(n_404)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g276 ( 
.A(n_105),
.Y(n_276)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_106),
.Y(n_195)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_106),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_106),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_106),
.Y(n_380)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_106),
.Y(n_420)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

AOI22x1_ASAP7_75t_L g190 ( 
.A1(n_108),
.A2(n_191),
.B1(n_192),
.B2(n_199),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_108),
.A2(n_191),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_113),
.Y(n_199)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_118),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_119),
.B(n_193),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_119),
.A2(n_415),
.B(n_421),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_120),
.Y(n_207)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_145),
.B(n_150),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_125),
.A2(n_145),
.B1(n_184),
.B2(n_189),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_126),
.B(n_151),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_126),
.A2(n_439),
.B(n_440),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_134),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_SL g255 ( 
.A(n_130),
.Y(n_255)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_138),
.B1(n_141),
.B2(n_143),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_137),
.Y(n_257)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_140),
.Y(n_212)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_149),
.Y(n_155)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_150),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_156),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_SL g439 ( 
.A1(n_153),
.A2(n_261),
.B(n_262),
.Y(n_439)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_156),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_156),
.B(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_164),
.B2(n_165),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_159),
.B(n_164),
.Y(n_224)
);

INVx3_ASAP7_75t_SL g161 ( 
.A(n_162),
.Y(n_161)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_164),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_164),
.A2(n_165),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_182),
.C(n_190),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_167),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_177),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_168),
.B(n_177),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_175),
.B2(n_176),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_169),
.A2(n_288),
.B(n_295),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_169),
.A2(n_175),
.B1(n_326),
.B2(n_372),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_169),
.A2(n_295),
.B(n_372),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_170),
.A2(n_175),
.B(n_330),
.Y(n_443)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_178),
.Y(n_272)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_182),
.A2(n_183),
.B1(n_190),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_184),
.A2(n_189),
.B(n_234),
.Y(n_247)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_189),
.B(n_262),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_190),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_191),
.A2(n_274),
.B(n_277),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_191),
.A2(n_277),
.B(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_191),
.B(n_192),
.Y(n_421)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_198),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_222),
.B2(n_223),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_213),
.B(n_221),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_214),
.Y(n_221)
);

INVx6_ASAP7_75t_SL g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_219),
.Y(n_300)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_234),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_279),
.B(n_468),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_278),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_239),
.B(n_278),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_244),
.C(n_245),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_240),
.A2(n_241),
.B1(n_244),
.B2(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_244),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_245),
.B(n_458),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.C(n_273),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_246),
.A2(n_247),
.B1(n_273),
.B2(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_248),
.B(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_266),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_249),
.A2(n_266),
.B1(n_267),
.B2(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_249),
.Y(n_432)
);

OAI32xp33_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_252),
.A3(n_254),
.B1(n_256),
.B2(n_261),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

OAI21xp33_ASAP7_75t_SL g376 ( 
.A1(n_262),
.A2(n_377),
.B(n_381),
.Y(n_376)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_273),
.Y(n_453)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

AOI32xp33_ASAP7_75t_L g391 ( 
.A1(n_276),
.A2(n_382),
.A3(n_392),
.B1(n_394),
.B2(n_398),
.Y(n_391)
);

BUFx24_ASAP7_75t_SL g471 ( 
.A(n_278),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_446),
.B(n_465),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

AOI21x1_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_427),
.B(n_445),
.Y(n_281)
);

AO21x1_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_406),
.B(n_426),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_366),
.B(n_405),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_333),
.B(n_365),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_306),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_286),
.B(n_306),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_297),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_287),
.A2(n_297),
.B1(n_298),
.B2(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_287),
.Y(n_363)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx6_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_294),
.Y(n_393)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_294),
.Y(n_401)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_323),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_307),
.B(n_324),
.C(n_332),
.Y(n_367)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_308),
.Y(n_359)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx4_ASAP7_75t_SL g312 ( 
.A(n_313),
.Y(n_312)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_318),
.Y(n_315)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_324),
.A2(n_325),
.B1(n_331),
.B2(n_332),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_356),
.B(n_364),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_344),
.B(n_355),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_343),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_341),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_338),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

BUFx5_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_354),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_345),
.B(n_354),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_350),
.B(n_353),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_346),
.Y(n_358)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx6_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx3_ASAP7_75t_SL g350 ( 
.A(n_351),
.Y(n_350)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_352),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_353),
.A2(n_385),
.B(n_389),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_362),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_357),
.B(n_362),
.Y(n_364)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_367),
.B(n_368),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_383),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_370),
.A2(n_371),
.B1(n_374),
.B2(n_375),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_371),
.B(n_374),
.C(n_383),
.Y(n_407)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_380),
.Y(n_417)
);

INVxp33_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_391),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_384),
.B(n_391),
.Y(n_412)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

NAND2xp33_ASAP7_75t_SL g398 ( 
.A(n_399),
.B(n_402),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_407),
.B(n_408),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_409),
.A2(n_410),
.B1(n_413),
.B2(n_425),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_412),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_411),
.B(n_412),
.C(n_425),
.Y(n_428)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_413),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_414),
.B(n_422),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_414),
.B(n_423),
.C(n_424),
.Y(n_433)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_429),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_428),
.B(n_429),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_436),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_431),
.A2(n_433),
.B1(n_434),
.B2(n_435),
.Y(n_430)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_431),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_433),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_433),
.B(n_434),
.C(n_436),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_437),
.A2(n_438),
.B1(n_441),
.B2(n_444),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_437),
.B(n_442),
.C(n_443),
.Y(n_456)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_441),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_442),
.B(n_443),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_448),
.B(n_460),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_449),
.A2(n_466),
.B(n_467),
.Y(n_465)
);

NOR2x1_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_457),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_450),
.B(n_457),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_454),
.C(n_456),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_451),
.B(n_463),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_454),
.A2(n_455),
.B1(n_456),
.B2(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_456),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_462),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_461),
.B(n_462),
.Y(n_466)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);


endmodule