module fake_jpeg_29628_n_154 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_154);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_154;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_34),
.B(n_47),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_12),
.B(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_12),
.B(n_11),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_40),
.Y(n_60)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_0),
.C(n_1),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_0),
.B(n_2),
.Y(n_52)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_46),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_16),
.B(n_11),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

AO22x2_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_18),
.B1(n_21),
.B2(n_19),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_59),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_30),
.A2(n_21),
.B1(n_22),
.B2(n_19),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_26),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_67),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_21),
.B1(n_22),
.B2(n_26),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_14),
.B1(n_23),
.B2(n_20),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_31),
.A2(n_13),
.B1(n_23),
.B2(n_20),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_35),
.A2(n_17),
.B1(n_14),
.B2(n_24),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_61),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_43),
.B1(n_17),
.B2(n_44),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_67),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_47),
.A2(n_24),
.B1(n_13),
.B2(n_7),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_65),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_25),
.B1(n_6),
.B2(n_4),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_33),
.B(n_9),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_45),
.A2(n_25),
.B1(n_4),
.B2(n_10),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_71),
.Y(n_77)
);

OR2x4_ASAP7_75t_L g71 ( 
.A(n_33),
.B(n_25),
.Y(n_71)
);

AND2x4_ASAP7_75t_L g73 ( 
.A(n_33),
.B(n_25),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_51),
.B(n_4),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_79),
.B(n_82),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_86),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_66),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_95),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_63),
.B1(n_48),
.B2(n_71),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_108),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_76),
.A2(n_89),
.B(n_88),
.C(n_94),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_99),
.B(n_94),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_73),
.B(n_74),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_80),
.B(n_52),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_102),
.B(n_109),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_78),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_84),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_64),
.B1(n_70),
.B2(n_73),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_95),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_93),
.C(n_89),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_117),
.Y(n_127)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

AO221x1_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_114),
.B1(n_118),
.B2(n_119),
.C(n_120),
.Y(n_125)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_123),
.B(n_98),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_76),
.C(n_77),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_80),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_77),
.Y(n_123)
);

AOI221xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_99),
.B1(n_110),
.B2(n_97),
.C(n_98),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_126),
.B(n_132),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_98),
.B(n_108),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_130),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_121),
.A2(n_90),
.B1(n_85),
.B2(n_75),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_131),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_90),
.B1(n_114),
.B2(n_117),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_124),
.A2(n_112),
.B1(n_111),
.B2(n_107),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_134),
.A2(n_92),
.B1(n_70),
.B2(n_111),
.Y(n_144)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_101),
.Y(n_140)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_138),
.B(n_139),
.Y(n_141)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_140),
.B(n_142),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_127),
.C(n_107),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_134),
.B(n_103),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_144),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_127),
.C(n_135),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_147),
.A2(n_148),
.B1(n_136),
.B2(n_144),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_135),
.C(n_137),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_150),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_145),
.A2(n_91),
.B1(n_105),
.B2(n_87),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_149),
.A2(n_146),
.B(n_83),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_151),
.A2(n_54),
.B1(n_56),
.B2(n_72),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_152),
.Y(n_154)
);


endmodule