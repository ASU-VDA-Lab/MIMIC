module fake_jpeg_19068_n_254 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_254);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_155;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_100;
wire n_96;

INVx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_25),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_37),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx5_ASAP7_75t_SL g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_1),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_18),
.Y(n_54)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_27),
.B1(n_17),
.B2(n_28),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_49),
.B1(n_53),
.B2(n_56),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_24),
.B(n_23),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_27),
.B1(n_17),
.B2(n_16),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_39),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_36),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_33),
.A2(n_27),
.B1(n_17),
.B2(n_28),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_54),
.B(n_35),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_33),
.A2(n_16),
.B1(n_28),
.B2(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_61),
.Y(n_98)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_63),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_64),
.B(n_71),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_33),
.B1(n_37),
.B2(n_24),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_67),
.A2(n_29),
.B1(n_23),
.B2(n_24),
.Y(n_112)
);

AO22x1_ASAP7_75t_SL g69 ( 
.A1(n_57),
.A2(n_39),
.B1(n_34),
.B2(n_36),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_69),
.A2(n_89),
.B1(n_55),
.B2(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_70),
.B(n_75),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_39),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_46),
.B(n_18),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_78),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_56),
.B(n_22),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_53),
.B(n_21),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_36),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_81),
.A2(n_55),
.B(n_52),
.Y(n_90)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_21),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_84),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_47),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_34),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_31),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_43),
.B(n_22),
.Y(n_88)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_83),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_85),
.A2(n_52),
.B1(n_55),
.B2(n_44),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_111),
.B1(n_112),
.B2(n_74),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_36),
.C(n_43),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_113),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_29),
.B(n_23),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_97),
.A2(n_26),
.B(n_20),
.Y(n_137)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_41),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_114),
.B(n_81),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_74),
.A2(n_44),
.B1(n_29),
.B2(n_32),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_115),
.A2(n_82),
.B1(n_89),
.B2(n_78),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_108),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_127),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_71),
.B1(n_73),
.B2(n_72),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_107),
.A2(n_59),
.B1(n_69),
.B2(n_80),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_120),
.B(n_124),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_103),
.B(n_77),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_121),
.B(n_2),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_109),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_81),
.B1(n_69),
.B2(n_86),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_140),
.B1(n_100),
.B2(n_99),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_70),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_60),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_125),
.B(n_129),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_126),
.A2(n_136),
.B1(n_92),
.B2(n_102),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_115),
.A2(n_66),
.B1(n_68),
.B2(n_65),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_104),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_62),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_137),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_61),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_131),
.B(n_132),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_95),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_97),
.A2(n_109),
.B1(n_90),
.B2(n_106),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

AND2x6_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_41),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_98),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_32),
.B1(n_26),
.B2(n_68),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_141),
.Y(n_155)
);

OA21x2_ASAP7_75t_L g140 ( 
.A1(n_105),
.A2(n_65),
.B(n_20),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_30),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_31),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_100),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_162),
.B1(n_164),
.B2(n_140),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_118),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_146),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_126),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_99),
.C(n_104),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_2),
.C(n_3),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_138),
.Y(n_154)
);

NAND2x1_ASAP7_75t_SL g175 ( 
.A(n_154),
.B(n_160),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_159),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_92),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_L g161 ( 
.A1(n_124),
.A2(n_91),
.A3(n_30),
.B1(n_31),
.B2(n_102),
.C1(n_6),
.C2(n_7),
.Y(n_161)
);

OAI321xp33_ASAP7_75t_L g172 ( 
.A1(n_161),
.A2(n_140),
.A3(n_137),
.B1(n_133),
.B2(n_127),
.C(n_117),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_128),
.Y(n_163)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

OAI22x1_ASAP7_75t_L g164 ( 
.A1(n_134),
.A2(n_91),
.B1(n_30),
.B2(n_4),
.Y(n_164)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_139),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_166),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_30),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_167),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_119),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_168),
.A2(n_116),
.B1(n_149),
.B2(n_136),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_170),
.A2(n_173),
.B1(n_174),
.B2(n_188),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_171),
.B(n_182),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_172),
.A2(n_164),
.B1(n_150),
.B2(n_168),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_145),
.A2(n_123),
.B1(n_130),
.B2(n_135),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_149),
.A2(n_135),
.B1(n_120),
.B2(n_126),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_178),
.Y(n_200)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_183),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_144),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_5),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_143),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_14),
.C(n_9),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_162),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_147),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_189),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_195),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_180),
.A2(n_185),
.B1(n_147),
.B2(n_152),
.Y(n_194)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_152),
.B(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_189),
.Y(n_196)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_184),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_180),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_198),
.B(n_199),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_176),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_202),
.B(n_204),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_143),
.B(n_160),
.Y(n_203)
);

AOI211xp5_ASAP7_75t_L g208 ( 
.A1(n_203),
.A2(n_206),
.B(n_174),
.C(n_188),
.Y(n_208)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_205),
.A2(n_186),
.B1(n_178),
.B2(n_181),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_179),
.A2(n_167),
.B(n_158),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_177),
.C(n_163),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_211),
.Y(n_220)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_201),
.A2(n_185),
.B1(n_173),
.B2(n_170),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_201),
.B1(n_191),
.B2(n_198),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_167),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_217),
.C(n_218),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_144),
.C(n_166),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_183),
.Y(n_221)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_213),
.A2(n_195),
.B(n_192),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_224),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_190),
.C(n_203),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_210),
.A2(n_193),
.B(n_196),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_225),
.B(n_226),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_210),
.A2(n_191),
.B(n_154),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_229),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_219),
.A2(n_155),
.B(n_206),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_228),
.A2(n_209),
.B1(n_218),
.B2(n_208),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_235),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_215),
.C(n_212),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_234),
.C(n_230),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_194),
.Y(n_233)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_233),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_220),
.B(n_211),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_155),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_239),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_216),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_240),
.A2(n_8),
.B(n_11),
.Y(n_247)
);

AOI21x1_ASAP7_75t_L g241 ( 
.A1(n_237),
.A2(n_231),
.B(n_11),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_241),
.A2(n_8),
.B(n_11),
.Y(n_246)
);

INVxp67_ASAP7_75t_SL g244 ( 
.A(n_242),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_246),
.Y(n_250)
);

NOR2xp67_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_12),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_SL g248 ( 
.A1(n_245),
.A2(n_243),
.B(n_240),
.C(n_239),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_248),
.A2(n_249),
.B(n_12),
.Y(n_252)
);

OAI311xp33_ASAP7_75t_L g251 ( 
.A1(n_250),
.A2(n_12),
.A3(n_13),
.B1(n_14),
.C1(n_244),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_252),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_13),
.Y(n_254)
);


endmodule