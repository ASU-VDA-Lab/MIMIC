module fake_netlist_1_12098_n_1067 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_300, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_292, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_297, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_291, n_170, n_294, n_40, n_111, n_157, n_296, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_295, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_298, n_283, n_299, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_293, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_301, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1067);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_300;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_292;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_297;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_291;
input n_170;
input n_294;
input n_40;
input n_111;
input n_157;
input n_296;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_295;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_298;
input n_283;
input n_299;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_293;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_301;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1067;
wire n_663;
wire n_707;
wire n_791;
wire n_513;
wire n_361;
wire n_963;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_964;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_938;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_572;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_975;
wire n_303;
wire n_1042;
wire n_968;
wire n_437;
wire n_512;
wire n_326;
wire n_333;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_529;
wire n_455;
wire n_1011;
wire n_1025;
wire n_630;
wire n_511;
wire n_1002;
wire n_467;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_844;
wire n_818;
wire n_1018;
wire n_738;
wire n_979;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_506;
wire n_533;
wire n_490;
wire n_393;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_950;
wire n_935;
wire n_460;
wire n_1046;
wire n_478;
wire n_482;
wire n_415;
wire n_703;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_995;
wire n_813;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_501;
wire n_871;
wire n_803;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_1020;
wire n_982;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_990;
wire n_751;
wire n_941;
wire n_626;
wire n_800;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_621;
wire n_423;
wire n_342;
wire n_666;
wire n_880;
wire n_799;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_806;
wire n_881;
wire n_539;
wire n_1055;
wire n_1066;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_363;
wire n_315;
wire n_409;
wire n_733;
wire n_861;
wire n_654;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_1060;
wire n_908;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_553;
wire n_440;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_811;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_924;
wire n_947;
wire n_1043;
wire n_912;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_1007;
wire n_1027;
wire n_831;
wire n_859;
wire n_1040;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_967;
wire n_504;
wire n_581;
wire n_458;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_819;
wire n_405;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_992;
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_118), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_27), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_124), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_135), .Y(n_305) );
BUFx3_ASAP7_75t_L g306 ( .A(n_282), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_178), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_295), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_182), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_143), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_31), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_25), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_223), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_188), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_241), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_206), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_112), .Y(n_317) );
CKINVDCx16_ASAP7_75t_R g318 ( .A(n_216), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_221), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_68), .Y(n_320) );
INVxp67_ASAP7_75t_L g321 ( .A(n_4), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_298), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_281), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_18), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_3), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_286), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_197), .Y(n_327) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_233), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_63), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_37), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_70), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_265), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_210), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_77), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_132), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_71), .Y(n_336) );
INVx2_ASAP7_75t_SL g337 ( .A(n_201), .Y(n_337) );
BUFx3_ASAP7_75t_L g338 ( .A(n_29), .Y(n_338) );
INVx1_ASAP7_75t_SL g339 ( .A(n_45), .Y(n_339) );
CKINVDCx16_ASAP7_75t_R g340 ( .A(n_260), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_164), .B(n_94), .Y(n_341) );
INVx1_ASAP7_75t_SL g342 ( .A(n_189), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_8), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_31), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_155), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_122), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_121), .B(n_249), .Y(n_347) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_44), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_86), .Y(n_349) );
BUFx2_ASAP7_75t_L g350 ( .A(n_84), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_151), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_195), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_280), .Y(n_353) );
BUFx10_ASAP7_75t_L g354 ( .A(n_113), .Y(n_354) );
INVxp33_ASAP7_75t_SL g355 ( .A(n_252), .Y(n_355) );
CKINVDCx20_ASAP7_75t_R g356 ( .A(n_287), .Y(n_356) );
INVxp67_ASAP7_75t_SL g357 ( .A(n_52), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_78), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_34), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_8), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_212), .Y(n_361) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_38), .Y(n_362) );
CKINVDCx14_ASAP7_75t_R g363 ( .A(n_40), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_158), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_239), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_203), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_17), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_104), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_33), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_215), .Y(n_370) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_146), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_248), .Y(n_372) );
INVxp67_ASAP7_75t_L g373 ( .A(n_23), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_120), .Y(n_374) );
CKINVDCx20_ASAP7_75t_R g375 ( .A(n_184), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_159), .Y(n_376) );
INVx1_ASAP7_75t_SL g377 ( .A(n_172), .Y(n_377) );
NOR2xp67_ASAP7_75t_L g378 ( .A(n_22), .B(n_217), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_108), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_190), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_236), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_148), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_131), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_272), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_199), .Y(n_385) );
CKINVDCx14_ASAP7_75t_R g386 ( .A(n_245), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_51), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_76), .Y(n_388) );
CKINVDCx14_ASAP7_75t_R g389 ( .A(n_279), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_227), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_293), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_264), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_114), .Y(n_393) );
NOR2xp67_ASAP7_75t_L g394 ( .A(n_55), .B(n_46), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_128), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_27), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_246), .Y(n_397) );
BUFx10_ASAP7_75t_L g398 ( .A(n_299), .Y(n_398) );
INVxp67_ASAP7_75t_SL g399 ( .A(n_105), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_251), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_255), .Y(n_401) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_288), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_127), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_26), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_93), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_41), .Y(n_406) );
INVx4_ASAP7_75t_R g407 ( .A(n_6), .Y(n_407) );
CKINVDCx14_ASAP7_75t_R g408 ( .A(n_261), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_74), .Y(n_409) );
INVxp67_ASAP7_75t_L g410 ( .A(n_247), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_205), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_225), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_213), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_130), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_4), .Y(n_415) );
CKINVDCx5p33_ASAP7_75t_R g416 ( .A(n_87), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_193), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_161), .Y(n_418) );
NOR2xp67_ASAP7_75t_L g419 ( .A(n_183), .B(n_48), .Y(n_419) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_254), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_99), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_250), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_269), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_156), .Y(n_424) );
BUFx2_ASAP7_75t_L g425 ( .A(n_67), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_301), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_97), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_115), .Y(n_428) );
CKINVDCx5p33_ASAP7_75t_R g429 ( .A(n_207), .Y(n_429) );
CKINVDCx5p33_ASAP7_75t_R g430 ( .A(n_32), .Y(n_430) );
CKINVDCx5p33_ASAP7_75t_R g431 ( .A(n_2), .Y(n_431) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_294), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_244), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_176), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_79), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_157), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_277), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_297), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_242), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_75), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_166), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_17), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_142), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_234), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_119), .Y(n_445) );
INVx2_ASAP7_75t_SL g446 ( .A(n_117), .Y(n_446) );
CKINVDCx5p33_ASAP7_75t_R g447 ( .A(n_259), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_7), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_25), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_13), .Y(n_450) );
CKINVDCx5p33_ASAP7_75t_R g451 ( .A(n_88), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g452 ( .A(n_18), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_137), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_141), .Y(n_454) );
CKINVDCx5p33_ASAP7_75t_R g455 ( .A(n_109), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_59), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_162), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_202), .Y(n_458) );
BUFx3_ASAP7_75t_L g459 ( .A(n_14), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_35), .Y(n_460) );
INVx1_ASAP7_75t_SL g461 ( .A(n_95), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_14), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_318), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_326), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_358), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_372), .Y(n_466) );
BUFx3_ASAP7_75t_L g467 ( .A(n_306), .Y(n_467) );
AND2x4_ASAP7_75t_L g468 ( .A(n_362), .B(n_0), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_303), .B(n_0), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_362), .Y(n_470) );
INVx3_ASAP7_75t_L g471 ( .A(n_354), .Y(n_471) );
AND2x4_ASAP7_75t_L g472 ( .A(n_387), .B(n_1), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_426), .Y(n_473) );
BUFx2_ASAP7_75t_L g474 ( .A(n_338), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_387), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_336), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_335), .B(n_1), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_350), .B(n_2), .Y(n_478) );
INVx3_ASAP7_75t_L g479 ( .A(n_354), .Y(n_479) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_313), .Y(n_480) );
OA21x2_ASAP7_75t_L g481 ( .A1(n_305), .A2(n_39), .B(n_36), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_427), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_321), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_425), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_450), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_340), .B(n_3), .Y(n_486) );
INVx3_ASAP7_75t_L g487 ( .A(n_398), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_337), .B(n_446), .Y(n_488) );
OAI21x1_ASAP7_75t_L g489 ( .A1(n_456), .A2(n_43), .B(n_42), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_321), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_363), .B(n_5), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_307), .Y(n_492) );
XNOR2xp5_ASAP7_75t_L g493 ( .A(n_311), .B(n_5), .Y(n_493) );
INVx6_ASAP7_75t_L g494 ( .A(n_398), .Y(n_494) );
NAND3xp33_ASAP7_75t_L g495 ( .A(n_470), .B(n_373), .C(n_324), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_463), .Y(n_496) );
BUFx10_ASAP7_75t_L g497 ( .A(n_468), .Y(n_497) );
AO21x2_ASAP7_75t_L g498 ( .A1(n_489), .A2(n_314), .B(n_309), .Y(n_498) );
BUFx2_ASAP7_75t_L g499 ( .A(n_463), .Y(n_499) );
INVx2_ASAP7_75t_SL g500 ( .A(n_494), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_467), .Y(n_501) );
BUFx3_ASAP7_75t_L g502 ( .A(n_471), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_464), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_471), .B(n_410), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_464), .Y(n_505) );
INVx8_ASAP7_75t_L g506 ( .A(n_468), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_467), .Y(n_507) );
INVx3_ASAP7_75t_L g508 ( .A(n_468), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_465), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_472), .A2(n_373), .B1(n_367), .B2(n_312), .Y(n_510) );
INVx5_ASAP7_75t_L g511 ( .A(n_480), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_471), .B(n_410), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_465), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_466), .Y(n_514) );
AOI22xp33_ASAP7_75t_SL g515 ( .A1(n_472), .A2(n_343), .B1(n_344), .B2(n_325), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_466), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_473), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_472), .A2(n_396), .B1(n_431), .B2(n_404), .Y(n_518) );
INVx1_ASAP7_75t_SL g519 ( .A(n_486), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_473), .Y(n_520) );
INVx2_ASAP7_75t_SL g521 ( .A(n_506), .Y(n_521) );
INVx2_ASAP7_75t_SL g522 ( .A(n_506), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_498), .A2(n_488), .B(n_489), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_506), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_500), .B(n_502), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_502), .B(n_494), .Y(n_526) );
BUFx3_ASAP7_75t_L g527 ( .A(n_499), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_519), .B(n_483), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_508), .Y(n_529) );
INVxp67_ASAP7_75t_L g530 ( .A(n_519), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_497), .B(n_491), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_508), .B(n_475), .Y(n_532) );
INVx3_ASAP7_75t_L g533 ( .A(n_497), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_515), .B(n_491), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_515), .A2(n_478), .B1(n_490), .B2(n_492), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_504), .B(n_478), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_510), .A2(n_476), .B1(n_484), .B2(n_356), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_518), .A2(n_479), .B1(n_487), .B2(n_494), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_498), .A2(n_477), .B(n_481), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_495), .B(n_479), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_504), .B(n_479), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_503), .A2(n_492), .B1(n_482), .B2(n_360), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_512), .B(n_487), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_505), .Y(n_544) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_512), .A2(n_482), .B(n_469), .C(n_448), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_496), .B(n_474), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_514), .B(n_357), .Y(n_547) );
BUFx3_ASAP7_75t_L g548 ( .A(n_501), .Y(n_548) );
NAND2x1_ASAP7_75t_L g549 ( .A(n_507), .B(n_407), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_516), .B(n_485), .Y(n_550) );
INVx2_ASAP7_75t_SL g551 ( .A(n_509), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_513), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_517), .B(n_357), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_520), .Y(n_554) );
INVx3_ASAP7_75t_L g555 ( .A(n_511), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_511), .Y(n_556) );
AND2x4_ASAP7_75t_L g557 ( .A(n_511), .B(n_352), .Y(n_557) );
NAND2xp33_ASAP7_75t_L g558 ( .A(n_521), .B(n_371), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g559 ( .A1(n_536), .A2(n_399), .B(n_462), .C(n_415), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_529), .Y(n_560) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_527), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_530), .Y(n_562) );
OAI21xp33_ASAP7_75t_L g563 ( .A1(n_528), .A2(n_493), .B(n_449), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_523), .A2(n_481), .B(n_399), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_536), .B(n_442), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_546), .B(n_493), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_554), .Y(n_567) );
O2A1O1Ixp33_ASAP7_75t_SL g568 ( .A1(n_545), .A2(n_347), .B(n_316), .C(n_319), .Y(n_568) );
OAI21xp5_ASAP7_75t_L g569 ( .A1(n_539), .A2(n_481), .B(n_320), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_530), .B(n_452), .Y(n_570) );
A2O1A1Ixp33_ASAP7_75t_L g571 ( .A1(n_523), .A2(n_378), .B(n_459), .C(n_322), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_552), .Y(n_572) );
NOR3xp33_ASAP7_75t_L g573 ( .A(n_537), .B(n_389), .C(n_386), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_539), .A2(n_329), .B(n_315), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_532), .B(n_355), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_532), .B(n_375), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_541), .A2(n_332), .B(n_331), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_551), .Y(n_578) );
OAI21xp33_ASAP7_75t_L g579 ( .A1(n_535), .A2(n_408), .B(n_304), .Y(n_579) );
INVx3_ASAP7_75t_L g580 ( .A(n_548), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_543), .A2(n_345), .B(n_333), .Y(n_581) );
INVx3_ASAP7_75t_L g582 ( .A(n_555), .Y(n_582) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_522), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_538), .B(n_444), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_531), .A2(n_351), .B(n_349), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_544), .Y(n_586) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_540), .A2(n_359), .B(n_353), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_534), .A2(n_458), .B1(n_366), .B2(n_369), .Y(n_588) );
OAI21x1_ASAP7_75t_L g589 ( .A1(n_549), .A2(n_370), .B(n_361), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_547), .B(n_302), .Y(n_590) );
AOI21xp5_ASAP7_75t_L g591 ( .A1(n_547), .A2(n_379), .B(n_376), .Y(n_591) );
OA22x2_ASAP7_75t_L g592 ( .A1(n_557), .A2(n_382), .B1(n_390), .B2(n_381), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_553), .B(n_392), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_553), .A2(n_401), .B(n_395), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_533), .B(n_308), .Y(n_595) );
A2O1A1Ixp33_ASAP7_75t_L g596 ( .A1(n_550), .A2(n_403), .B(n_411), .C(n_405), .Y(n_596) );
O2A1O1Ixp33_ASAP7_75t_L g597 ( .A1(n_542), .A2(n_414), .B(n_422), .C(n_413), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_524), .B(n_310), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_533), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_562), .B(n_542), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_559), .B(n_526), .Y(n_601) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_574), .A2(n_525), .B(n_556), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_566), .B(n_555), .Y(n_603) );
AO31x2_ASAP7_75t_L g604 ( .A1(n_571), .A2(n_428), .A3(n_438), .B(n_434), .Y(n_604) );
AND2x4_ASAP7_75t_L g605 ( .A(n_578), .B(n_394), .Y(n_605) );
OAI22x1_ASAP7_75t_L g606 ( .A1(n_561), .A2(n_441), .B1(n_443), .B2(n_439), .Y(n_606) );
OAI22x1_ASAP7_75t_L g607 ( .A1(n_584), .A2(n_453), .B1(n_460), .B2(n_445), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g608 ( .A1(n_564), .A2(n_419), .B(n_341), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_586), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_567), .Y(n_610) );
OAI21xp5_ASAP7_75t_L g611 ( .A1(n_591), .A2(n_342), .B(n_339), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_576), .B(n_317), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_565), .B(n_323), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_560), .Y(n_614) );
O2A1O1Ixp5_ASAP7_75t_L g615 ( .A1(n_569), .A2(n_461), .B(n_377), .C(n_327), .Y(n_615) );
OAI21xp5_ASAP7_75t_L g616 ( .A1(n_594), .A2(n_334), .B(n_330), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_575), .B(n_346), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_572), .Y(n_618) );
AO31x2_ASAP7_75t_L g619 ( .A1(n_596), .A2(n_480), .A3(n_328), .B(n_348), .Y(n_619) );
OAI21x1_ASAP7_75t_L g620 ( .A1(n_589), .A2(n_328), .B(n_313), .Y(n_620) );
OAI21xp5_ASAP7_75t_SL g621 ( .A1(n_573), .A2(n_328), .B(n_313), .Y(n_621) );
A2O1A1Ixp33_ASAP7_75t_L g622 ( .A1(n_597), .A2(n_402), .B(n_420), .C(n_348), .Y(n_622) );
AO31x2_ASAP7_75t_L g623 ( .A1(n_593), .A2(n_480), .A3(n_402), .B(n_420), .Y(n_623) );
NOR2xp67_ASAP7_75t_SL g624 ( .A(n_583), .B(n_364), .Y(n_624) );
AOI221x1_ASAP7_75t_L g625 ( .A1(n_579), .A2(n_480), .B1(n_420), .B2(n_402), .C(n_348), .Y(n_625) );
NOR2xp67_ASAP7_75t_L g626 ( .A(n_563), .B(n_7), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_593), .A2(n_368), .B(n_365), .Y(n_627) );
OAI21x1_ASAP7_75t_L g628 ( .A1(n_582), .A2(n_49), .B(n_47), .Y(n_628) );
AO21x1_ASAP7_75t_L g629 ( .A1(n_587), .A2(n_53), .B(n_50), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g630 ( .A1(n_577), .A2(n_380), .B(n_374), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_588), .B(n_383), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_570), .B(n_384), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_580), .B(n_385), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_580), .B(n_388), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_590), .A2(n_393), .B(n_391), .Y(n_635) );
OAI21x1_ASAP7_75t_L g636 ( .A1(n_582), .A2(n_56), .B(n_54), .Y(n_636) );
OA21x2_ASAP7_75t_L g637 ( .A1(n_581), .A2(n_585), .B(n_599), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_592), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_568), .A2(n_400), .B(n_397), .Y(n_639) );
NOR2xp67_ASAP7_75t_L g640 ( .A(n_598), .B(n_9), .Y(n_640) );
INVxp67_ASAP7_75t_L g641 ( .A(n_558), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_583), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_595), .Y(n_643) );
INVx1_ASAP7_75t_SL g644 ( .A(n_561), .Y(n_644) );
OAI21x1_ASAP7_75t_L g645 ( .A1(n_620), .A2(n_58), .B(n_57), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_618), .Y(n_646) );
OAI21x1_ASAP7_75t_L g647 ( .A1(n_628), .A2(n_61), .B(n_60), .Y(n_647) );
OAI21x1_ASAP7_75t_L g648 ( .A1(n_636), .A2(n_64), .B(n_62), .Y(n_648) );
AO21x2_ASAP7_75t_L g649 ( .A1(n_608), .A2(n_66), .B(n_65), .Y(n_649) );
CKINVDCx5p33_ASAP7_75t_R g650 ( .A(n_642), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_610), .Y(n_651) );
AND2x2_ASAP7_75t_SL g652 ( .A(n_638), .B(n_9), .Y(n_652) );
OR2x2_ASAP7_75t_L g653 ( .A(n_644), .B(n_10), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_614), .Y(n_654) );
OAI21xp5_ASAP7_75t_L g655 ( .A1(n_615), .A2(n_409), .B(n_406), .Y(n_655) );
OA21x2_ASAP7_75t_L g656 ( .A1(n_625), .A2(n_416), .B(n_412), .Y(n_656) );
NOR2xp67_ASAP7_75t_L g657 ( .A(n_641), .B(n_69), .Y(n_657) );
INVx2_ASAP7_75t_SL g658 ( .A(n_603), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_643), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_600), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_626), .A2(n_457), .B1(n_455), .B2(n_454), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_602), .A2(n_601), .B(n_611), .Y(n_662) );
OAI21x1_ASAP7_75t_L g663 ( .A1(n_629), .A2(n_73), .B(n_72), .Y(n_663) );
NAND2x1p5_ASAP7_75t_L g664 ( .A(n_624), .B(n_10), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_637), .Y(n_665) );
OAI21x1_ASAP7_75t_L g666 ( .A1(n_621), .A2(n_81), .B(n_80), .Y(n_666) );
OAI21x1_ASAP7_75t_L g667 ( .A1(n_627), .A2(n_83), .B(n_82), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_640), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_607), .B(n_11), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_616), .B(n_12), .Y(n_670) );
BUFx10_ASAP7_75t_L g671 ( .A(n_605), .Y(n_671) );
OAI21x1_ASAP7_75t_L g672 ( .A1(n_639), .A2(n_89), .B(n_85), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_604), .B(n_12), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_622), .A2(n_418), .B(n_417), .Y(n_674) );
OA21x2_ASAP7_75t_L g675 ( .A1(n_623), .A2(n_423), .B(n_421), .Y(n_675) );
NOR2xp33_ASAP7_75t_R g676 ( .A(n_633), .B(n_13), .Y(n_676) );
OAI21x1_ASAP7_75t_L g677 ( .A1(n_635), .A2(n_91), .B(n_90), .Y(n_677) );
INVxp67_ASAP7_75t_L g678 ( .A(n_606), .Y(n_678) );
NOR2x1_ASAP7_75t_SL g679 ( .A(n_634), .B(n_15), .Y(n_679) );
OAI21x1_ASAP7_75t_L g680 ( .A1(n_630), .A2(n_96), .B(n_92), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g681 ( .A1(n_605), .A2(n_429), .B(n_424), .Y(n_681) );
OAI21x1_ASAP7_75t_L g682 ( .A1(n_623), .A2(n_632), .B(n_612), .Y(n_682) );
OA21x2_ASAP7_75t_L g683 ( .A1(n_623), .A2(n_432), .B(n_430), .Y(n_683) );
INVx2_ASAP7_75t_SL g684 ( .A(n_604), .Y(n_684) );
OA21x2_ASAP7_75t_L g685 ( .A1(n_619), .A2(n_435), .B(n_433), .Y(n_685) );
OA21x2_ASAP7_75t_L g686 ( .A1(n_619), .A2(n_437), .B(n_436), .Y(n_686) );
INVx3_ASAP7_75t_L g687 ( .A(n_613), .Y(n_687) );
OAI21x1_ASAP7_75t_L g688 ( .A1(n_617), .A2(n_100), .B(n_98), .Y(n_688) );
OR2x2_ASAP7_75t_L g689 ( .A(n_631), .B(n_16), .Y(n_689) );
OA21x2_ASAP7_75t_L g690 ( .A1(n_608), .A2(n_447), .B(n_440), .Y(n_690) );
OA21x2_ASAP7_75t_L g691 ( .A1(n_608), .A2(n_451), .B(n_102), .Y(n_691) );
NAND2x1p5_ASAP7_75t_L g692 ( .A(n_624), .B(n_19), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_609), .Y(n_693) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_609), .Y(n_694) );
INVx1_ASAP7_75t_SL g695 ( .A(n_642), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_609), .Y(n_696) );
AO21x2_ASAP7_75t_L g697 ( .A1(n_608), .A2(n_103), .B(n_101), .Y(n_697) );
AND2x4_ASAP7_75t_L g698 ( .A(n_643), .B(n_19), .Y(n_698) );
OAI21x1_ASAP7_75t_L g699 ( .A1(n_620), .A2(n_107), .B(n_106), .Y(n_699) );
BUFx3_ASAP7_75t_L g700 ( .A(n_642), .Y(n_700) );
AND2x4_ASAP7_75t_L g701 ( .A(n_654), .B(n_20), .Y(n_701) );
BUFx3_ASAP7_75t_L g702 ( .A(n_700), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_665), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_693), .Y(n_704) );
AND2x4_ASAP7_75t_L g705 ( .A(n_694), .B(n_20), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_646), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_696), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_646), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_651), .Y(n_709) );
OR2x2_ASAP7_75t_L g710 ( .A(n_695), .B(n_21), .Y(n_710) );
INVx3_ASAP7_75t_L g711 ( .A(n_698), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_694), .Y(n_712) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_700), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_660), .B(n_21), .Y(n_714) );
INVx3_ASAP7_75t_L g715 ( .A(n_698), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_673), .Y(n_716) );
INVx3_ASAP7_75t_L g717 ( .A(n_664), .Y(n_717) );
INVx3_ASAP7_75t_L g718 ( .A(n_664), .Y(n_718) );
INVxp67_ASAP7_75t_L g719 ( .A(n_652), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_673), .Y(n_720) );
AND2x4_ASAP7_75t_L g721 ( .A(n_658), .B(n_668), .Y(n_721) );
AND2x4_ASAP7_75t_L g722 ( .A(n_687), .B(n_23), .Y(n_722) );
OAI21xp33_ASAP7_75t_SL g723 ( .A1(n_652), .A2(n_24), .B(n_26), .Y(n_723) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_684), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_669), .B(n_24), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_695), .B(n_28), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_692), .Y(n_727) );
BUFx6f_ASAP7_75t_L g728 ( .A(n_666), .Y(n_728) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_678), .Y(n_729) );
INVx1_ASAP7_75t_SL g730 ( .A(n_671), .Y(n_730) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_678), .Y(n_731) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_685), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_662), .B(n_30), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_689), .Y(n_734) );
BUFx3_ASAP7_75t_L g735 ( .A(n_650), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_647), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_679), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_671), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_670), .B(n_30), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_670), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_653), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_685), .Y(n_742) );
BUFx3_ASAP7_75t_L g743 ( .A(n_677), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_661), .A2(n_110), .B1(n_111), .B2(n_116), .Y(n_744) );
BUFx2_ASAP7_75t_L g745 ( .A(n_676), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_648), .Y(n_746) );
AO21x2_ASAP7_75t_L g747 ( .A1(n_682), .A2(n_123), .B(n_125), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_676), .Y(n_748) );
BUFx3_ASAP7_75t_L g749 ( .A(n_667), .Y(n_749) );
OAI21x1_ASAP7_75t_L g750 ( .A1(n_645), .A2(n_126), .B(n_129), .Y(n_750) );
OA21x2_ASAP7_75t_L g751 ( .A1(n_663), .A2(n_133), .B(n_134), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_657), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_657), .Y(n_753) );
INVxp67_ASAP7_75t_L g754 ( .A(n_661), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_690), .Y(n_755) );
INVx8_ASAP7_75t_L g756 ( .A(n_681), .Y(n_756) );
AOI21x1_ASAP7_75t_L g757 ( .A1(n_691), .A2(n_300), .B(n_138), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_686), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_675), .Y(n_759) );
INVxp33_ASAP7_75t_SL g760 ( .A(n_655), .Y(n_760) );
AO21x2_ASAP7_75t_L g761 ( .A1(n_655), .A2(n_136), .B(n_139), .Y(n_761) );
OAI21x1_ASAP7_75t_L g762 ( .A1(n_699), .A2(n_140), .B(n_144), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_681), .B(n_145), .Y(n_763) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_683), .Y(n_764) );
INVx3_ASAP7_75t_L g765 ( .A(n_672), .Y(n_765) );
OR2x2_ASAP7_75t_L g766 ( .A(n_683), .B(n_697), .Y(n_766) );
AND2x4_ASAP7_75t_L g767 ( .A(n_688), .B(n_147), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_680), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_674), .B(n_149), .Y(n_769) );
INVxp67_ASAP7_75t_L g770 ( .A(n_697), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_649), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_649), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_674), .B(n_150), .Y(n_773) );
AND2x2_ASAP7_75t_L g774 ( .A(n_656), .B(n_152), .Y(n_774) );
AND2x2_ASAP7_75t_L g775 ( .A(n_656), .B(n_153), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_659), .Y(n_776) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_694), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_665), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_694), .B(n_154), .Y(n_779) );
INVx2_ASAP7_75t_L g780 ( .A(n_665), .Y(n_780) );
INVx2_ASAP7_75t_SL g781 ( .A(n_735), .Y(n_781) );
BUFx3_ASAP7_75t_L g782 ( .A(n_702), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_704), .Y(n_783) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_777), .Y(n_784) );
INVx2_ASAP7_75t_SL g785 ( .A(n_735), .Y(n_785) );
BUFx2_ASAP7_75t_L g786 ( .A(n_705), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_706), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_776), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_707), .Y(n_789) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_724), .Y(n_790) );
OR2x2_ASAP7_75t_L g791 ( .A(n_712), .B(n_160), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_725), .B(n_163), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_719), .A2(n_165), .B1(n_167), .B2(n_168), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_709), .Y(n_794) );
INVx2_ASAP7_75t_L g795 ( .A(n_708), .Y(n_795) );
INVx2_ASAP7_75t_L g796 ( .A(n_703), .Y(n_796) );
INVxp67_ASAP7_75t_L g797 ( .A(n_729), .Y(n_797) );
BUFx2_ASAP7_75t_L g798 ( .A(n_705), .Y(n_798) );
AND2x4_ASAP7_75t_L g799 ( .A(n_711), .B(n_169), .Y(n_799) );
AND2x4_ASAP7_75t_SL g800 ( .A(n_717), .B(n_170), .Y(n_800) );
AND2x2_ASAP7_75t_L g801 ( .A(n_726), .B(n_171), .Y(n_801) );
INVxp67_ASAP7_75t_L g802 ( .A(n_729), .Y(n_802) );
OAI21x1_ASAP7_75t_SL g803 ( .A1(n_727), .A2(n_173), .B(n_174), .Y(n_803) );
AND2x2_ASAP7_75t_L g804 ( .A(n_741), .B(n_175), .Y(n_804) );
AOI211x1_ASAP7_75t_L g805 ( .A1(n_748), .A2(n_177), .B(n_179), .C(n_180), .Y(n_805) );
BUFx2_ASAP7_75t_L g806 ( .A(n_702), .Y(n_806) );
AND2x2_ASAP7_75t_L g807 ( .A(n_734), .B(n_181), .Y(n_807) );
INVx2_ASAP7_75t_L g808 ( .A(n_778), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_722), .B(n_185), .Y(n_809) );
OAI221xp5_ASAP7_75t_L g810 ( .A1(n_723), .A2(n_186), .B1(n_187), .B2(n_191), .C(n_192), .Y(n_810) );
AND2x2_ASAP7_75t_L g811 ( .A(n_722), .B(n_194), .Y(n_811) );
OR2x2_ASAP7_75t_L g812 ( .A(n_731), .B(n_296), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_719), .A2(n_196), .B1(n_198), .B2(n_200), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_731), .Y(n_814) );
INVx2_ASAP7_75t_SL g815 ( .A(n_713), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_780), .Y(n_816) );
INVx3_ASAP7_75t_L g817 ( .A(n_717), .Y(n_817) );
INVxp33_ASAP7_75t_SL g818 ( .A(n_745), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_714), .Y(n_819) );
INVx3_ASAP7_75t_L g820 ( .A(n_718), .Y(n_820) );
BUFx2_ASAP7_75t_L g821 ( .A(n_713), .Y(n_821) );
INVx4_ASAP7_75t_L g822 ( .A(n_718), .Y(n_822) );
HB1xp67_ASAP7_75t_L g823 ( .A(n_724), .Y(n_823) );
BUFx3_ASAP7_75t_L g824 ( .A(n_713), .Y(n_824) );
AND2x2_ASAP7_75t_L g825 ( .A(n_701), .B(n_204), .Y(n_825) );
INVxp67_ASAP7_75t_SL g826 ( .A(n_764), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_740), .B(n_208), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_730), .B(n_209), .Y(n_828) );
INVx3_ASAP7_75t_L g829 ( .A(n_711), .Y(n_829) );
INVx4_ASAP7_75t_L g830 ( .A(n_715), .Y(n_830) );
AND2x2_ASAP7_75t_L g831 ( .A(n_730), .B(n_211), .Y(n_831) );
AND2x2_ASAP7_75t_L g832 ( .A(n_710), .B(n_214), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_714), .Y(n_833) );
AND2x2_ASAP7_75t_L g834 ( .A(n_721), .B(n_218), .Y(n_834) );
INVxp67_ASAP7_75t_SL g835 ( .A(n_764), .Y(n_835) );
NOR2xp67_ASAP7_75t_L g836 ( .A(n_737), .B(n_219), .Y(n_836) );
HB1xp67_ASAP7_75t_L g837 ( .A(n_716), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_739), .Y(n_838) );
AND2x2_ASAP7_75t_L g839 ( .A(n_754), .B(n_220), .Y(n_839) );
AND2x2_ASAP7_75t_L g840 ( .A(n_754), .B(n_222), .Y(n_840) );
NOR2x1_ASAP7_75t_SL g841 ( .A(n_779), .B(n_738), .Y(n_841) );
INVx2_ASAP7_75t_L g842 ( .A(n_736), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_739), .Y(n_843) );
AND2x4_ASAP7_75t_L g844 ( .A(n_755), .B(n_224), .Y(n_844) );
NOR2xp33_ASAP7_75t_L g845 ( .A(n_760), .B(n_226), .Y(n_845) );
NOR2xp67_ASAP7_75t_L g846 ( .A(n_744), .B(n_228), .Y(n_846) );
OR2x6_ASAP7_75t_L g847 ( .A(n_756), .B(n_229), .Y(n_847) );
AOI22xp33_ASAP7_75t_SL g848 ( .A1(n_760), .A2(n_230), .B1(n_231), .B2(n_232), .Y(n_848) );
HB1xp67_ASAP7_75t_L g849 ( .A(n_720), .Y(n_849) );
AND2x2_ASAP7_75t_L g850 ( .A(n_763), .B(n_235), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_733), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_756), .A2(n_237), .B1(n_238), .B2(n_240), .Y(n_852) );
AND2x2_ASAP7_75t_L g853 ( .A(n_773), .B(n_243), .Y(n_853) );
HB1xp67_ASAP7_75t_L g854 ( .A(n_732), .Y(n_854) );
BUFx6f_ASAP7_75t_L g855 ( .A(n_728), .Y(n_855) );
AOI22xp33_ASAP7_75t_SL g856 ( .A1(n_756), .A2(n_253), .B1(n_256), .B2(n_257), .Y(n_856) );
INVx2_ASAP7_75t_L g857 ( .A(n_746), .Y(n_857) );
NOR2x1_ASAP7_75t_L g858 ( .A(n_761), .B(n_258), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_752), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_753), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_732), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_769), .Y(n_862) );
INVx2_ASAP7_75t_L g863 ( .A(n_746), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_774), .Y(n_864) );
HB1xp67_ASAP7_75t_L g865 ( .A(n_759), .Y(n_865) );
INVxp67_ASAP7_75t_SL g866 ( .A(n_742), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_758), .B(n_262), .Y(n_867) );
INVx2_ASAP7_75t_L g868 ( .A(n_775), .Y(n_868) );
AND2x2_ASAP7_75t_SL g869 ( .A(n_766), .B(n_263), .Y(n_869) );
AND2x2_ASAP7_75t_L g870 ( .A(n_761), .B(n_266), .Y(n_870) );
HB1xp67_ASAP7_75t_L g871 ( .A(n_768), .Y(n_871) );
AND2x4_ASAP7_75t_L g872 ( .A(n_790), .B(n_749), .Y(n_872) );
AND2x2_ASAP7_75t_L g873 ( .A(n_806), .B(n_747), .Y(n_873) );
HB1xp67_ASAP7_75t_L g874 ( .A(n_790), .Y(n_874) );
INVx2_ASAP7_75t_L g875 ( .A(n_783), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_788), .Y(n_876) );
INVx1_ASAP7_75t_SL g877 ( .A(n_782), .Y(n_877) );
OR2x2_ASAP7_75t_L g878 ( .A(n_784), .B(n_772), .Y(n_878) );
INVx2_ASAP7_75t_L g879 ( .A(n_787), .Y(n_879) );
INVx2_ASAP7_75t_L g880 ( .A(n_795), .Y(n_880) );
OR2x2_ASAP7_75t_L g881 ( .A(n_784), .B(n_770), .Y(n_881) );
INVx2_ASAP7_75t_SL g882 ( .A(n_824), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_789), .Y(n_883) );
NOR2x1_ASAP7_75t_L g884 ( .A(n_822), .B(n_767), .Y(n_884) );
NOR2xp33_ASAP7_75t_L g885 ( .A(n_786), .B(n_767), .Y(n_885) );
NOR2x1_ASAP7_75t_L g886 ( .A(n_822), .B(n_749), .Y(n_886) );
INVx4_ASAP7_75t_L g887 ( .A(n_847), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_794), .Y(n_888) );
HB1xp67_ASAP7_75t_L g889 ( .A(n_823), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_814), .Y(n_890) );
BUFx2_ASAP7_75t_L g891 ( .A(n_824), .Y(n_891) );
INVx2_ASAP7_75t_L g892 ( .A(n_796), .Y(n_892) );
HB1xp67_ASAP7_75t_L g893 ( .A(n_854), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_851), .B(n_771), .Y(n_894) );
NOR2xp33_ASAP7_75t_SL g895 ( .A(n_869), .B(n_743), .Y(n_895) );
AND2x2_ASAP7_75t_L g896 ( .A(n_798), .B(n_771), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_837), .Y(n_897) );
HB1xp67_ASAP7_75t_L g898 ( .A(n_854), .Y(n_898) );
AND2x2_ASAP7_75t_L g899 ( .A(n_821), .B(n_765), .Y(n_899) );
NAND2x1_ASAP7_75t_L g900 ( .A(n_847), .B(n_765), .Y(n_900) );
INVx2_ASAP7_75t_L g901 ( .A(n_808), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_849), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_849), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_797), .B(n_728), .Y(n_904) );
NOR2xp33_ASAP7_75t_L g905 ( .A(n_838), .B(n_757), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_802), .Y(n_906) );
HB1xp67_ASAP7_75t_L g907 ( .A(n_865), .Y(n_907) );
AND2x2_ASAP7_75t_L g908 ( .A(n_802), .B(n_751), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_781), .B(n_751), .Y(n_909) );
INVx2_ASAP7_75t_L g910 ( .A(n_816), .Y(n_910) );
INVx3_ASAP7_75t_L g911 ( .A(n_830), .Y(n_911) );
AND2x2_ASAP7_75t_L g912 ( .A(n_785), .B(n_762), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_843), .B(n_750), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_859), .Y(n_914) );
AND2x2_ASAP7_75t_L g915 ( .A(n_860), .B(n_267), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_819), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_833), .Y(n_917) );
AND2x4_ASAP7_75t_L g918 ( .A(n_841), .B(n_268), .Y(n_918) );
AND2x4_ASAP7_75t_SL g919 ( .A(n_830), .B(n_270), .Y(n_919) );
INVx3_ASAP7_75t_L g920 ( .A(n_844), .Y(n_920) );
OR2x2_ASAP7_75t_L g921 ( .A(n_815), .B(n_271), .Y(n_921) );
HB1xp67_ASAP7_75t_L g922 ( .A(n_826), .Y(n_922) );
INVx2_ASAP7_75t_L g923 ( .A(n_861), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_871), .Y(n_924) );
AND2x2_ASAP7_75t_L g925 ( .A(n_839), .B(n_273), .Y(n_925) );
NAND2xp5_ASAP7_75t_SL g926 ( .A(n_869), .B(n_274), .Y(n_926) );
AND2x2_ASAP7_75t_L g927 ( .A(n_840), .B(n_275), .Y(n_927) );
AND2x4_ASAP7_75t_L g928 ( .A(n_829), .B(n_276), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_818), .A2(n_278), .B1(n_283), .B2(n_284), .Y(n_929) );
BUFx3_ASAP7_75t_L g930 ( .A(n_817), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_812), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_862), .B(n_285), .Y(n_932) );
INVxp67_ASAP7_75t_SL g933 ( .A(n_826), .Y(n_933) );
AND2x2_ASAP7_75t_L g934 ( .A(n_829), .B(n_289), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_835), .Y(n_935) );
AND2x2_ASAP7_75t_L g936 ( .A(n_864), .B(n_290), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_835), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_868), .B(n_291), .Y(n_938) );
OR2x2_ASAP7_75t_L g939 ( .A(n_907), .B(n_866), .Y(n_939) );
NOR2x1_ASAP7_75t_L g940 ( .A(n_887), .B(n_820), .Y(n_940) );
AND2x2_ASAP7_75t_L g941 ( .A(n_877), .B(n_817), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_894), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_916), .B(n_818), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_914), .Y(n_944) );
OAI21xp5_ASAP7_75t_L g945 ( .A1(n_926), .A2(n_845), .B(n_848), .Y(n_945) );
NAND4xp25_ASAP7_75t_L g946 ( .A(n_885), .B(n_845), .C(n_805), .D(n_792), .Y(n_946) );
OR2x2_ASAP7_75t_L g947 ( .A(n_874), .B(n_842), .Y(n_947) );
AND2x2_ASAP7_75t_L g948 ( .A(n_876), .B(n_834), .Y(n_948) );
BUFx2_ASAP7_75t_L g949 ( .A(n_911), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_894), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_887), .A2(n_810), .B1(n_848), .B2(n_825), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_875), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_917), .B(n_804), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_879), .Y(n_954) );
OR2x2_ASAP7_75t_L g955 ( .A(n_889), .B(n_857), .Y(n_955) );
AND2x2_ASAP7_75t_L g956 ( .A(n_883), .B(n_832), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_880), .Y(n_957) );
INVxp67_ASAP7_75t_SL g958 ( .A(n_922), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_888), .Y(n_959) );
AND2x4_ASAP7_75t_L g960 ( .A(n_933), .B(n_872), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_896), .B(n_811), .Y(n_961) );
AND2x2_ASAP7_75t_L g962 ( .A(n_890), .B(n_809), .Y(n_962) );
BUFx3_ASAP7_75t_L g963 ( .A(n_891), .Y(n_963) );
INVx1_ASAP7_75t_L g964 ( .A(n_923), .Y(n_964) );
INVx1_ASAP7_75t_L g965 ( .A(n_897), .Y(n_965) );
AND2x4_ASAP7_75t_L g966 ( .A(n_933), .B(n_855), .Y(n_966) );
INVx3_ASAP7_75t_L g967 ( .A(n_911), .Y(n_967) );
AND2x4_ASAP7_75t_L g968 ( .A(n_872), .B(n_855), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_910), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_910), .Y(n_970) );
BUFx2_ASAP7_75t_L g971 ( .A(n_882), .Y(n_971) );
OR2x6_ASAP7_75t_L g972 ( .A(n_900), .B(n_799), .Y(n_972) );
OR2x2_ASAP7_75t_L g973 ( .A(n_902), .B(n_863), .Y(n_973) );
OR2x2_ASAP7_75t_L g974 ( .A(n_903), .B(n_863), .Y(n_974) );
BUFx2_ASAP7_75t_L g975 ( .A(n_930), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_906), .B(n_801), .Y(n_976) );
OR2x2_ASAP7_75t_L g977 ( .A(n_893), .B(n_791), .Y(n_977) );
NAND2x1p5_ASAP7_75t_L g978 ( .A(n_918), .B(n_799), .Y(n_978) );
AND2x4_ASAP7_75t_L g979 ( .A(n_899), .B(n_855), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_892), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_931), .B(n_807), .Y(n_981) );
AOI22xp5_ASAP7_75t_L g982 ( .A1(n_946), .A2(n_895), .B1(n_926), .B2(n_920), .Y(n_982) );
INVx2_ASAP7_75t_L g983 ( .A(n_939), .Y(n_983) );
INVx1_ASAP7_75t_SL g984 ( .A(n_949), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_961), .B(n_904), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g986 ( .A(n_942), .B(n_924), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_942), .B(n_898), .Y(n_987) );
INVx1_ASAP7_75t_SL g988 ( .A(n_963), .Y(n_988) );
INVx1_ASAP7_75t_SL g989 ( .A(n_971), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_950), .B(n_898), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_950), .B(n_935), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_965), .B(n_937), .Y(n_992) );
AND2x2_ASAP7_75t_L g993 ( .A(n_960), .B(n_873), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_959), .Y(n_994) );
OR2x2_ASAP7_75t_L g995 ( .A(n_958), .B(n_881), .Y(n_995) );
INVx2_ASAP7_75t_L g996 ( .A(n_947), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_964), .B(n_878), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_959), .Y(n_998) );
AND2x4_ASAP7_75t_L g999 ( .A(n_967), .B(n_886), .Y(n_999) );
INVxp67_ASAP7_75t_L g1000 ( .A(n_975), .Y(n_1000) );
INVx2_ASAP7_75t_SL g1001 ( .A(n_967), .Y(n_1001) );
INVx1_ASAP7_75t_L g1002 ( .A(n_944), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_964), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_952), .B(n_901), .Y(n_1004) );
INVx2_ASAP7_75t_L g1005 ( .A(n_955), .Y(n_1005) );
INVx2_ASAP7_75t_L g1006 ( .A(n_969), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_987), .Y(n_1007) );
NAND3xp33_ASAP7_75t_L g1008 ( .A(n_982), .B(n_951), .C(n_945), .Y(n_1008) );
BUFx2_ASAP7_75t_L g1009 ( .A(n_988), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_987), .Y(n_1010) );
INVx1_ASAP7_75t_L g1011 ( .A(n_986), .Y(n_1011) );
OAI211xp5_ASAP7_75t_L g1012 ( .A1(n_989), .A2(n_940), .B(n_943), .C(n_884), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_986), .Y(n_1013) );
OAI322xp33_ASAP7_75t_L g1014 ( .A1(n_1000), .A2(n_981), .A3(n_953), .B1(n_977), .B2(n_895), .C1(n_954), .C2(n_957), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_991), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_997), .B(n_954), .Y(n_1016) );
AOI22xp5_ASAP7_75t_L g1017 ( .A1(n_985), .A2(n_976), .B1(n_948), .B2(n_956), .Y(n_1017) );
OR2x2_ASAP7_75t_L g1018 ( .A(n_983), .B(n_973), .Y(n_1018) );
AOI21xp33_ASAP7_75t_SL g1019 ( .A1(n_1001), .A2(n_978), .B(n_972), .Y(n_1019) );
OAI21xp33_ASAP7_75t_L g1020 ( .A1(n_984), .A2(n_972), .B(n_962), .Y(n_1020) );
INVx2_ASAP7_75t_L g1021 ( .A(n_1006), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_991), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_1009), .B(n_993), .Y(n_1023) );
AOI221x1_ASAP7_75t_L g1024 ( .A1(n_1008), .A2(n_1002), .B1(n_990), .B2(n_992), .C(n_1003), .Y(n_1024) );
OAI21xp33_ASAP7_75t_L g1025 ( .A1(n_1020), .A2(n_997), .B(n_995), .Y(n_1025) );
AOI21xp5_ASAP7_75t_L g1026 ( .A1(n_1012), .A2(n_999), .B(n_919), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_1016), .Y(n_1027) );
OAI211xp5_ASAP7_75t_L g1028 ( .A1(n_1019), .A2(n_929), .B(n_992), .C(n_941), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_1015), .Y(n_1029) );
AOI221x1_ASAP7_75t_SL g1030 ( .A1(n_1007), .A2(n_994), .B1(n_998), .B2(n_996), .C(n_1005), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1022), .Y(n_1031) );
NOR3xp33_ASAP7_75t_L g1032 ( .A(n_1014), .B(n_810), .C(n_856), .Y(n_1032) );
A2O1A1Ixp33_ASAP7_75t_L g1033 ( .A1(n_1017), .A2(n_800), .B(n_929), .C(n_836), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1034 ( .A(n_1030), .B(n_1011), .Y(n_1034) );
NAND4xp25_ASAP7_75t_L g1035 ( .A(n_1033), .B(n_813), .C(n_793), .D(n_856), .Y(n_1035) );
NAND4xp25_ASAP7_75t_L g1036 ( .A(n_1032), .B(n_793), .C(n_813), .D(n_852), .Y(n_1036) );
AOI21xp5_ASAP7_75t_L g1037 ( .A1(n_1026), .A2(n_1010), .B(n_1013), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_1027), .B(n_1021), .Y(n_1038) );
A2O1A1Ixp33_ASAP7_75t_SL g1039 ( .A1(n_1028), .A2(n_852), .B(n_905), .C(n_831), .Y(n_1039) );
OAI211xp5_ASAP7_75t_L g1040 ( .A1(n_1025), .A2(n_846), .B(n_905), .C(n_1004), .Y(n_1040) );
NOR3xp33_ASAP7_75t_L g1041 ( .A(n_1040), .B(n_1029), .C(n_1031), .Y(n_1041) );
AOI22xp5_ASAP7_75t_L g1042 ( .A1(n_1037), .A2(n_1023), .B1(n_979), .B2(n_1018), .Y(n_1042) );
NOR2x1_ASAP7_75t_L g1043 ( .A(n_1035), .B(n_928), .Y(n_1043) );
OR2x2_ASAP7_75t_L g1044 ( .A(n_1038), .B(n_957), .Y(n_1044) );
NOR3x1_ASAP7_75t_L g1045 ( .A(n_1039), .B(n_1024), .C(n_921), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1034), .Y(n_1046) );
NOR2x1_ASAP7_75t_L g1047 ( .A(n_1043), .B(n_1036), .Y(n_1047) );
NAND5xp2_ASAP7_75t_L g1048 ( .A(n_1046), .B(n_927), .C(n_925), .D(n_828), .E(n_850), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1044), .Y(n_1049) );
INVx2_ASAP7_75t_L g1050 ( .A(n_1045), .Y(n_1050) );
O2A1O1Ixp5_ASAP7_75t_L g1051 ( .A1(n_1050), .A2(n_1041), .B(n_928), .C(n_827), .Y(n_1051) );
AOI22xp5_ASAP7_75t_L g1052 ( .A1(n_1047), .A2(n_1042), .B1(n_912), .B2(n_979), .Y(n_1052) );
NOR2xp67_ASAP7_75t_L g1053 ( .A(n_1049), .B(n_292), .Y(n_1053) );
AOI22xp5_ASAP7_75t_L g1054 ( .A1(n_1053), .A2(n_1048), .B1(n_913), .B2(n_853), .Y(n_1054) );
INVx2_ASAP7_75t_SL g1055 ( .A(n_1052), .Y(n_1055) );
XNOR2xp5_ASAP7_75t_L g1056 ( .A(n_1055), .B(n_1051), .Y(n_1056) );
OR2x2_ASAP7_75t_L g1057 ( .A(n_1054), .B(n_974), .Y(n_1057) );
OAI22x1_ASAP7_75t_L g1058 ( .A1(n_1056), .A2(n_934), .B1(n_870), .B2(n_915), .Y(n_1058) );
HB1xp67_ASAP7_75t_L g1059 ( .A(n_1057), .Y(n_1059) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1059), .Y(n_1060) );
OAI21x1_ASAP7_75t_SL g1061 ( .A1(n_1058), .A2(n_803), .B(n_938), .Y(n_1061) );
OA21x2_ASAP7_75t_L g1062 ( .A1(n_1060), .A2(n_932), .B(n_938), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_1061), .B(n_936), .Y(n_1063) );
AOI22xp5_ASAP7_75t_SL g1064 ( .A1(n_1063), .A2(n_966), .B1(n_909), .B2(n_968), .Y(n_1064) );
OAI22x1_ASAP7_75t_L g1065 ( .A1(n_1062), .A2(n_858), .B1(n_968), .B2(n_980), .Y(n_1065) );
OR2x6_ASAP7_75t_L g1066 ( .A(n_1065), .B(n_867), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_1066), .A2(n_1064), .B1(n_970), .B2(n_908), .Y(n_1067) );
endmodule