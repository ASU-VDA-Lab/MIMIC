module fake_jpeg_15920_n_316 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_316);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_316;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_0),
.C(n_1),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_17),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_32),
.A2(n_18),
.B1(n_15),
.B2(n_23),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_48),
.B1(n_51),
.B2(n_15),
.Y(n_65)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_14),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_30),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_32),
.A2(n_18),
.B1(n_24),
.B2(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_31),
.A2(n_18),
.B1(n_28),
.B2(n_22),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_31),
.A2(n_18),
.B1(n_28),
.B2(n_22),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_52),
.A2(n_35),
.B1(n_31),
.B2(n_15),
.Y(n_57)
);

NAND2xp33_ASAP7_75t_SL g54 ( 
.A(n_38),
.B(n_21),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_55),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_34),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_50),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_58),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_52),
.B(n_35),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_62),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_50),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_66),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_55),
.B(n_34),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_68),
.B(n_72),
.Y(n_90)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_73),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_35),
.B1(n_38),
.B2(n_33),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_53),
.B1(n_43),
.B2(n_41),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_22),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_39),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_28),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_76),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_23),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

AOI32xp33_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_45),
.A3(n_49),
.B1(n_40),
.B2(n_38),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_80),
.A2(n_84),
.B(n_97),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_76),
.B1(n_75),
.B2(n_72),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_83),
.A2(n_86),
.B1(n_88),
.B2(n_96),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_41),
.B1(n_42),
.B2(n_33),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_67),
.A2(n_57),
.B1(n_63),
.B2(n_42),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_SL g89 ( 
.A(n_68),
.B(n_48),
.C(n_51),
.Y(n_89)
);

NOR2xp67_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_21),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_65),
.B(n_55),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_62),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_67),
.A2(n_42),
.B1(n_41),
.B2(n_29),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_63),
.A2(n_41),
.B1(n_60),
.B2(n_29),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_71),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_103),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_59),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_56),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_107),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_61),
.C(n_73),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_92),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_112),
.B(n_127),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_53),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_114),
.A2(n_115),
.B1(n_128),
.B2(n_89),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_53),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_90),
.B(n_77),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_64),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_120),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_87),
.Y(n_120)
);

OR2x2_ASAP7_75t_SL g121 ( 
.A(n_90),
.B(n_24),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_116),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_79),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_43),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_83),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_141),
.B(n_114),
.Y(n_156)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_137),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_121),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_101),
.Y(n_136)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_153),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_93),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_150),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_80),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_106),
.C(n_109),
.Y(n_164)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_84),
.B1(n_88),
.B2(n_89),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_148),
.A2(n_114),
.B1(n_113),
.B2(n_115),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_83),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_101),
.Y(n_151)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_104),
.B(n_60),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_154),
.Y(n_170)
);

AND2x6_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_99),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_156),
.A2(n_178),
.B(n_179),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_157),
.B(n_177),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_161),
.A2(n_165),
.B1(n_168),
.B2(n_169),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_133),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_134),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_166),
.C(n_172),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_148),
.A2(n_126),
.B1(n_99),
.B2(n_114),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_119),
.C(n_115),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_118),
.B1(n_124),
.B2(n_112),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_167),
.A2(n_181),
.B1(n_140),
.B2(n_25),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_142),
.A2(n_97),
.B1(n_96),
.B2(n_85),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_145),
.A2(n_125),
.B1(n_111),
.B2(n_98),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_78),
.C(n_74),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_180),
.C(n_182),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_145),
.A2(n_101),
.B1(n_29),
.B2(n_30),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_174),
.A2(n_183),
.B1(n_37),
.B2(n_16),
.Y(n_205)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_175),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_132),
.Y(n_177)
);

OA21x2_ASAP7_75t_L g178 ( 
.A1(n_144),
.A2(n_107),
.B(n_36),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_129),
.B(n_149),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_78),
.C(n_74),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_16),
.B1(n_20),
.B2(n_25),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_36),
.C(n_29),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_141),
.A2(n_37),
.B1(n_36),
.B2(n_23),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_156),
.A2(n_131),
.B(n_129),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_187),
.A2(n_192),
.B(n_195),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_159),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_149),
.Y(n_189)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_152),
.Y(n_190)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_134),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_130),
.Y(n_193)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_193),
.Y(n_223)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

AOI22x1_ASAP7_75t_SL g195 ( 
.A1(n_161),
.A2(n_153),
.B1(n_137),
.B2(n_131),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_166),
.B(n_155),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_172),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_133),
.Y(n_198)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_198),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_155),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_206),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_140),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_200),
.B(n_209),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_147),
.C(n_139),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_204),
.C(n_183),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_202),
.A2(n_24),
.B1(n_25),
.B2(n_20),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_164),
.B(n_139),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_205),
.B(n_26),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_159),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_174),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_170),
.A2(n_0),
.B(n_1),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_208),
.A2(n_199),
.B(n_194),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_158),
.B(n_27),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_195),
.A2(n_163),
.B1(n_157),
.B2(n_158),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_214),
.A2(n_226),
.B1(n_228),
.B2(n_13),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_196),
.A2(n_165),
.B1(n_180),
.B2(n_168),
.Y(n_215)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_184),
.Y(n_236)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_0),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_160),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_222),
.C(n_224),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_182),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_186),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_27),
.C(n_19),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_225),
.B(n_26),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_192),
.A2(n_37),
.B1(n_1),
.B2(n_2),
.Y(n_228)
);

INVxp33_ASAP7_75t_SL g230 ( 
.A(n_188),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_230),
.A2(n_231),
.B(n_192),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_201),
.B(n_191),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_241),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_SL g235 ( 
.A1(n_217),
.A2(n_187),
.B(n_196),
.C(n_203),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_235),
.A2(n_243),
.B(n_231),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_238),
.C(n_239),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_188),
.Y(n_237)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_184),
.C(n_197),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_185),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_213),
.A2(n_208),
.B(n_207),
.Y(n_240)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_240),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_185),
.C(n_186),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_248),
.B(n_211),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_217),
.A2(n_205),
.B1(n_202),
.B2(n_16),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_246),
.B(n_250),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_213),
.A2(n_13),
.B(n_12),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_249),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_19),
.C(n_27),
.Y(n_249)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_255),
.A2(n_257),
.B(n_264),
.Y(n_268)
);

OAI321xp33_ASAP7_75t_L g257 ( 
.A1(n_243),
.A2(n_211),
.A3(n_219),
.B1(n_223),
.B2(n_228),
.C(n_229),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_210),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_260),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_239),
.B(n_212),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_248),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_262),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_241),
.B(n_215),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_216),
.Y(n_264)
);

BUFx24_ASAP7_75t_SL g265 ( 
.A(n_236),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_265),
.B(n_13),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_232),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_272),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_251),
.A2(n_235),
.B(n_232),
.Y(n_269)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_263),
.A2(n_235),
.B(n_249),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_270),
.A2(n_11),
.B(n_1),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_238),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_235),
.C(n_19),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_274),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_26),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_277),
.B(n_279),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_26),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_278),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_11),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_17),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_258),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_283),
.Y(n_300)
);

AO21x1_ASAP7_75t_L g284 ( 
.A1(n_275),
.A2(n_255),
.B(n_271),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_8),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_280),
.B(n_267),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_285),
.A2(n_3),
.B(n_7),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_256),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_291),
.Y(n_299)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_289),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_17),
.Y(n_291)
);

AOI322xp5_ASAP7_75t_L g292 ( 
.A1(n_274),
.A2(n_272),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_7),
.Y(n_298)
);

AOI211x1_ASAP7_75t_L g293 ( 
.A1(n_290),
.A2(n_0),
.B(n_3),
.C(n_4),
.Y(n_293)
);

OAI321xp33_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_298),
.A3(n_302),
.B1(n_288),
.B2(n_10),
.C(n_9),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_295),
.B(n_301),
.Y(n_306)
);

A2O1A1Ixp33_ASAP7_75t_L g296 ( 
.A1(n_286),
.A2(n_3),
.B(n_7),
.C(n_8),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_297),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_7),
.B(n_8),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_17),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_282),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_304),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_287),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_307),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_291),
.B(n_10),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_299),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_9),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_310),
.A2(n_10),
.B1(n_17),
.B2(n_311),
.Y(n_314)
);

AOI321xp33_ASAP7_75t_L g313 ( 
.A1(n_312),
.A2(n_306),
.A3(n_308),
.B1(n_9),
.B2(n_10),
.C(n_17),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_314),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_315),
.Y(n_316)
);


endmodule