module fake_jpeg_20473_n_345 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_28),
.Y(n_55)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_62),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_32),
.B1(n_35),
.B2(n_18),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_63),
.B1(n_37),
.B2(n_40),
.Y(n_72)
);

INVxp67_ASAP7_75t_SL g58 ( 
.A(n_38),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_31),
.B1(n_18),
.B2(n_20),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_29),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_47),
.A2(n_49),
.B1(n_32),
.B2(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_73),
.Y(n_113)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_47),
.C(n_43),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_80),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_72),
.A2(n_89),
.B1(n_90),
.B2(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

CKINVDCx6p67_ASAP7_75t_R g112 ( 
.A(n_75),
.Y(n_112)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_81),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_43),
.C(n_40),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_61),
.A2(n_26),
.B1(n_18),
.B2(n_31),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_82),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_85),
.B(n_96),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_92),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_62),
.A2(n_31),
.B1(n_19),
.B2(n_20),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_41),
.B1(n_40),
.B2(n_37),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_24),
.Y(n_91)
);

NAND3xp33_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_15),
.C(n_12),
.Y(n_103)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_67),
.A2(n_65),
.B1(n_66),
.B2(n_52),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_94),
.A2(n_21),
.B1(n_34),
.B2(n_36),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_60),
.A2(n_41),
.B1(n_37),
.B2(n_19),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_95),
.A2(n_97),
.B1(n_23),
.B2(n_27),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g96 ( 
.A(n_60),
.B(n_38),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_57),
.A2(n_41),
.B1(n_28),
.B2(n_27),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_100),
.Y(n_128)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_101),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_103),
.B(n_107),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_105),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_106),
.A2(n_121),
.B1(n_126),
.B2(n_25),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_21),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_71),
.A2(n_48),
.B1(n_45),
.B2(n_42),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_110),
.A2(n_120),
.B1(n_95),
.B2(n_84),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_48),
.B1(n_45),
.B2(n_42),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_117),
.A2(n_124),
.B1(n_70),
.B2(n_84),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_21),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_131),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_48),
.B1(n_45),
.B2(n_42),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_94),
.A2(n_36),
.B1(n_34),
.B2(n_21),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_96),
.A2(n_44),
.B1(n_33),
.B2(n_17),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_87),
.A2(n_21),
.B1(n_24),
.B2(n_15),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_83),
.A2(n_24),
.B(n_15),
.C(n_14),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_91),
.C(n_99),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_135),
.B(n_129),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_83),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_137),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_86),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_78),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_140),
.Y(n_188)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_44),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_77),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_141),
.B(n_146),
.Y(n_192)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_147),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_125),
.B(n_88),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_125),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_148),
.B(n_150),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_149),
.A2(n_153),
.B1(n_112),
.B2(n_132),
.Y(n_185)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_75),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_155),
.B(n_157),
.Y(n_166)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_156),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_123),
.B(n_110),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_104),
.B(n_10),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_158),
.B(n_104),
.Y(n_163)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_116),
.Y(n_159)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_160),
.B(n_161),
.Y(n_190)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_163),
.B(n_178),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_152),
.A2(n_115),
.B1(n_123),
.B2(n_118),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_164),
.A2(n_167),
.B1(n_187),
.B2(n_189),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_118),
.B(n_148),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_165),
.A2(n_175),
.B(n_182),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_152),
.A2(n_115),
.B1(n_120),
.B2(n_105),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_131),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_177),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_146),
.A2(n_112),
.B1(n_108),
.B2(n_132),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_173),
.A2(n_185),
.B1(n_191),
.B2(n_142),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_134),
.A2(n_133),
.B(n_130),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_130),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_136),
.B(n_129),
.Y(n_178)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_157),
.A2(n_102),
.B(n_108),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_186),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_184),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_144),
.A2(n_112),
.B1(n_114),
.B2(n_33),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_140),
.A2(n_112),
.B1(n_114),
.B2(n_74),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_153),
.A2(n_112),
.B1(n_109),
.B2(n_116),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_150),
.A2(n_109),
.B1(n_10),
.B2(n_11),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_193),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_195),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_190),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_198),
.Y(n_230)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_197),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_185),
.A2(n_139),
.B1(n_151),
.B2(n_155),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_168),
.B(n_138),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_200),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_141),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_209),
.Y(n_234)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_203),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_162),
.B(n_158),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_206),
.Y(n_243)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_172),
.A2(n_151),
.B1(n_161),
.B2(n_156),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_166),
.B(n_160),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_212),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_184),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_211),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_172),
.A2(n_151),
.B1(n_143),
.B2(n_147),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_159),
.Y(n_213)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_169),
.B(n_143),
.Y(n_214)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_214),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_162),
.B(n_109),
.Y(n_215)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_170),
.B(n_25),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_216),
.A2(n_221),
.B1(n_222),
.B2(n_0),
.Y(n_249)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_217),
.A2(n_218),
.B(n_223),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_192),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_25),
.C(n_33),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_177),
.C(n_186),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_165),
.A2(n_33),
.B1(n_17),
.B2(n_2),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_175),
.A2(n_17),
.B1(n_16),
.B2(n_14),
.Y(n_222)
);

AND2x2_ASAP7_75t_SL g223 ( 
.A(n_192),
.B(n_17),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_187),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_224),
.A2(n_182),
.B1(n_179),
.B2(n_164),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_225),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_219),
.A2(n_167),
.B1(n_188),
.B2(n_189),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_227),
.A2(n_198),
.B1(n_224),
.B2(n_226),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_231),
.C(n_220),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_171),
.C(n_188),
.Y(n_231)
);

AO22x2_ASAP7_75t_L g235 ( 
.A1(n_219),
.A2(n_179),
.B1(n_163),
.B2(n_176),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_240),
.Y(n_256)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_208),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_217),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_199),
.Y(n_237)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_204),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_202),
.A2(n_180),
.B(n_176),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_241),
.A2(n_202),
.B(n_214),
.Y(n_253)
);

OAI21xp33_ASAP7_75t_L g245 ( 
.A1(n_196),
.A2(n_16),
.B(n_13),
.Y(n_245)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_245),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_201),
.Y(n_258)
);

BUFx4f_ASAP7_75t_SL g251 ( 
.A(n_240),
.Y(n_251)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_252),
.A2(n_257),
.B1(n_265),
.B2(n_225),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_253),
.A2(n_254),
.B(n_235),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_230),
.A2(n_212),
.B(n_209),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_231),
.B(n_194),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_259),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_227),
.A2(n_205),
.B1(n_221),
.B2(n_218),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_258),
.A2(n_234),
.B1(n_248),
.B2(n_244),
.Y(n_272)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_243),
.B(n_204),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_261),
.B(n_270),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_230),
.B(n_205),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_254),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_247),
.A2(n_223),
.B1(n_210),
.B2(n_197),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_271),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_247),
.A2(n_207),
.B1(n_203),
.B2(n_216),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_269),
.A2(n_246),
.B1(n_248),
.B2(n_223),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_232),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_232),
.Y(n_271)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_272),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_228),
.C(n_241),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_283),
.C(n_288),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_258),
.A2(n_229),
.B1(n_234),
.B2(n_244),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_275),
.A2(n_277),
.B1(n_285),
.B2(n_235),
.Y(n_294)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_282),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_246),
.C(n_242),
.Y(n_283)
);

A2O1A1Ixp33_ASAP7_75t_L g284 ( 
.A1(n_256),
.A2(n_235),
.B(n_239),
.C(n_238),
.Y(n_284)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_284),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_267),
.A2(n_256),
.B1(n_268),
.B2(n_257),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_289),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_268),
.A2(n_235),
.B1(n_239),
.B2(n_238),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_287),
.A2(n_289),
.B1(n_273),
.B2(n_282),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_233),
.C(n_193),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_253),
.B(n_233),
.C(n_250),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_265),
.C(n_269),
.Y(n_292)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_292),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_252),
.C(n_251),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_297),
.C(n_279),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_301),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_280),
.A2(n_251),
.B1(n_260),
.B2(n_263),
.Y(n_295)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_295),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_208),
.C(n_263),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_290),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_303),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_236),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_283),
.B(n_13),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_281),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_305),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_276),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_277),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_293),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_308),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_291),
.A2(n_281),
.B(n_278),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_309),
.A2(n_292),
.B1(n_298),
.B2(n_302),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_296),
.A2(n_284),
.B(n_287),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_310),
.A2(n_9),
.B1(n_1),
.B2(n_2),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_314),
.C(n_316),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_12),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_12),
.C(n_11),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_313),
.B(n_291),
.Y(n_319)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_319),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_321),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_315),
.A2(n_299),
.B1(n_296),
.B2(n_9),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_326),
.C(n_316),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_307),
.A2(n_0),
.B(n_1),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_324),
.A2(n_327),
.B(n_4),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_0),
.C(n_1),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_314),
.B(n_3),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_317),
.Y(n_328)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_328),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_330),
.B(n_332),
.Y(n_336)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_325),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_333),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_311),
.C(n_308),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_329),
.B(n_332),
.Y(n_338)
);

AO21x1_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_336),
.B(n_334),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_335),
.C(n_331),
.Y(n_340)
);

AOI322xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_328),
.A3(n_320),
.B1(n_326),
.B2(n_318),
.C1(n_7),
.C2(n_6),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_4),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_342),
.A2(n_4),
.B(n_5),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_4),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_5),
.Y(n_345)
);


endmodule