module fake_jpeg_27447_n_308 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_30),
.C(n_25),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_46),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_16),
.Y(n_46)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_32),
.B1(n_26),
.B2(n_22),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_56),
.B1(n_38),
.B2(n_35),
.Y(n_70)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx2_ASAP7_75t_SL g78 ( 
.A(n_53),
.Y(n_78)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_35),
.A2(n_32),
.B1(n_38),
.B2(n_34),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_32),
.B1(n_22),
.B2(n_26),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_38),
.B1(n_35),
.B2(n_34),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_56),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_62),
.Y(n_106)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_48),
.A2(n_32),
.B1(n_39),
.B2(n_22),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_65),
.A2(n_74),
.B1(n_53),
.B2(n_50),
.Y(n_110)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_72),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_70),
.A2(n_77),
.B1(n_86),
.B2(n_57),
.Y(n_113)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_71),
.A2(n_75),
.B(n_76),
.Y(n_112)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_34),
.B1(n_33),
.B2(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_20),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_20),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_20),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_84),
.Y(n_107)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_40),
.Y(n_84)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_59),
.A2(n_16),
.B1(n_27),
.B2(n_31),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_52),
.Y(n_87)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_17),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_88),
.B(n_111),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_92),
.B(n_101),
.Y(n_136)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_93),
.Y(n_126)
);

AO22x1_ASAP7_75t_SL g94 ( 
.A1(n_79),
.A2(n_57),
.B1(n_33),
.B2(n_40),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_94),
.A2(n_110),
.B1(n_80),
.B2(n_87),
.Y(n_123)
);

FAx1_ASAP7_75t_SL g95 ( 
.A(n_68),
.B(n_82),
.CI(n_84),
.CON(n_95),
.SN(n_95)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_102),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_0),
.B(n_1),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_97),
.A2(n_0),
.B(n_1),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_33),
.C(n_37),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_37),
.C(n_49),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_71),
.B(n_29),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_104),
.B(n_23),
.Y(n_135)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_114),
.Y(n_117)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_69),
.A2(n_29),
.B1(n_28),
.B2(n_17),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_SL g124 ( 
.A1(n_111),
.A2(n_113),
.B(n_17),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_66),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_114),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_91),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_116),
.B(n_121),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_125),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_119),
.B(n_141),
.Y(n_160)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_122),
.B(n_133),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_124),
.B1(n_139),
.B2(n_102),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_98),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_98),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_138),
.Y(n_147)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_130),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_66),
.C(n_76),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_105),
.C(n_33),
.Y(n_152)
);

OR2x2_ASAP7_75t_SL g132 ( 
.A(n_95),
.B(n_28),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_132),
.A2(n_137),
.B(n_140),
.Y(n_163)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_135),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_75),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_101),
.A2(n_106),
.B1(n_97),
.B2(n_110),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_72),
.B(n_63),
.C(n_83),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_103),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_143),
.B(n_152),
.Y(n_196)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_149),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_118),
.B(n_136),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_145),
.A2(n_154),
.B(n_165),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_148),
.A2(n_158),
.B1(n_167),
.B2(n_170),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_100),
.B(n_1),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_100),
.B1(n_99),
.B2(n_93),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_156),
.A2(n_121),
.B1(n_115),
.B2(n_129),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_96),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_159),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_137),
.A2(n_90),
.B1(n_99),
.B2(n_109),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_109),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_73),
.Y(n_161)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

AO21x2_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_44),
.B(n_73),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_162),
.A2(n_165),
.B1(n_150),
.B2(n_168),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_37),
.Y(n_166)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_59),
.B1(n_31),
.B2(n_16),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_126),
.Y(n_168)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_168),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_0),
.B(n_1),
.Y(n_169)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_134),
.A2(n_31),
.B1(n_23),
.B2(n_27),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_161),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_172),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_173),
.A2(n_176),
.B1(n_182),
.B2(n_164),
.Y(n_208)
);

OAI211xp5_ASAP7_75t_L g175 ( 
.A1(n_162),
.A2(n_27),
.B(n_23),
.C(n_130),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_178),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_162),
.A2(n_134),
.B1(n_126),
.B2(n_120),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_177),
.A2(n_183),
.B1(n_164),
.B2(n_166),
.Y(n_215)
);

BUFx24_ASAP7_75t_SL g178 ( 
.A(n_151),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_115),
.B1(n_21),
.B2(n_18),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_162),
.A2(n_21),
.B1(n_18),
.B2(n_30),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_194),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_146),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_187),
.B(n_189),
.Y(n_217)
);

AOI32xp33_ASAP7_75t_L g189 ( 
.A1(n_149),
.A2(n_19),
.A3(n_25),
.B1(n_4),
.B2(n_5),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_153),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_190),
.B(n_197),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_148),
.A2(n_154),
.B1(n_156),
.B2(n_169),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_192),
.A2(n_21),
.B1(n_18),
.B2(n_25),
.Y(n_220)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_142),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_153),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_188),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_199),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_143),
.C(n_160),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_200),
.B(n_25),
.C(n_19),
.Y(n_240)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_142),
.Y(n_203)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_205),
.Y(n_223)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_182),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_209),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_208),
.A2(n_220),
.B1(n_198),
.B2(n_179),
.Y(n_235)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_160),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_186),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_211),
.A2(n_212),
.B(n_185),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_179),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_191),
.A2(n_163),
.B(n_147),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_213),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_191),
.Y(n_214)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_215),
.A2(n_219),
.B1(n_174),
.B2(n_180),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_147),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_216),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_145),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_218),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_184),
.A2(n_166),
.B1(n_152),
.B2(n_163),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_230),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_174),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_229),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_180),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_198),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_238),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_213),
.B(n_183),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_240),
.Y(n_256)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_235),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_185),
.Y(n_238)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_239),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_19),
.C(n_9),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_201),
.C(n_199),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_221),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_216),
.Y(n_269)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_245),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_240),
.C(n_227),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_249),
.C(n_232),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_212),
.C(n_209),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_255),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_206),
.Y(n_252)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_242),
.Y(n_253)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_222),
.Y(n_254)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_254),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_222),
.Y(n_255)
);

NOR2xp67_ASAP7_75t_R g258 ( 
.A(n_226),
.B(n_217),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_258),
.A2(n_203),
.B1(n_211),
.B2(n_208),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_248),
.A2(n_234),
.B(n_237),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_263),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_269),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_223),
.C(n_204),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_9),
.C(n_5),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_225),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_11),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_243),
.A2(n_205),
.B1(n_228),
.B2(n_215),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_249),
.A2(n_202),
.B(n_236),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_270),
.A2(n_257),
.B(n_247),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_271),
.Y(n_275)
);

OAI321xp33_ASAP7_75t_L g272 ( 
.A1(n_263),
.A2(n_245),
.A3(n_256),
.B1(n_247),
.B2(n_244),
.C(n_251),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_282),
.Y(n_284)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_260),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_276),
.A2(n_281),
.B1(n_270),
.B2(n_265),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_13),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_9),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_280),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_10),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_262),
.A2(n_11),
.B(n_7),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_283),
.A2(n_261),
.B(n_259),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_277),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_276),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_290),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_288),
.A2(n_289),
.B1(n_285),
.B2(n_286),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_266),
.Y(n_290)
);

AO21x1_ASAP7_75t_L g292 ( 
.A1(n_275),
.A2(n_267),
.B(n_268),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_292),
.B(n_282),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_293),
.A2(n_294),
.B(n_296),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_291),
.A2(n_273),
.B(n_279),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_298),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_8),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_10),
.C(n_11),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_299),
.A2(n_10),
.B(n_12),
.Y(n_302)
);

OAI21x1_ASAP7_75t_L g303 ( 
.A1(n_302),
.A2(n_297),
.B(n_295),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_301),
.C(n_300),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_12),
.C(n_13),
.Y(n_305)
);

OAI21x1_ASAP7_75t_SL g306 ( 
.A1(n_305),
.A2(n_15),
.B(n_3),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_15),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_307),
.B(n_15),
.Y(n_308)
);


endmodule