module real_jpeg_29824_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_0),
.A2(n_46),
.B1(n_47),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_52),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_0),
.A2(n_52),
.B1(n_62),
.B2(n_63),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_0),
.A2(n_34),
.B1(n_35),
.B2(n_52),
.Y(n_153)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_1),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_1),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_1),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_1),
.A2(n_127),
.B(n_185),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_2),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_2),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_64),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_64),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_64),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_3),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_3),
.B(n_46),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g212 ( 
.A1(n_3),
.A2(n_46),
.B(n_208),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_168),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_3),
.A2(n_11),
.B(n_34),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_3),
.B(n_134),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_3),
.A2(n_85),
.B1(n_86),
.B2(n_256),
.Y(n_258)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_7),
.A2(n_62),
.B1(n_63),
.B2(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_7),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_7),
.A2(n_46),
.B1(n_47),
.B2(n_138),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_138),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_138),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_8),
.A2(n_46),
.B1(n_47),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_8),
.A2(n_55),
.B1(n_62),
.B2(n_63),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_55),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_55),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_9),
.A2(n_38),
.B1(n_62),
.B2(n_63),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_9),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_10),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_10),
.A2(n_62),
.B1(n_63),
.B2(n_164),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_164),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_164),
.Y(n_248)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_12),
.A2(n_62),
.B1(n_63),
.B2(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_12),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_12),
.A2(n_46),
.B1(n_47),
.B2(n_170),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_170),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_170),
.Y(n_256)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_49),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_15),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_114),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_113),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_97),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_20),
.B(n_97),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_72),
.C(n_82),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_21),
.A2(n_22),
.B1(n_72),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_56),
.B1(n_70),
.B2(n_71),
.Y(n_22)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_24),
.A2(n_25),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_24),
.B(n_40),
.C(n_56),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_33),
.B(n_36),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_26),
.A2(n_92),
.B(n_93),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_26),
.A2(n_33),
.B1(n_92),
.B2(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_26),
.A2(n_36),
.B(n_93),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_26),
.A2(n_33),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_26),
.A2(n_77),
.B(n_216),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_26),
.A2(n_33),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_26),
.A2(n_33),
.B1(n_215),
.B2(n_233),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_33),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g207 ( 
.A1(n_28),
.A2(n_47),
.A3(n_49),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g209 ( 
.A(n_29),
.B(n_44),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_29),
.A2(n_32),
.B(n_168),
.C(n_235),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_33),
.A2(n_79),
.B(n_132),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_33),
.B(n_168),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_34),
.B(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_35),
.B(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_37),
.B(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_50),
.B(n_53),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_41),
.A2(n_107),
.B(n_179),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_41),
.A2(n_53),
.B(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_48),
.B1(n_51),
.B2(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_42),
.B(n_54),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_42),
.A2(n_48),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_42),
.A2(n_48),
.B1(n_163),
.B2(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_42),
.A2(n_48),
.B1(n_194),
.B2(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_48),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_43)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_47),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_46),
.B(n_59),
.Y(n_182)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_47),
.A2(n_67),
.B1(n_167),
.B2(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_48),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_48),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_56),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_56),
.A2(n_71),
.B1(n_99),
.B2(n_111),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_61),
.B(n_65),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_69),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_57),
.A2(n_61),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_57),
.A2(n_101),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_57),
.B(n_168),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_57),
.A2(n_101),
.B1(n_137),
.B2(n_176),
.Y(n_291)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_59),
.B(n_63),
.C(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_58),
.B(n_95),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_58),
.A2(n_66),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_63),
.Y(n_67)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

HAxp5_ASAP7_75t_SL g167 ( 
.A(n_63),
.B(n_168),
.CON(n_167),
.SN(n_167)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_66),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_72),
.A2(n_73),
.B(n_76),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_72),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_75),
.A2(n_109),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_78),
.B(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_82),
.A2(n_83),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_90),
.B(n_94),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_84),
.A2(n_94),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_84),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_84),
.A2(n_91),
.B1(n_120),
.B2(n_308),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_87),
.B(n_88),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_85),
.A2(n_153),
.B(n_154),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_85),
.A2(n_87),
.B1(n_153),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_85),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_85),
.A2(n_129),
.B(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_85),
.A2(n_87),
.B1(n_248),
.B2(n_256),
.Y(n_255)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_86),
.B(n_168),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_130),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_89),
.A2(n_155),
.B(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_91),
.Y(n_308)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_112),
.Y(n_97)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_103),
.B1(n_104),
.B2(n_110),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_100),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_101),
.A2(n_137),
.B(n_139),
.Y(n_136)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_108),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_144),
.B(n_317),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_140),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_116),
.B(n_140),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.C(n_122),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_117),
.B(n_121),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_122),
.A2(n_123),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_133),
.C(n_135),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_124),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_131),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_125),
.B(n_131),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_130),
.A2(n_206),
.B1(n_247),
.B2(n_249),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_133),
.A2(n_135),
.B1(n_136),
.B2(n_305),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_133),
.Y(n_305)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_311),
.B(n_316),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_298),
.B(n_310),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_198),
.B(n_279),
.C(n_297),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_186),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_148),
.B(n_186),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_171),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_158),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_150),
.B(n_158),
.C(n_171),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_151),
.B(n_152),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.C(n_166),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_166),
.B(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_169),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_180),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_177),
.B2(n_178),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_173),
.B(n_178),
.C(n_180),
.Y(n_295)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_183),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.C(n_192),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_187),
.A2(n_188),
.B1(n_274),
.B2(n_276),
.Y(n_273)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_275),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_192),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.C(n_196),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_193),
.B(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_221),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_195),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_278),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_271),
.B(n_277),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_226),
.B(n_270),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_217),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_202),
.B(n_217),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_210),
.C(n_213),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_203),
.A2(n_204),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_207),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_222),
.B2(n_223),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_218),
.B(n_224),
.C(n_225),
.Y(n_272)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_264),
.B(n_269),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_244),
.B(n_263),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_236),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_229),
.B(n_236),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_234),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_230),
.A2(n_231),
.B1(n_234),
.B2(n_251),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_234),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_242),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_241),
.C(n_242),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_243),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_252),
.B(n_262),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_250),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_246),
.B(n_250),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_257),
.B(n_261),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_254),
.B(n_255),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_265),
.B(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_272),
.B(n_273),
.Y(n_277)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_274),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_280),
.B(n_281),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_295),
.B2(n_296),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_287),
.C(n_296),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_290),
.C(n_293),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_295),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_299),
.B(n_300),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_309),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_306),
.B2(n_307),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_307),
.C(n_309),
.Y(n_312)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_312),
.B(n_313),
.Y(n_316)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);


endmodule