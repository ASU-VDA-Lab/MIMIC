module fake_jpeg_20630_n_10 (n_3, n_2, n_1, n_0, n_4, n_10);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_10;

wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

OAI22xp5_ASAP7_75t_SL g5 ( 
.A1(n_2),
.A2(n_4),
.B1(n_3),
.B2(n_0),
.Y(n_5)
);

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_1),
.Y(n_6)
);

OAI21xp5_ASAP7_75t_L g7 ( 
.A1(n_3),
.A2(n_2),
.B(n_0),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_1),
.B(n_0),
.Y(n_8)
);

AOI22xp5_ASAP7_75t_L g9 ( 
.A1(n_5),
.A2(n_4),
.B1(n_8),
.B2(n_7),
.Y(n_9)
);

A2O1A1Ixp33_ASAP7_75t_SL g10 ( 
.A1(n_9),
.A2(n_5),
.B(n_7),
.C(n_6),
.Y(n_10)
);


endmodule