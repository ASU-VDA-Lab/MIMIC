module real_aes_8480_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_505;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_0), .B(n_85), .C(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g120 ( .A(n_0), .Y(n_120) );
INVx1_ASAP7_75t_L g534 ( .A(n_1), .Y(n_534) );
INVx1_ASAP7_75t_L g154 ( .A(n_2), .Y(n_154) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_3), .A2(n_38), .B1(n_179), .B2(n_480), .Y(n_503) );
AOI21xp33_ASAP7_75t_L g186 ( .A1(n_4), .A2(n_170), .B(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_5), .B(n_168), .Y(n_546) );
AND2x6_ASAP7_75t_L g147 ( .A(n_6), .B(n_148), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_7), .A2(n_257), .B(n_258), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_8), .B(n_108), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_8), .B(n_39), .Y(n_121) );
INVx1_ASAP7_75t_L g192 ( .A(n_9), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_10), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g139 ( .A(n_11), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_12), .B(n_160), .Y(n_489) );
INVx1_ASAP7_75t_L g263 ( .A(n_13), .Y(n_263) );
INVx1_ASAP7_75t_L g528 ( .A(n_14), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_15), .B(n_135), .Y(n_517) );
AO32x2_ASAP7_75t_L g501 ( .A1(n_16), .A2(n_134), .A3(n_168), .B1(n_482), .B2(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_17), .B(n_179), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_18), .B(n_175), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_19), .B(n_135), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_20), .A2(n_49), .B1(n_179), .B2(n_480), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_21), .B(n_170), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_22), .A2(n_98), .B1(n_736), .B2(n_737), .Y(n_735) );
INVx1_ASAP7_75t_L g737 ( .A(n_22), .Y(n_737) );
AOI22xp33_ASAP7_75t_SL g481 ( .A1(n_23), .A2(n_76), .B1(n_160), .B2(n_179), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_24), .B(n_179), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_25), .B(n_182), .Y(n_181) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_26), .A2(n_261), .B(n_262), .C(n_264), .Y(n_260) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_27), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_28), .B(n_165), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_29), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_30), .B(n_115), .Y(n_441) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_31), .A2(n_88), .B1(n_125), .B2(n_126), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_31), .Y(n_125) );
INVx1_ASAP7_75t_L g207 ( .A(n_32), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_33), .B(n_165), .Y(n_473) );
INVx2_ASAP7_75t_L g145 ( .A(n_34), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_35), .B(n_179), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_36), .B(n_165), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_37), .A2(n_147), .B(n_150), .C(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g108 ( .A(n_39), .Y(n_108) );
INVx1_ASAP7_75t_L g205 ( .A(n_40), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_41), .B(n_158), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_42), .B(n_179), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_43), .A2(n_86), .B1(n_227), .B2(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_44), .B(n_179), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_45), .B(n_179), .Y(n_529) );
CKINVDCx16_ASAP7_75t_R g208 ( .A(n_46), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_47), .B(n_533), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_48), .B(n_170), .Y(n_251) );
AOI22xp33_ASAP7_75t_SL g521 ( .A1(n_50), .A2(n_61), .B1(n_160), .B2(n_179), .Y(n_521) );
OAI22xp5_ASAP7_75t_SL g733 ( .A1(n_51), .A2(n_734), .B1(n_735), .B2(n_738), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_51), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_52), .A2(n_150), .B1(n_160), .B2(n_203), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_53), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_54), .B(n_179), .Y(n_488) );
CKINVDCx16_ASAP7_75t_R g141 ( .A(n_55), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_56), .B(n_179), .Y(n_554) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_57), .A2(n_178), .B(n_190), .C(n_191), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_58), .A2(n_104), .B1(n_113), .B2(n_744), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_59), .Y(n_240) );
INVx1_ASAP7_75t_L g188 ( .A(n_60), .Y(n_188) );
INVx1_ASAP7_75t_L g148 ( .A(n_62), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_63), .B(n_179), .Y(n_535) );
INVx1_ASAP7_75t_L g138 ( .A(n_64), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_65), .Y(n_444) );
AO32x2_ASAP7_75t_L g477 ( .A1(n_66), .A2(n_168), .A3(n_243), .B1(n_478), .B2(n_482), .Y(n_477) );
INVx1_ASAP7_75t_L g553 ( .A(n_67), .Y(n_553) );
INVx1_ASAP7_75t_L g468 ( .A(n_68), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g122 ( .A1(n_69), .A2(n_123), .B1(n_439), .B2(n_440), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_69), .Y(n_439) );
A2O1A1Ixp33_ASAP7_75t_SL g174 ( .A1(n_70), .A2(n_175), .B(n_176), .C(n_178), .Y(n_174) );
INVxp67_ASAP7_75t_L g177 ( .A(n_71), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_72), .B(n_160), .Y(n_469) );
INVx1_ASAP7_75t_L g112 ( .A(n_73), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_74), .Y(n_210) );
INVx1_ASAP7_75t_L g233 ( .A(n_75), .Y(n_233) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_77), .A2(n_147), .B(n_150), .C(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_78), .B(n_480), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_79), .B(n_160), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_80), .B(n_155), .Y(n_223) );
INVx2_ASAP7_75t_L g136 ( .A(n_81), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_82), .B(n_175), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_83), .B(n_160), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g149 ( .A1(n_84), .A2(n_147), .B(n_150), .C(n_153), .Y(n_149) );
OR2x2_ASAP7_75t_L g117 ( .A(n_85), .B(n_118), .Y(n_117) );
OR2x2_ASAP7_75t_L g450 ( .A(n_85), .B(n_119), .Y(n_450) );
INVx2_ASAP7_75t_L g455 ( .A(n_85), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_87), .A2(n_102), .B1(n_160), .B2(n_161), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_88), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_89), .B(n_165), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_90), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_91), .A2(n_147), .B(n_150), .C(n_246), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g253 ( .A(n_92), .Y(n_253) );
INVx1_ASAP7_75t_L g173 ( .A(n_93), .Y(n_173) );
CKINVDCx16_ASAP7_75t_R g259 ( .A(n_94), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_95), .B(n_155), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_96), .B(n_160), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_97), .B(n_168), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_98), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_99), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_100), .A2(n_170), .B(n_171), .Y(n_169) );
AOI222xp33_ASAP7_75t_L g446 ( .A1(n_101), .A2(n_447), .B1(n_732), .B2(n_733), .C1(n_739), .C2(n_742), .Y(n_446) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx6p67_ASAP7_75t_R g745 ( .A(n_106), .Y(n_745) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AO21x1_ASAP7_75t_SL g113 ( .A1(n_114), .A2(n_442), .B(n_445), .Y(n_113) );
OAI21xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_122), .B(n_441), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NOR2x2_ASAP7_75t_L g741 ( .A(n_118), .B(n_455), .Y(n_741) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OR2x2_ASAP7_75t_L g454 ( .A(n_119), .B(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
INVx1_ASAP7_75t_L g440 ( .A(n_123), .Y(n_440) );
XNOR2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_127), .Y(n_123) );
INVx1_ASAP7_75t_L g451 ( .A(n_127), .Y(n_451) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_127), .A2(n_452), .B1(n_457), .B2(n_743), .Y(n_742) );
NAND2x1_ASAP7_75t_L g127 ( .A(n_128), .B(n_355), .Y(n_127) );
NOR5xp2_ASAP7_75t_L g128 ( .A(n_129), .B(n_278), .C(n_310), .D(n_325), .E(n_342), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_194), .B(n_215), .C(n_266), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_166), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_131), .B(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_131), .B(n_330), .Y(n_393) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_132), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_132), .B(n_212), .Y(n_279) );
AND2x2_ASAP7_75t_L g320 ( .A(n_132), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_132), .B(n_289), .Y(n_324) );
OR2x2_ASAP7_75t_L g361 ( .A(n_132), .B(n_200), .Y(n_361) );
INVx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g199 ( .A(n_133), .B(n_200), .Y(n_199) );
INVx3_ASAP7_75t_L g269 ( .A(n_133), .Y(n_269) );
OR2x2_ASAP7_75t_L g432 ( .A(n_133), .B(n_272), .Y(n_432) );
AO21x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_140), .B(n_162), .Y(n_133) );
AO21x2_ASAP7_75t_L g200 ( .A1(n_134), .A2(n_201), .B(n_209), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_134), .B(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g228 ( .A(n_134), .Y(n_228) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_135), .Y(n_168) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x2_ASAP7_75t_SL g165 ( .A(n_136), .B(n_137), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
OAI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_142), .B(n_149), .Y(n_140) );
OAI22xp33_ASAP7_75t_L g201 ( .A1(n_142), .A2(n_180), .B1(n_202), .B2(n_208), .Y(n_201) );
OAI21xp5_ASAP7_75t_L g232 ( .A1(n_142), .A2(n_233), .B(n_234), .Y(n_232) );
NAND2x1p5_ASAP7_75t_L g142 ( .A(n_143), .B(n_147), .Y(n_142) );
AND2x4_ASAP7_75t_L g170 ( .A(n_143), .B(n_147), .Y(n_170) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_146), .Y(n_143) );
INVx1_ASAP7_75t_L g533 ( .A(n_144), .Y(n_533) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g151 ( .A(n_145), .Y(n_151) );
INVx1_ASAP7_75t_L g161 ( .A(n_145), .Y(n_161) );
INVx1_ASAP7_75t_L g152 ( .A(n_146), .Y(n_152) );
INVx3_ASAP7_75t_L g156 ( .A(n_146), .Y(n_156) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_146), .Y(n_158) );
INVx1_ASAP7_75t_L g175 ( .A(n_146), .Y(n_175) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_146), .Y(n_204) );
INVx4_ASAP7_75t_SL g180 ( .A(n_147), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_147), .A2(n_467), .B(n_470), .Y(n_466) );
BUFx3_ASAP7_75t_L g482 ( .A(n_147), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g486 ( .A1(n_147), .A2(n_487), .B(n_491), .Y(n_486) );
OAI21xp5_ASAP7_75t_L g526 ( .A1(n_147), .A2(n_527), .B(n_531), .Y(n_526) );
OAI21xp5_ASAP7_75t_L g539 ( .A1(n_147), .A2(n_540), .B(n_543), .Y(n_539) );
INVx5_ASAP7_75t_L g172 ( .A(n_150), .Y(n_172) );
AND2x6_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_151), .Y(n_179) );
BUFx3_ASAP7_75t_L g227 ( .A(n_151), .Y(n_227) );
INVx1_ASAP7_75t_L g480 ( .A(n_151), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_157), .C(n_159), .Y(n_153) );
O2A1O1Ixp5_ASAP7_75t_SL g467 ( .A1(n_155), .A2(n_178), .B(n_468), .C(n_469), .Y(n_467) );
INVx2_ASAP7_75t_L g504 ( .A(n_155), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_155), .A2(n_541), .B(n_542), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_155), .A2(n_550), .B(n_551), .Y(n_549) );
INVx5_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_156), .B(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_156), .B(n_192), .Y(n_191) );
OAI22xp5_ASAP7_75t_SL g478 ( .A1(n_156), .A2(n_158), .B1(n_479), .B2(n_481), .Y(n_478) );
INVx2_ASAP7_75t_L g190 ( .A(n_158), .Y(n_190) );
INVx4_ASAP7_75t_L g249 ( .A(n_158), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_158), .A2(n_503), .B1(n_504), .B2(n_505), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_158), .A2(n_504), .B1(n_520), .B2(n_521), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_159), .A2(n_528), .B(n_529), .C(n_530), .Y(n_527) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_164), .B(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_164), .B(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g243 ( .A(n_165), .Y(n_243) );
OA21x2_ASAP7_75t_L g255 ( .A1(n_165), .A2(n_256), .B(n_265), .Y(n_255) );
OA21x2_ASAP7_75t_L g465 ( .A1(n_165), .A2(n_466), .B(n_473), .Y(n_465) );
OA21x2_ASAP7_75t_L g485 ( .A1(n_165), .A2(n_486), .B(n_494), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g334 ( .A1(n_166), .A2(n_335), .B1(n_336), .B2(n_339), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_166), .B(n_269), .Y(n_418) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_184), .Y(n_166) );
AND2x2_ASAP7_75t_L g214 ( .A(n_167), .B(n_200), .Y(n_214) );
AND2x2_ASAP7_75t_L g271 ( .A(n_167), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g276 ( .A(n_167), .Y(n_276) );
INVx3_ASAP7_75t_L g289 ( .A(n_167), .Y(n_289) );
OR2x2_ASAP7_75t_L g309 ( .A(n_167), .B(n_272), .Y(n_309) );
AND2x2_ASAP7_75t_L g328 ( .A(n_167), .B(n_185), .Y(n_328) );
BUFx2_ASAP7_75t_L g360 ( .A(n_167), .Y(n_360) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_181), .Y(n_167) );
INVx4_ASAP7_75t_L g183 ( .A(n_168), .Y(n_183) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_168), .A2(n_539), .B(n_546), .Y(n_538) );
BUFx2_ASAP7_75t_L g257 ( .A(n_170), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_174), .C(n_180), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_L g187 ( .A1(n_172), .A2(n_180), .B(n_188), .C(n_189), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g258 ( .A1(n_172), .A2(n_180), .B(n_259), .C(n_260), .Y(n_258) );
INVx1_ASAP7_75t_L g490 ( .A(n_175), .Y(n_490) );
INVx3_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_179), .Y(n_250) );
OA21x2_ASAP7_75t_L g185 ( .A1(n_182), .A2(n_186), .B(n_193), .Y(n_185) );
INVx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_SL g229 ( .A(n_183), .B(n_230), .Y(n_229) );
NAND3xp33_ASAP7_75t_L g518 ( .A(n_183), .B(n_482), .C(n_519), .Y(n_518) );
AO21x1_ASAP7_75t_L g608 ( .A1(n_183), .A2(n_519), .B(n_609), .Y(n_608) );
AND2x4_ASAP7_75t_L g275 ( .A(n_184), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_SL g184 ( .A(n_185), .Y(n_184) );
BUFx2_ASAP7_75t_L g198 ( .A(n_185), .Y(n_198) );
INVx2_ASAP7_75t_L g213 ( .A(n_185), .Y(n_213) );
OR2x2_ASAP7_75t_L g291 ( .A(n_185), .B(n_272), .Y(n_291) );
AND2x2_ASAP7_75t_L g321 ( .A(n_185), .B(n_200), .Y(n_321) );
AND2x2_ASAP7_75t_L g338 ( .A(n_185), .B(n_269), .Y(n_338) );
AND2x2_ASAP7_75t_L g378 ( .A(n_185), .B(n_289), .Y(n_378) );
AND2x2_ASAP7_75t_SL g414 ( .A(n_185), .B(n_214), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_190), .A2(n_492), .B(n_493), .Y(n_491) );
O2A1O1Ixp5_ASAP7_75t_L g552 ( .A1(n_190), .A2(n_532), .B(n_553), .C(n_554), .Y(n_552) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2xp33_ASAP7_75t_SL g195 ( .A(n_196), .B(n_211), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_197), .B(n_199), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_197), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_SL g197 ( .A(n_198), .Y(n_197) );
OAI21xp33_ASAP7_75t_L g352 ( .A1(n_198), .A2(n_214), .B(n_353), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_198), .B(n_200), .Y(n_408) );
AND2x2_ASAP7_75t_L g344 ( .A(n_199), .B(n_345), .Y(n_344) );
INVx3_ASAP7_75t_L g272 ( .A(n_200), .Y(n_272) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_200), .Y(n_370) );
OAI22xp5_ASAP7_75t_SL g203 ( .A1(n_204), .A2(n_205), .B1(n_206), .B2(n_207), .Y(n_203) );
INVx2_ASAP7_75t_L g206 ( .A(n_204), .Y(n_206) );
INVx4_ASAP7_75t_L g261 ( .A(n_204), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_211), .B(n_269), .Y(n_437) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_212), .A2(n_380), .B1(n_381), .B2(n_386), .Y(n_379) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
AND2x2_ASAP7_75t_L g270 ( .A(n_213), .B(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g308 ( .A(n_213), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_SL g345 ( .A(n_213), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_214), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g399 ( .A(n_214), .Y(n_399) );
CKINVDCx16_ASAP7_75t_R g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_241), .Y(n_216) );
INVx4_ASAP7_75t_L g285 ( .A(n_217), .Y(n_285) );
AND2x2_ASAP7_75t_L g363 ( .A(n_217), .B(n_330), .Y(n_363) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_231), .Y(n_217) );
INVx3_ASAP7_75t_L g282 ( .A(n_218), .Y(n_282) );
AND2x2_ASAP7_75t_L g296 ( .A(n_218), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g300 ( .A(n_218), .Y(n_300) );
INVx2_ASAP7_75t_L g314 ( .A(n_218), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_218), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g371 ( .A(n_218), .B(n_366), .Y(n_371) );
AND2x2_ASAP7_75t_L g436 ( .A(n_218), .B(n_406), .Y(n_436) );
OR2x6_ASAP7_75t_L g218 ( .A(n_219), .B(n_229), .Y(n_218) );
AOI21xp5_ASAP7_75t_SL g219 ( .A1(n_220), .A2(n_221), .B(n_228), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_225), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_225), .A2(n_236), .B(n_237), .Y(n_235) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g264 ( .A(n_227), .Y(n_264) );
INVx1_ASAP7_75t_L g238 ( .A(n_228), .Y(n_238) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_228), .A2(n_526), .B(n_536), .Y(n_525) );
OA21x2_ASAP7_75t_L g547 ( .A1(n_228), .A2(n_548), .B(n_555), .Y(n_547) );
AND2x2_ASAP7_75t_L g277 ( .A(n_231), .B(n_255), .Y(n_277) );
INVx2_ASAP7_75t_L g297 ( .A(n_231), .Y(n_297) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_238), .B(n_239), .Y(n_231) );
INVx1_ASAP7_75t_L g302 ( .A(n_241), .Y(n_302) );
AND2x2_ASAP7_75t_L g348 ( .A(n_241), .B(n_296), .Y(n_348) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_254), .Y(n_241) );
INVx2_ASAP7_75t_L g287 ( .A(n_242), .Y(n_287) );
INVx1_ASAP7_75t_L g295 ( .A(n_242), .Y(n_295) );
AND2x2_ASAP7_75t_L g313 ( .A(n_242), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_242), .B(n_297), .Y(n_351) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_252), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_251), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_248), .B(n_250), .Y(n_246) );
AND2x2_ASAP7_75t_L g330 ( .A(n_254), .B(n_287), .Y(n_330) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g283 ( .A(n_255), .Y(n_283) );
AND2x2_ASAP7_75t_L g366 ( .A(n_255), .B(n_297), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_261), .B(n_263), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_261), .A2(n_471), .B(n_472), .Y(n_470) );
INVx1_ASAP7_75t_L g530 ( .A(n_261), .Y(n_530) );
OAI21xp5_ASAP7_75t_SL g266 ( .A1(n_267), .A2(n_273), .B(n_277), .Y(n_266) );
INVx1_ASAP7_75t_SL g311 ( .A(n_267), .Y(n_311) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_268), .B(n_275), .Y(n_368) );
INVx1_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g317 ( .A(n_269), .B(n_272), .Y(n_317) );
AND2x2_ASAP7_75t_L g346 ( .A(n_269), .B(n_290), .Y(n_346) );
OR2x2_ASAP7_75t_L g349 ( .A(n_269), .B(n_309), .Y(n_349) );
AOI222xp33_ASAP7_75t_L g413 ( .A1(n_270), .A2(n_362), .B1(n_414), .B2(n_415), .C1(n_417), .C2(n_419), .Y(n_413) );
BUFx2_ASAP7_75t_L g327 ( .A(n_272), .Y(n_327) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g316 ( .A(n_275), .B(n_317), .Y(n_316) );
INVx3_ASAP7_75t_SL g333 ( .A(n_275), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_275), .B(n_327), .Y(n_387) );
AND2x2_ASAP7_75t_L g322 ( .A(n_277), .B(n_282), .Y(n_322) );
INVx1_ASAP7_75t_L g341 ( .A(n_277), .Y(n_341) );
OAI221xp5_ASAP7_75t_SL g278 ( .A1(n_279), .A2(n_280), .B1(n_284), .B2(n_288), .C(n_292), .Y(n_278) );
OR2x2_ASAP7_75t_L g350 ( .A(n_280), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x2_ASAP7_75t_L g335 ( .A(n_282), .B(n_305), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_282), .B(n_295), .Y(n_375) );
AND2x2_ASAP7_75t_L g380 ( .A(n_282), .B(n_330), .Y(n_380) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_282), .Y(n_390) );
NAND2x1_ASAP7_75t_SL g401 ( .A(n_282), .B(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g286 ( .A(n_283), .B(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g306 ( .A(n_283), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_283), .B(n_301), .Y(n_332) );
INVx1_ASAP7_75t_L g398 ( .A(n_283), .Y(n_398) );
INVx1_ASAP7_75t_L g373 ( .A(n_284), .Y(n_373) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_L g385 ( .A(n_285), .Y(n_385) );
NOR2xp67_ASAP7_75t_L g397 ( .A(n_285), .B(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g402 ( .A(n_286), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_286), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g305 ( .A(n_287), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_287), .B(n_297), .Y(n_318) );
INVx1_ASAP7_75t_L g384 ( .A(n_287), .Y(n_384) );
INVx1_ASAP7_75t_L g405 ( .A(n_288), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OAI21xp5_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_298), .B(n_307), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
AND2x2_ASAP7_75t_L g438 ( .A(n_294), .B(n_371), .Y(n_438) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g406 ( .A(n_295), .B(n_366), .Y(n_406) );
AOI32xp33_ASAP7_75t_L g319 ( .A1(n_296), .A2(n_302), .A3(n_320), .B1(n_322), .B2(n_323), .Y(n_319) );
AOI322xp5_ASAP7_75t_L g421 ( .A1(n_296), .A2(n_328), .A3(n_411), .B1(n_422), .B2(n_423), .C1(n_424), .C2(n_426), .Y(n_421) );
INVx2_ASAP7_75t_L g301 ( .A(n_297), .Y(n_301) );
INVx1_ASAP7_75t_L g411 ( .A(n_297), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_302), .B1(n_303), .B2(n_304), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_299), .B(n_305), .Y(n_354) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_300), .B(n_366), .Y(n_416) );
INVx1_ASAP7_75t_L g303 ( .A(n_301), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_301), .B(n_330), .Y(n_420) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_309), .B(n_404), .Y(n_403) );
OAI221xp5_ASAP7_75t_SL g310 ( .A1(n_311), .A2(n_312), .B1(n_315), .B2(n_318), .C(n_319), .Y(n_310) );
OR2x2_ASAP7_75t_L g331 ( .A(n_312), .B(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g340 ( .A(n_312), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g365 ( .A(n_313), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g369 ( .A(n_323), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI221xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_329), .B1(n_331), .B2(n_333), .C(n_334), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_327), .A2(n_358), .B1(n_362), .B2(n_363), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_328), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g433 ( .A(n_328), .Y(n_433) );
INVx1_ASAP7_75t_L g427 ( .A(n_330), .Y(n_427) );
INVx1_ASAP7_75t_SL g362 ( .A(n_331), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_333), .B(n_361), .Y(n_423) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_338), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g404 ( .A(n_338), .Y(n_404) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
OAI221xp5_ASAP7_75t_SL g342 ( .A1(n_343), .A2(n_347), .B1(n_349), .B2(n_350), .C(n_352), .Y(n_342) );
NOR2xp33_ASAP7_75t_SL g343 ( .A(n_344), .B(n_346), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_344), .A2(n_362), .B1(n_408), .B2(n_409), .Y(n_407) );
CKINVDCx14_ASAP7_75t_R g347 ( .A(n_348), .Y(n_347) );
OAI21xp33_ASAP7_75t_L g426 ( .A1(n_349), .A2(n_427), .B(n_428), .Y(n_426) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR3xp33_ASAP7_75t_SL g355 ( .A(n_356), .B(n_388), .C(n_412), .Y(n_355) );
NAND4xp25_ASAP7_75t_L g356 ( .A(n_357), .B(n_364), .C(n_372), .D(n_379), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g435 ( .A(n_360), .Y(n_435) );
INVx3_ASAP7_75t_SL g429 ( .A(n_361), .Y(n_429) );
OR2x2_ASAP7_75t_L g434 ( .A(n_361), .B(n_435), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_367), .B1(n_369), .B2(n_371), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_366), .B(n_384), .Y(n_425) );
INVxp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI21xp5_ASAP7_75t_SL g372 ( .A1(n_373), .A2(n_374), .B(n_376), .Y(n_372) );
INVxp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
INVxp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI211xp5_ASAP7_75t_SL g388 ( .A1(n_389), .A2(n_391), .B(n_394), .C(n_407), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g422 ( .A(n_393), .Y(n_422) );
AOI222xp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_399), .B1(n_400), .B2(n_403), .C1(n_405), .C2(n_406), .Y(n_394) );
INVxp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NAND4xp25_ASAP7_75t_SL g431 ( .A(n_404), .B(n_432), .C(n_433), .D(n_434), .Y(n_431) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NAND3xp33_ASAP7_75t_SL g412 ( .A(n_413), .B(n_421), .C(n_430), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_436), .B1(n_437), .B2(n_438), .Y(n_430) );
AOI21xp33_ASAP7_75t_L g445 ( .A1(n_441), .A2(n_442), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_451), .B1(n_452), .B2(n_456), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g743 ( .A(n_449), .Y(n_743) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_653), .Y(n_457) );
NAND3xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_602), .C(n_644), .Y(n_458) );
AOI211xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_511), .B(n_556), .C(n_578), .Y(n_459) );
OAI211xp5_ASAP7_75t_SL g460 ( .A1(n_461), .A2(n_474), .B(n_495), .C(n_506), .Y(n_460) );
INVxp67_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_462), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g665 ( .A(n_462), .B(n_582), .Y(n_665) );
BUFx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g567 ( .A(n_463), .B(n_498), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_463), .B(n_485), .Y(n_684) );
INVx1_ASAP7_75t_L g702 ( .A(n_463), .Y(n_702) );
AND2x2_ASAP7_75t_L g711 ( .A(n_463), .B(n_599), .Y(n_711) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OR2x2_ASAP7_75t_L g594 ( .A(n_464), .B(n_485), .Y(n_594) );
AND2x2_ASAP7_75t_L g652 ( .A(n_464), .B(n_599), .Y(n_652) );
INVx1_ASAP7_75t_L g696 ( .A(n_464), .Y(n_696) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g573 ( .A(n_465), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g581 ( .A(n_465), .Y(n_581) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_465), .Y(n_621) );
INVxp67_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_483), .Y(n_475) );
AND2x2_ASAP7_75t_L g560 ( .A(n_476), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g593 ( .A(n_476), .Y(n_593) );
OR2x2_ASAP7_75t_L g719 ( .A(n_476), .B(n_720), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_476), .B(n_485), .Y(n_723) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g498 ( .A(n_477), .Y(n_498) );
INVx1_ASAP7_75t_L g509 ( .A(n_477), .Y(n_509) );
AND2x2_ASAP7_75t_L g582 ( .A(n_477), .B(n_500), .Y(n_582) );
AND2x2_ASAP7_75t_L g622 ( .A(n_477), .B(n_501), .Y(n_622) );
OAI21xp5_ASAP7_75t_L g548 ( .A1(n_482), .A2(n_549), .B(n_552), .Y(n_548) );
INVxp67_ASAP7_75t_L g664 ( .A(n_483), .Y(n_664) );
AND2x4_ASAP7_75t_L g689 ( .A(n_483), .B(n_582), .Y(n_689) );
BUFx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_SL g580 ( .A(n_484), .B(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g499 ( .A(n_485), .B(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g568 ( .A(n_485), .B(n_501), .Y(n_568) );
INVx1_ASAP7_75t_L g574 ( .A(n_485), .Y(n_574) );
INVx2_ASAP7_75t_L g600 ( .A(n_485), .Y(n_600) );
AND2x2_ASAP7_75t_L g616 ( .A(n_485), .B(n_617), .Y(n_616) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_489), .B(n_490), .Y(n_487) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_496), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_499), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx2_ASAP7_75t_L g571 ( .A(n_498), .Y(n_571) );
AND2x2_ASAP7_75t_L g679 ( .A(n_498), .B(n_500), .Y(n_679) );
AND2x2_ASAP7_75t_L g596 ( .A(n_499), .B(n_581), .Y(n_596) );
AND2x2_ASAP7_75t_L g695 ( .A(n_499), .B(n_696), .Y(n_695) );
NOR2xp67_ASAP7_75t_L g617 ( .A(n_500), .B(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g720 ( .A(n_500), .B(n_581), .Y(n_720) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx2_ASAP7_75t_L g510 ( .A(n_501), .Y(n_510) );
AND2x2_ASAP7_75t_L g599 ( .A(n_501), .B(n_600), .Y(n_599) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_504), .A2(n_532), .B(n_534), .C(n_535), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_504), .A2(n_544), .B(n_545), .Y(n_543) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_510), .Y(n_507) );
AND2x2_ASAP7_75t_L g645 ( .A(n_508), .B(n_580), .Y(n_645) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_509), .B(n_581), .Y(n_630) );
INVx2_ASAP7_75t_L g629 ( .A(n_510), .Y(n_629) );
OAI222xp33_ASAP7_75t_L g633 ( .A1(n_510), .A2(n_573), .B1(n_634), .B2(n_636), .C1(n_637), .C2(n_640), .Y(n_633) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_522), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g558 ( .A(n_515), .Y(n_558) );
OR2x2_ASAP7_75t_L g669 ( .A(n_515), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx3_ASAP7_75t_L g591 ( .A(n_516), .Y(n_591) );
NOR2x1_ASAP7_75t_L g642 ( .A(n_516), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g648 ( .A(n_516), .B(n_562), .Y(n_648) );
AND2x4_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
INVx1_ASAP7_75t_L g609 ( .A(n_517), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_522), .A2(n_612), .B1(n_651), .B2(n_652), .Y(n_650) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_537), .Y(n_522) );
INVx3_ASAP7_75t_L g584 ( .A(n_523), .Y(n_584) );
OR2x2_ASAP7_75t_L g717 ( .A(n_523), .B(n_593), .Y(n_717) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g590 ( .A(n_524), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g606 ( .A(n_524), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g614 ( .A(n_524), .B(n_562), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_524), .B(n_538), .Y(n_670) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g561 ( .A(n_525), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g565 ( .A(n_525), .B(n_538), .Y(n_565) );
AND2x2_ASAP7_75t_L g641 ( .A(n_525), .B(n_588), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_525), .B(n_547), .Y(n_681) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_537), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g597 ( .A(n_537), .B(n_558), .Y(n_597) );
AND2x2_ASAP7_75t_L g601 ( .A(n_537), .B(n_591), .Y(n_601) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_547), .Y(n_537) );
INVx3_ASAP7_75t_L g562 ( .A(n_538), .Y(n_562) );
AND2x2_ASAP7_75t_L g587 ( .A(n_538), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g722 ( .A(n_538), .B(n_705), .Y(n_722) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_547), .Y(n_576) );
INVx2_ASAP7_75t_L g588 ( .A(n_547), .Y(n_588) );
AND2x2_ASAP7_75t_L g632 ( .A(n_547), .B(n_608), .Y(n_632) );
INVx1_ASAP7_75t_L g675 ( .A(n_547), .Y(n_675) );
OR2x2_ASAP7_75t_L g706 ( .A(n_547), .B(n_608), .Y(n_706) );
AND2x2_ASAP7_75t_L g726 ( .A(n_547), .B(n_562), .Y(n_726) );
OAI21xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_559), .B(n_563), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g564 ( .A(n_558), .B(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_558), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g683 ( .A(n_560), .Y(n_683) );
INVx2_ASAP7_75t_SL g577 ( .A(n_561), .Y(n_577) );
AND2x2_ASAP7_75t_L g697 ( .A(n_561), .B(n_591), .Y(n_697) );
INVx2_ASAP7_75t_L g643 ( .A(n_562), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_562), .B(n_675), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_566), .B1(n_569), .B2(n_575), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_565), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_SL g731 ( .A(n_565), .Y(n_731) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx1_ASAP7_75t_L g656 ( .A(n_567), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_567), .B(n_599), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_568), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g672 ( .A(n_568), .B(n_621), .Y(n_672) );
INVx2_ASAP7_75t_L g728 ( .A(n_568), .Y(n_728) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
AND2x2_ASAP7_75t_L g598 ( .A(n_571), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_571), .B(n_616), .Y(n_649) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_573), .B(n_593), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
INVx1_ASAP7_75t_L g710 ( .A(n_576), .Y(n_710) );
O2A1O1Ixp33_ASAP7_75t_SL g660 ( .A1(n_577), .A2(n_661), .B(n_663), .C(n_666), .Y(n_660) );
OR2x2_ASAP7_75t_L g687 ( .A(n_577), .B(n_591), .Y(n_687) );
OAI221xp5_ASAP7_75t_SL g578 ( .A1(n_579), .A2(n_583), .B1(n_585), .B2(n_592), .C(n_595), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_580), .B(n_582), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_580), .B(n_629), .Y(n_636) );
AND2x2_ASAP7_75t_L g678 ( .A(n_580), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g714 ( .A(n_580), .Y(n_714) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_581), .Y(n_605) );
INVx1_ASAP7_75t_L g618 ( .A(n_581), .Y(n_618) );
NOR2xp67_ASAP7_75t_L g638 ( .A(n_584), .B(n_639), .Y(n_638) );
INVxp67_ASAP7_75t_L g692 ( .A(n_584), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_584), .B(n_632), .Y(n_708) );
INVx2_ASAP7_75t_L g694 ( .A(n_585), .Y(n_694) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_589), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g635 ( .A(n_587), .B(n_606), .Y(n_635) );
O2A1O1Ixp33_ASAP7_75t_L g644 ( .A1(n_587), .A2(n_603), .B(n_645), .C(n_646), .Y(n_644) );
AND2x2_ASAP7_75t_L g613 ( .A(n_588), .B(n_608), .Y(n_613) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_592), .B(n_691), .Y(n_690) );
OR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
OR2x2_ASAP7_75t_L g661 ( .A(n_593), .B(n_662), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_597), .B1(n_598), .B2(n_601), .Y(n_595) );
INVx1_ASAP7_75t_L g715 ( .A(n_597), .Y(n_715) );
INVx1_ASAP7_75t_L g662 ( .A(n_599), .Y(n_662) );
INVx1_ASAP7_75t_L g713 ( .A(n_601), .Y(n_713) );
AOI211xp5_ASAP7_75t_SL g602 ( .A1(n_603), .A2(n_606), .B(n_610), .C(n_633), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g625 ( .A(n_605), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g676 ( .A(n_606), .Y(n_676) );
AND2x2_ASAP7_75t_L g725 ( .A(n_606), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OAI21xp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_615), .B(n_623), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx2_ASAP7_75t_L g639 ( .A(n_613), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_613), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g631 ( .A(n_614), .B(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g707 ( .A(n_614), .Y(n_707) );
OAI32xp33_ASAP7_75t_L g718 ( .A1(n_614), .A2(n_666), .A3(n_673), .B1(n_714), .B2(n_719), .Y(n_718) );
NOR2xp33_ASAP7_75t_SL g615 ( .A(n_616), .B(n_619), .Y(n_615) );
INVx1_ASAP7_75t_SL g686 ( .A(n_616), .Y(n_686) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_SL g626 ( .A(n_622), .Y(n_626) );
OAI21xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_627), .B(n_631), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI22xp33_ASAP7_75t_L g698 ( .A1(n_625), .A2(n_673), .B1(n_699), .B2(n_701), .Y(n_698) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_629), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g666 ( .A(n_632), .Y(n_666) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2x1p5_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
INVx1_ASAP7_75t_L g659 ( .A(n_643), .Y(n_659) );
OAI21xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_649), .B(n_650), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_652), .A2(n_694), .B1(n_695), .B2(n_697), .C(n_698), .Y(n_693) );
NAND5xp2_ASAP7_75t_L g653 ( .A(n_654), .B(n_677), .C(n_693), .D(n_703), .E(n_721), .Y(n_653) );
AOI211xp5_ASAP7_75t_SL g654 ( .A1(n_655), .A2(n_657), .B(n_660), .C(n_667), .Y(n_654) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g724 ( .A(n_661), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
OAI22xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B1(n_671), .B2(n_673), .Y(n_667) );
INVx1_ASAP7_75t_SL g700 ( .A(n_670), .Y(n_700) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OAI322xp33_ASAP7_75t_L g682 ( .A1(n_673), .A2(n_683), .A3(n_684), .B1(n_685), .B2(n_686), .C1(n_687), .C2(n_688), .Y(n_682) );
OR2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_676), .Y(n_673) );
INVx1_ASAP7_75t_L g685 ( .A(n_675), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_675), .B(n_700), .Y(n_699) );
AOI211xp5_ASAP7_75t_SL g677 ( .A1(n_678), .A2(n_680), .B(n_682), .C(n_690), .Y(n_677) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OAI22xp33_ASAP7_75t_L g712 ( .A1(n_686), .A2(n_713), .B1(n_714), .B2(n_715), .Y(n_712) );
INVx1_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g729 ( .A(n_696), .Y(n_729) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_711), .B1(n_712), .B2(n_716), .C(n_718), .Y(n_703) );
OAI211xp5_ASAP7_75t_SL g704 ( .A1(n_705), .A2(n_707), .B(n_708), .C(n_709), .Y(n_704) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
OR2x2_ASAP7_75t_L g730 ( .A(n_706), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B1(n_724), .B2(n_725), .C(n_727), .Y(n_721) );
AOI21xp33_ASAP7_75t_SL g727 ( .A1(n_728), .A2(n_729), .B(n_730), .Y(n_727) );
CKINVDCx16_ASAP7_75t_R g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_745), .Y(n_744) );
endmodule