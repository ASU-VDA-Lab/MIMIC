module fake_jpeg_14094_n_250 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_1),
.B(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_40),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_41),
.B(n_44),
.Y(n_97)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_46),
.Y(n_79)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g96 ( 
.A(n_51),
.Y(n_96)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_29),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_61),
.Y(n_83)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_63),
.Y(n_67)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_0),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_64),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_19),
.B(n_16),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_23),
.B(n_15),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_66),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_38),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_70),
.B(n_72),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_22),
.B1(n_38),
.B2(n_23),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g127 ( 
.A1(n_71),
.A2(n_78),
.B1(n_95),
.B2(n_99),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_35),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_36),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_73),
.B(n_80),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_22),
.B1(n_35),
.B2(n_28),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_36),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_40),
.A2(n_22),
.B1(n_25),
.B2(n_31),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_84),
.B1(n_91),
.B2(n_58),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_43),
.A2(n_25),
.B1(n_31),
.B2(n_29),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_28),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_43),
.B(n_26),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_46),
.A2(n_25),
.B1(n_31),
.B2(n_33),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_60),
.A2(n_37),
.B1(n_34),
.B2(n_33),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_51),
.B1(n_48),
.B2(n_57),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_45),
.A2(n_26),
.B1(n_34),
.B2(n_30),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_49),
.A2(n_37),
.B1(n_30),
.B2(n_18),
.Y(n_99)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_105),
.A2(n_76),
.B1(n_101),
.B2(n_94),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_106),
.A2(n_111),
.B1(n_98),
.B2(n_93),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_17),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_110),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_66),
.C(n_51),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_123),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_1),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_121),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_15),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_76),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_47),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_115),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_2),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g152 ( 
.A1(n_113),
.A2(n_120),
.B(n_122),
.Y(n_152)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

NOR2x1_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_3),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_128),
.B1(n_130),
.B2(n_76),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_3),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_5),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_5),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_79),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_90),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_131),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_89),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_85),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g130 ( 
.A1(n_93),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_11),
.Y(n_132)
);

AOI21xp33_ASAP7_75t_L g138 ( 
.A1(n_132),
.A2(n_96),
.B(n_13),
.Y(n_138)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_133),
.Y(n_136)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_134),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_135),
.Y(n_162)
);

NOR3xp33_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_145),
.C(n_149),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_75),
.B(n_96),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_141),
.A2(n_158),
.B(n_159),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_125),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_120),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_109),
.B(n_115),
.C(n_103),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_105),
.B1(n_126),
.B2(n_127),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_160),
.Y(n_172)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_SL g149 ( 
.A(n_119),
.B(n_89),
.C(n_75),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_113),
.A2(n_93),
.B(n_94),
.C(n_101),
.Y(n_153)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_154),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_98),
.B(n_69),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_122),
.A2(n_98),
.B(n_13),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_69),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_167),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_137),
.B(n_118),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_152),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_142),
.B(n_116),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_137),
.B(n_127),
.Y(n_169)
);

A2O1A1O1Ixp25_ASAP7_75t_L g197 ( 
.A1(n_169),
.A2(n_176),
.B(n_177),
.C(n_135),
.D(n_153),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_151),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_181),
.Y(n_186)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_146),
.A2(n_157),
.B1(n_141),
.B2(n_158),
.Y(n_175)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_157),
.B(n_124),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_104),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_114),
.C(n_131),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_179),
.C(n_156),
.Y(n_194)
);

AND2x2_ASAP7_75t_SL g179 ( 
.A(n_139),
.B(n_117),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_133),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_136),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_171),
.A2(n_147),
.B(n_159),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_183),
.A2(n_199),
.B(n_166),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_167),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_191),
.Y(n_210)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_172),
.A2(n_147),
.A3(n_145),
.B1(n_160),
.B2(n_159),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_197),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_187),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_194),
.C(n_198),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_176),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_144),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_192),
.B(n_195),
.Y(n_204)
);

NOR3xp33_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_149),
.C(n_156),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_153),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_130),
.B(n_136),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_162),
.B1(n_168),
.B2(n_172),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_199),
.B1(n_166),
.B2(n_193),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_200),
.A2(n_163),
.B(n_179),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_212),
.B(n_180),
.Y(n_224)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_190),
.Y(n_203)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_211),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_178),
.C(n_179),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_209),
.C(n_213),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_179),
.C(n_177),
.Y(n_209)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_188),
.A2(n_186),
.A3(n_168),
.B1(n_196),
.B2(n_198),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_164),
.C(n_162),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_210),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_217),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_205),
.B(n_188),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_150),
.Y(n_231)
);

NOR3xp33_ASAP7_75t_SL g217 ( 
.A(n_206),
.B(n_165),
.C(n_183),
.Y(n_217)
);

NAND3xp33_ASAP7_75t_SL g221 ( 
.A(n_206),
.B(n_185),
.C(n_197),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_211),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_222),
.A2(n_202),
.B1(n_209),
.B2(n_208),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_193),
.C(n_174),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_173),
.C(n_181),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_224),
.A2(n_123),
.B1(n_140),
.B2(n_129),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_226),
.A2(n_217),
.B(n_230),
.C(n_220),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_219),
.A2(n_214),
.B1(n_204),
.B2(n_212),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_228),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_219),
.A2(n_180),
.B1(n_213),
.B2(n_207),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_229),
.A2(n_218),
.B1(n_224),
.B2(n_223),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_232),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_216),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_235),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_220),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_237),
.A2(n_226),
.B1(n_229),
.B2(n_232),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_238),
.A2(n_218),
.B1(n_231),
.B2(n_140),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_241),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_235),
.A2(n_233),
.B(n_236),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_240),
.B(n_242),
.Y(n_245)
);

BUFx24_ASAP7_75t_SL g242 ( 
.A(n_235),
.Y(n_242)
);

NAND2xp33_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_143),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_69),
.B(n_82),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_150),
.C(n_134),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_247),
.A2(n_248),
.B(n_246),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_249),
.B(n_82),
.Y(n_250)
);


endmodule