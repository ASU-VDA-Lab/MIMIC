module fake_jpeg_21735_n_299 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_299);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_299;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_247;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_273;
wire n_200;
wire n_86;
wire n_156;
wire n_265;
wire n_115;
wire n_123;
wire n_192;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_14),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_26),
.Y(n_57)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_48),
.Y(n_64)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_52),
.B(n_37),
.Y(n_78)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_24),
.B1(n_23),
.B2(n_15),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_56),
.A2(n_16),
.B1(n_31),
.B2(n_30),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_57),
.B(n_78),
.Y(n_102)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_73),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_67),
.B1(n_82),
.B2(n_28),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_66),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_41),
.A2(n_23),
.B1(n_26),
.B2(n_28),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_45),
.A2(n_23),
.B1(n_22),
.B2(n_35),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_69),
.A2(n_75),
.B(n_36),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx2_ASAP7_75t_SL g74 ( 
.A(n_46),
.Y(n_74)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_37),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_80),
.Y(n_94)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_15),
.B1(n_31),
.B2(n_30),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_28),
.B1(n_25),
.B2(n_20),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_47),
.A2(n_16),
.B1(n_31),
.B2(n_30),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_46),
.Y(n_83)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_15),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_89),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_16),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_0),
.B(n_1),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_104),
.B(n_99),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_37),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_95),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_93),
.A2(n_99),
.B1(n_20),
.B2(n_71),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_36),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_96),
.B(n_21),
.Y(n_129)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_68),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_103),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_104),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_68),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_36),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_60),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_35),
.C(n_17),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_17),
.C(n_27),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_105),
.A2(n_69),
.B1(n_45),
.B2(n_76),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_114),
.A2(n_120),
.B1(n_137),
.B2(n_111),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_69),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_118),
.B(n_108),
.Y(n_143)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_116),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_121),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_106),
.A2(n_69),
.B1(n_80),
.B2(n_77),
.Y(n_120)
);

NOR3xp33_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_20),
.C(n_25),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_85),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_134),
.Y(n_144)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_127),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_126),
.B(n_129),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_35),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_138),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_102),
.B(n_87),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_130),
.B(n_109),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_90),
.A2(n_61),
.B1(n_55),
.B2(n_83),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_131),
.A2(n_108),
.B(n_107),
.Y(n_146)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_64),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_136),
.B(n_29),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_96),
.A2(n_72),
.B1(n_70),
.B2(n_19),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_109),
.B(n_72),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_17),
.C(n_22),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_147),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_143),
.A2(n_152),
.B(n_153),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_145),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_146),
.A2(n_139),
.B1(n_136),
.B2(n_132),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_135),
.B(n_14),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_97),
.B1(n_84),
.B2(n_88),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_148),
.A2(n_155),
.B1(n_158),
.B2(n_162),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_113),
.A2(n_124),
.B1(n_116),
.B2(n_119),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_160),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_115),
.A2(n_84),
.B1(n_88),
.B2(n_101),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_150),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_117),
.A2(n_107),
.B1(n_101),
.B2(n_111),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_151),
.A2(n_169),
.B1(n_5),
.B2(n_6),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_113),
.B(n_115),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_118),
.A2(n_111),
.B(n_98),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_119),
.A2(n_22),
.B(n_100),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_156),
.A2(n_0),
.B(n_1),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_114),
.A2(n_100),
.B1(n_11),
.B2(n_12),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_120),
.B(n_27),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_159),
.A2(n_123),
.B(n_122),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_129),
.A2(n_21),
.B1(n_19),
.B2(n_29),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_29),
.B1(n_27),
.B2(n_21),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_127),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_165),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_196)
);

NOR3xp33_ASAP7_75t_SL g166 ( 
.A(n_138),
.B(n_21),
.C(n_19),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_167),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_126),
.A2(n_19),
.B1(n_27),
.B2(n_29),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_9),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_112),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_133),
.C(n_17),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g171 ( 
.A1(n_157),
.A2(n_130),
.A3(n_133),
.B1(n_131),
.B2(n_112),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_156),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_144),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_175),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_176),
.A2(n_177),
.B(n_184),
.Y(n_219)
);

NOR2x1_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_170),
.C(n_153),
.Y(n_204)
);

OA21x2_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_22),
.B(n_17),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_182),
.A2(n_190),
.B1(n_193),
.B2(n_194),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_10),
.Y(n_183)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_186),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_147),
.Y(n_187)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_187),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_0),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_189),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_2),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_2),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_2),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_195),
.A2(n_198),
.B1(n_158),
.B2(n_146),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_196),
.A2(n_197),
.B1(n_160),
.B2(n_167),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_155),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_143),
.B(n_5),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_165),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_205),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_219),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_149),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_210),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_142),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_142),
.C(n_159),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_176),
.C(n_177),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_213),
.A2(n_215),
.B1(n_220),
.B2(n_180),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_172),
.A2(n_200),
.B1(n_178),
.B2(n_159),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_173),
.B(n_148),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_172),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_199),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_223),
.Y(n_242)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_217),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_218),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_230),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_227),
.C(n_231),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_175),
.C(n_186),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_202),
.B(n_212),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_228),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_178),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_193),
.C(n_180),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_232),
.A2(n_159),
.B1(n_214),
.B2(n_197),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_216),
.B(n_174),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_234),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_201),
.C(n_221),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_238),
.C(n_182),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_203),
.B(n_141),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_237),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_203),
.B(n_141),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_207),
.B(n_190),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_230),
.A2(n_206),
.B(n_200),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_248),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_SL g243 ( 
.A1(n_234),
.A2(n_215),
.B(n_219),
.C(n_220),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

XOR2x1_ASAP7_75t_SL g244 ( 
.A(n_226),
.B(n_222),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_246),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_189),
.Y(n_245)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_245),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_227),
.A2(n_213),
.B1(n_181),
.B2(n_157),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_250),
.A2(n_229),
.B1(n_224),
.B2(n_195),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_235),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_229),
.A2(n_184),
.B(n_181),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_224),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_261),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_251),
.C(n_245),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_250),
.C(n_248),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_264),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_253),
.C(n_243),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_252),
.A2(n_194),
.B(n_188),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_263),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_249),
.Y(n_264)
);

FAx1_ASAP7_75t_SL g265 ( 
.A(n_240),
.B(n_182),
.CI(n_168),
.CON(n_265),
.SN(n_265)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_265),
.B(n_196),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_209),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_243),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_255),
.A2(n_244),
.B(n_241),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_267),
.A2(n_256),
.B(n_264),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_269),
.B(n_276),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_271),
.B(n_273),
.Y(n_277)
);

XOR2x1_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_243),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_275),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_192),
.C(n_191),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_272),
.A2(n_247),
.B1(n_260),
.B2(n_268),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_279),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_273),
.A2(n_247),
.B1(n_266),
.B2(n_257),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_281),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_265),
.B(n_192),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_269),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_275),
.A2(n_166),
.B(n_192),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_284),
.A2(n_166),
.B(n_162),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_277),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_287),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_145),
.C(n_7),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_282),
.C(n_277),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_292),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_285),
.C(n_288),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_288),
.B(n_8),
.C(n_9),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_295),
.A2(n_293),
.B(n_8),
.Y(n_296)
);

OAI21x1_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_9),
.B(n_6),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_6),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_8),
.B(n_277),
.Y(n_299)
);


endmodule