module fake_ariane_1163_n_1840 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_387, n_406, n_117, n_139, n_85, n_130, n_349, n_391, n_346, n_214, n_348, n_2, n_462, n_32, n_410, n_379, n_445, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_267, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_398, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_439, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_432, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_390, n_104, n_438, n_314, n_16, n_440, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_17, n_225, n_235, n_464, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_135, n_409, n_171, n_384, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_460, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_454, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_418, n_223, n_403, n_25, n_83, n_389, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_430, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_428, n_159, n_358, n_105, n_30, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_457, n_164, n_157, n_184, n_177, n_364, n_258, n_425, n_431, n_118, n_121, n_411, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_80, n_211, n_97, n_408, n_322, n_251, n_116, n_397, n_351, n_39, n_393, n_359, n_155, n_127, n_1840);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_387;
input n_406;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_346;
input n_214;
input n_348;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_267;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_398;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_439;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_432;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_104;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_464;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_135;
input n_409;
input n_171;
input n_384;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_460;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_430;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_425;
input n_431;
input n_118;
input n_121;
input n_411;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_80;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_116;
input n_397;
input n_351;
input n_39;
input n_393;
input n_359;
input n_155;
input n_127;

output n_1840;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_1383;
wire n_603;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_1713;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_764;
wire n_1503;
wire n_1196;
wire n_1181;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_813;
wire n_995;
wire n_1184;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_1703;
wire n_899;
wire n_611;
wire n_1295;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_1751;
wire n_533;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_1396;
wire n_1230;
wire n_612;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1716;
wire n_1585;
wire n_1432;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1555;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1680;
wire n_964;
wire n_1627;
wire n_489;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_471;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_698;
wire n_1674;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_706;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_1817;
wire n_552;
wire n_670;
wire n_1826;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_1467;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_1726;
wire n_1015;
wire n_545;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_1156;
wire n_501;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_1402;
wire n_957;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_1708;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_1733;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1208;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_673;
wire n_1038;
wire n_571;
wire n_1521;
wire n_1694;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_519;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_1687;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_621;
wire n_1587;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_1735;
wire n_1788;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_765;
wire n_1809;
wire n_1268;
wire n_917;
wire n_1271;
wire n_1530;
wire n_631;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_1813;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1344;
wire n_1390;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1136;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_946;
wire n_757;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_1434;
wire n_1569;
wire n_548;
wire n_523;
wire n_1662;
wire n_1299;
wire n_782;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_484;
wire n_849;
wire n_1820;
wire n_1251;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_159),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_404),
.Y(n_466)
);

BUFx10_ASAP7_75t_L g467 ( 
.A(n_392),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_348),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_105),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_375),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_10),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_446),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_120),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_37),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_43),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_432),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_346),
.Y(n_477)
);

BUFx10_ASAP7_75t_L g478 ( 
.A(n_415),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_296),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_462),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_205),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_449),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_320),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_62),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_138),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_184),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_350),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_36),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_322),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_340),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_132),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_372),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_457),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_254),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_402),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_255),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_317),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_403),
.Y(n_498)
);

BUFx5_ASAP7_75t_L g499 ( 
.A(n_460),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_154),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_74),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_267),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_218),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_344),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_363),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_121),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_122),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_82),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_133),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_135),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_416),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_452),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_345),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_422),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_331),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_82),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_64),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_79),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_302),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_96),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_11),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_178),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_108),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_179),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_171),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_335),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_48),
.Y(n_527)
);

BUFx10_ASAP7_75t_L g528 ( 
.A(n_433),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_359),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_353),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_21),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_319),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_389),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_417),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_9),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_461),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_229),
.Y(n_537)
);

CKINVDCx16_ASAP7_75t_R g538 ( 
.A(n_57),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_248),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_130),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_102),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_418),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g543 ( 
.A(n_242),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_341),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_164),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_455),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_220),
.Y(n_547)
);

BUFx5_ASAP7_75t_L g548 ( 
.A(n_107),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_60),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_312),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_194),
.Y(n_551)
);

CKINVDCx6p67_ASAP7_75t_R g552 ( 
.A(n_227),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_77),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_111),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_285),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_38),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_456),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_219),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_202),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_193),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_31),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_450),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_291),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_286),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_22),
.Y(n_565)
);

CKINVDCx16_ASAP7_75t_R g566 ( 
.A(n_441),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_385),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_115),
.Y(n_568)
);

BUFx8_ASAP7_75t_SL g569 ( 
.A(n_213),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_156),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_91),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_241),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_216),
.Y(n_573)
);

CKINVDCx14_ASAP7_75t_R g574 ( 
.A(n_77),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_257),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_141),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_91),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_1),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_18),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_56),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_83),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_306),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_412),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_459),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_185),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_354),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_25),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_32),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_97),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_95),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_14),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_391),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_35),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_163),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_454),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_447),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_238),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_300),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_436),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_239),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_448),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_362),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_83),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_256),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_49),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_327),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_5),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_207),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_121),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_234),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_182),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_71),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_288),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_260),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_35),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_31),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_463),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_195),
.Y(n_618)
);

CKINVDCx14_ASAP7_75t_R g619 ( 
.A(n_269),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_107),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_186),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_458),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_5),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_377),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_68),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_443),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_124),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_333),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_25),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_29),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_409),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_378),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_73),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_86),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_84),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_224),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_51),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_453),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_73),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_451),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_569),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_569),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_574),
.Y(n_643)
);

INVxp33_ASAP7_75t_SL g644 ( 
.A(n_535),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_538),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_574),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_568),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_519),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_568),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_571),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_479),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_552),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_571),
.Y(n_653)
);

CKINVDCx16_ASAP7_75t_R g654 ( 
.A(n_483),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_548),
.Y(n_655)
);

INVxp67_ASAP7_75t_SL g656 ( 
.A(n_471),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_548),
.Y(n_657)
);

INVx4_ASAP7_75t_R g658 ( 
.A(n_479),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_519),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_548),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_556),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_548),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_548),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_548),
.Y(n_664)
);

INVxp67_ASAP7_75t_SL g665 ( 
.A(n_473),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_517),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_520),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_486),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_523),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_549),
.Y(n_670)
);

INVxp67_ASAP7_75t_SL g671 ( 
.A(n_553),
.Y(n_671)
);

XOR2x2_ASAP7_75t_L g672 ( 
.A(n_612),
.B(n_0),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_561),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_565),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_485),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_485),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_579),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_515),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_589),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_515),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_593),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_633),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_615),
.Y(n_683)
);

INVxp67_ASAP7_75t_SL g684 ( 
.A(n_620),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_532),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_532),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_623),
.Y(n_687)
);

CKINVDCx14_ASAP7_75t_R g688 ( 
.A(n_619),
.Y(n_688)
);

INVxp33_ASAP7_75t_L g689 ( 
.A(n_630),
.Y(n_689)
);

CKINVDCx14_ASAP7_75t_R g690 ( 
.A(n_619),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_639),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_513),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_547),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_542),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_467),
.Y(n_695)
);

BUFx10_ASAP7_75t_L g696 ( 
.A(n_469),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_467),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_478),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_478),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_528),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_528),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_547),
.Y(n_702)
);

INVxp33_ASAP7_75t_L g703 ( 
.A(n_497),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_466),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_472),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_476),
.Y(n_706)
);

CKINVDCx14_ASAP7_75t_R g707 ( 
.A(n_494),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_499),
.Y(n_708)
);

CKINVDCx16_ASAP7_75t_R g709 ( 
.A(n_566),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_499),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_490),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_492),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_474),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_495),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_500),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_502),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_505),
.Y(n_717)
);

INVxp33_ASAP7_75t_L g718 ( 
.A(n_497),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_499),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_512),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_526),
.Y(n_721)
);

INVxp33_ASAP7_75t_SL g722 ( 
.A(n_475),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_530),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_536),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_537),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_539),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_499),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_558),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_499),
.Y(n_729)
);

INVxp67_ASAP7_75t_SL g730 ( 
.A(n_524),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_563),
.Y(n_731)
);

INVxp33_ASAP7_75t_SL g732 ( 
.A(n_484),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_501),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_576),
.Y(n_734)
);

INVxp67_ASAP7_75t_SL g735 ( 
.A(n_524),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_583),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_516),
.Y(n_737)
);

INVxp33_ASAP7_75t_SL g738 ( 
.A(n_506),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_507),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_629),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_508),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_655),
.Y(n_742)
);

AND2x6_ASAP7_75t_L g743 ( 
.A(n_708),
.B(n_525),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_651),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_651),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_651),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_657),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_660),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_696),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_651),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_739),
.Y(n_751)
);

INVx6_ASAP7_75t_L g752 ( 
.A(n_686),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_662),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_663),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_688),
.B(n_488),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_686),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_737),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_675),
.B(n_596),
.Y(n_758)
);

OA21x2_ASAP7_75t_L g759 ( 
.A1(n_664),
.A2(n_529),
.B(n_525),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_666),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_695),
.B(n_529),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_688),
.B(n_590),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_697),
.B(n_698),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_667),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_708),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_686),
.Y(n_766)
);

INVx5_ASAP7_75t_L g767 ( 
.A(n_686),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_699),
.B(n_640),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_669),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_675),
.B(n_599),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_670),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_710),
.Y(n_772)
);

BUFx2_ASAP7_75t_L g773 ( 
.A(n_645),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_L g774 ( 
.A1(n_644),
.A2(n_603),
.B1(n_521),
.B2(n_527),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_SL g775 ( 
.A1(n_648),
.A2(n_531),
.B1(n_541),
.B2(n_518),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_676),
.B(n_678),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_710),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_693),
.Y(n_778)
);

BUFx12f_ASAP7_75t_L g779 ( 
.A(n_641),
.Y(n_779)
);

XNOR2xp5_ASAP7_75t_L g780 ( 
.A(n_659),
.B(n_554),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_703),
.B(n_567),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_719),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_661),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_674),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_661),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_690),
.B(n_577),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_693),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_677),
.Y(n_788)
);

INVx4_ASAP7_75t_L g789 ( 
.A(n_652),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_679),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_676),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_719),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_678),
.B(n_602),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_642),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_668),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_727),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_680),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_727),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_694),
.B(n_578),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_729),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_729),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_700),
.B(n_567),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_690),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_680),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_685),
.Y(n_805)
);

OA21x2_ASAP7_75t_L g806 ( 
.A1(n_704),
.A2(n_595),
.B(n_573),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_681),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_685),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_739),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_702),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_683),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_702),
.B(n_611),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_647),
.Y(n_813)
);

BUFx12f_ASAP7_75t_L g814 ( 
.A(n_696),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_649),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_740),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_654),
.A2(n_581),
.B1(n_587),
.B2(n_580),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_650),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_709),
.A2(n_591),
.B1(n_605),
.B2(n_588),
.Y(n_819)
);

INVx5_ASAP7_75t_L g820 ( 
.A(n_658),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_653),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_705),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_687),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_707),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_722),
.A2(n_609),
.B1(n_616),
.B2(n_607),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_706),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_707),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_776),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_751),
.B(n_713),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_776),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_813),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_818),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_742),
.B(n_703),
.Y(n_833)
);

BUFx2_ASAP7_75t_L g834 ( 
.A(n_795),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_765),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_783),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_765),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_747),
.B(n_718),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_821),
.Y(n_839)
);

AND2x6_ASAP7_75t_L g840 ( 
.A(n_755),
.B(n_573),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_791),
.Y(n_841)
);

NAND2xp33_ASAP7_75t_SL g842 ( 
.A(n_749),
.B(n_718),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_744),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_801),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_791),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_804),
.Y(n_846)
);

OA21x2_ASAP7_75t_L g847 ( 
.A1(n_801),
.A2(n_712),
.B(n_711),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_751),
.B(n_741),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_820),
.B(n_792),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_809),
.B(n_689),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_772),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_792),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_748),
.B(n_730),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_792),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_783),
.Y(n_855)
);

OAI21x1_ASAP7_75t_L g856 ( 
.A1(n_777),
.A2(n_796),
.B(n_782),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_753),
.B(n_735),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_797),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_797),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_760),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_754),
.B(n_701),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_800),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_798),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_800),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_764),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_744),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_744),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_800),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_769),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_759),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_771),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_820),
.B(n_714),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_784),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_788),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_790),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_757),
.Y(n_876)
);

OR2x6_ASAP7_75t_L g877 ( 
.A(n_779),
.B(n_673),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_759),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_805),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_785),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_807),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_763),
.B(n_762),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_811),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_805),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_805),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_808),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_808),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_809),
.B(n_689),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_820),
.B(n_715),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_823),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_785),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_815),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_815),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_820),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_808),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_810),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_795),
.Y(n_897)
);

INVx6_ASAP7_75t_L g898 ( 
.A(n_778),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_810),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_746),
.Y(n_900)
);

NAND2xp33_ASAP7_75t_SL g901 ( 
.A(n_803),
.B(n_643),
.Y(n_901)
);

NAND2x1_ASAP7_75t_L g902 ( 
.A(n_743),
.B(n_716),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_746),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_810),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_822),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_746),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_822),
.B(n_717),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_826),
.B(n_720),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_752),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_773),
.B(n_646),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_826),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_745),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_745),
.Y(n_913)
);

NAND2xp33_ASAP7_75t_SL g914 ( 
.A(n_803),
.B(n_625),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_750),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_766),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_766),
.Y(n_917)
);

BUFx2_ASAP7_75t_L g918 ( 
.A(n_824),
.Y(n_918)
);

CKINVDCx16_ASAP7_75t_R g919 ( 
.A(n_814),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_778),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_860),
.Y(n_921)
);

BUFx10_ASAP7_75t_L g922 ( 
.A(n_882),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_835),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_829),
.B(n_732),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_865),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_850),
.Y(n_926)
);

BUFx4f_ASAP7_75t_L g927 ( 
.A(n_877),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_869),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_847),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_835),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_871),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_828),
.B(n_781),
.Y(n_932)
);

XOR2xp5_ASAP7_75t_SL g933 ( 
.A(n_897),
.B(n_825),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_876),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_888),
.B(n_794),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_SL g936 ( 
.A(n_840),
.B(n_789),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_847),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_847),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_848),
.B(n_789),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_830),
.B(n_781),
.Y(n_940)
);

INVx4_ASAP7_75t_L g941 ( 
.A(n_894),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_882),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_837),
.B(n_806),
.Y(n_943)
);

INVx2_ASAP7_75t_SL g944 ( 
.A(n_836),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_876),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_L g946 ( 
.A1(n_840),
.A2(n_774),
.B1(n_802),
.B2(n_761),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_837),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_855),
.B(n_824),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_844),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_844),
.B(n_806),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_834),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_918),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_R g953 ( 
.A(n_919),
.B(n_827),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_873),
.Y(n_954)
);

NAND2xp33_ASAP7_75t_L g955 ( 
.A(n_905),
.B(n_743),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_874),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_875),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_877),
.B(n_763),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_852),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_843),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_881),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_855),
.B(n_738),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_883),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_843),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_870),
.B(n_761),
.Y(n_965)
);

INVxp67_ASAP7_75t_L g966 ( 
.A(n_836),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_851),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_880),
.B(n_891),
.Y(n_968)
);

AOI22xp33_ASAP7_75t_L g969 ( 
.A1(n_840),
.A2(n_774),
.B1(n_802),
.B2(n_775),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_880),
.B(n_827),
.Y(n_970)
);

OR2x6_ASAP7_75t_L g971 ( 
.A(n_877),
.B(n_778),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_891),
.B(n_897),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_851),
.Y(n_973)
);

BUFx8_ASAP7_75t_SL g974 ( 
.A(n_910),
.Y(n_974)
);

NAND2xp33_ASAP7_75t_L g975 ( 
.A(n_911),
.B(n_743),
.Y(n_975)
);

NAND2xp33_ASAP7_75t_SL g976 ( 
.A(n_861),
.B(n_786),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_842),
.B(n_817),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_842),
.B(n_819),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_833),
.B(n_733),
.Y(n_979)
);

INVx2_ASAP7_75t_SL g980 ( 
.A(n_898),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_901),
.Y(n_981)
);

OR2x6_ASAP7_75t_L g982 ( 
.A(n_838),
.B(n_787),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_866),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_892),
.B(n_799),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_890),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_863),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_893),
.B(n_787),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_846),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_L g989 ( 
.A1(n_840),
.A2(n_692),
.B1(n_743),
.B2(n_672),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_SL g990 ( 
.A1(n_840),
.A2(n_673),
.B1(n_768),
.B2(n_665),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_870),
.B(n_768),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_914),
.B(n_787),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_914),
.B(n_721),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_878),
.B(n_758),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_894),
.B(n_723),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_863),
.Y(n_996)
);

BUFx8_ASAP7_75t_SL g997 ( 
.A(n_901),
.Y(n_997)
);

INVxp33_ASAP7_75t_L g998 ( 
.A(n_907),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_898),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_908),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_831),
.B(n_780),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_832),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_839),
.B(n_682),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_920),
.B(n_841),
.Y(n_1004)
);

INVx5_ASAP7_75t_L g1005 ( 
.A(n_852),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_858),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_898),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_859),
.Y(n_1008)
);

BUFx10_ASAP7_75t_L g1009 ( 
.A(n_895),
.Y(n_1009)
);

AND2x6_ASAP7_75t_L g1010 ( 
.A(n_878),
.B(n_595),
.Y(n_1010)
);

INVxp67_ASAP7_75t_SL g1011 ( 
.A(n_852),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_853),
.B(n_857),
.Y(n_1012)
);

OAI22xp33_ASAP7_75t_SL g1013 ( 
.A1(n_845),
.A2(n_770),
.B1(n_793),
.B2(n_758),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_872),
.B(n_724),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_864),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_912),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_889),
.B(n_725),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_849),
.B(n_656),
.Y(n_1018)
);

INVx4_ASAP7_75t_L g1019 ( 
.A(n_852),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_953),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_959),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_959),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_991),
.B(n_932),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_952),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_991),
.B(n_864),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_977),
.A2(n_849),
.B1(n_899),
.B2(n_896),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_945),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_979),
.B(n_879),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_924),
.B(n_932),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_951),
.Y(n_1030)
);

OR2x2_ASAP7_75t_L g1031 ( 
.A(n_968),
.B(n_757),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_921),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_944),
.B(n_854),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_925),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_936),
.B(n_854),
.Y(n_1035)
);

INVxp67_ASAP7_75t_L g1036 ( 
.A(n_935),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_SL g1037 ( 
.A(n_936),
.B(n_546),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_923),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_940),
.B(n_879),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_940),
.B(n_885),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_928),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_931),
.Y(n_1042)
);

AND2x6_ASAP7_75t_SL g1043 ( 
.A(n_970),
.B(n_691),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_962),
.B(n_816),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_1000),
.B(n_885),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_972),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_990),
.A2(n_969),
.B1(n_978),
.B2(n_954),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_990),
.A2(n_816),
.B1(n_904),
.B2(n_886),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_956),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_927),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_948),
.B(n_854),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_957),
.Y(n_1052)
);

NOR2x1p5_ASAP7_75t_L g1053 ( 
.A(n_958),
.B(n_671),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_989),
.A2(n_887),
.B1(n_884),
.B2(n_868),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1018),
.B(n_868),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_930),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1018),
.B(n_770),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_942),
.B(n_909),
.Y(n_1058)
);

AOI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_926),
.A2(n_916),
.B1(n_917),
.B2(n_913),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_947),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_966),
.B(n_958),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_994),
.B(n_854),
.Y(n_1062)
);

INVxp67_ASAP7_75t_L g1063 ( 
.A(n_934),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_961),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1012),
.B(n_966),
.Y(n_1065)
);

NAND2xp33_ASAP7_75t_L g1066 ( 
.A(n_963),
.B(n_862),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_998),
.B(n_862),
.Y(n_1067)
);

OR2x6_ASAP7_75t_L g1068 ( 
.A(n_971),
.B(n_902),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_984),
.A2(n_862),
.B1(n_909),
.B2(n_867),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_1001),
.B(n_862),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_959),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_985),
.B(n_793),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_922),
.B(n_866),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_949),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1002),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_967),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_922),
.B(n_867),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_973),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_946),
.B(n_812),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_981),
.B(n_900),
.Y(n_1080)
);

NAND2xp33_ASAP7_75t_L g1081 ( 
.A(n_1005),
.B(n_915),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_965),
.B(n_812),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_SL g1083 ( 
.A(n_971),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_1003),
.B(n_684),
.Y(n_1084)
);

OR2x2_ASAP7_75t_L g1085 ( 
.A(n_933),
.B(n_726),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_941),
.B(n_900),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_988),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_965),
.B(n_728),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_986),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_996),
.Y(n_1090)
);

NAND2xp33_ASAP7_75t_L g1091 ( 
.A(n_1005),
.B(n_915),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_993),
.B(n_915),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_1006),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_994),
.B(n_915),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_976),
.A2(n_743),
.B1(n_734),
.B2(n_736),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1013),
.B(n_856),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1029),
.B(n_982),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_1044),
.B(n_974),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1093),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1047),
.A2(n_1008),
.B1(n_939),
.B2(n_1016),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_1020),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1084),
.B(n_982),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1047),
.B(n_982),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1023),
.B(n_1013),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1023),
.B(n_1015),
.Y(n_1105)
);

INVxp67_ASAP7_75t_L g1106 ( 
.A(n_1046),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1057),
.B(n_1015),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1076),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_1024),
.B(n_927),
.Y(n_1109)
);

OR2x2_ASAP7_75t_L g1110 ( 
.A(n_1031),
.B(n_971),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1036),
.B(n_1004),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1032),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_1050),
.Y(n_1113)
);

NOR2xp67_ASAP7_75t_L g1114 ( 
.A(n_1079),
.B(n_941),
.Y(n_1114)
);

INVx1_ASAP7_75t_SL g1115 ( 
.A(n_1027),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1065),
.B(n_987),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_1053),
.B(n_999),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1070),
.B(n_1072),
.Y(n_1118)
);

BUFx2_ASAP7_75t_L g1119 ( 
.A(n_1030),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_1061),
.Y(n_1120)
);

INVx4_ASAP7_75t_L g1121 ( 
.A(n_1083),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1021),
.Y(n_1122)
);

INVx5_ASAP7_75t_L g1123 ( 
.A(n_1021),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_1028),
.B(n_1005),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1034),
.B(n_980),
.Y(n_1125)
);

BUFx4f_ASAP7_75t_SL g1126 ( 
.A(n_1085),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_1058),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_1021),
.Y(n_1128)
);

OR2x6_ASAP7_75t_L g1129 ( 
.A(n_1063),
.B(n_1007),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_1037),
.B(n_1005),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1041),
.B(n_992),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_1022),
.Y(n_1132)
);

INVxp67_ASAP7_75t_L g1133 ( 
.A(n_1083),
.Y(n_1133)
);

NAND2x1p5_ASAP7_75t_L g1134 ( 
.A(n_1022),
.B(n_1019),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1042),
.B(n_929),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1049),
.B(n_929),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_1022),
.Y(n_1137)
);

CKINVDCx8_ASAP7_75t_R g1138 ( 
.A(n_1043),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1071),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1052),
.B(n_1064),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1078),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_1071),
.Y(n_1142)
);

AND2x4_ASAP7_75t_SL g1143 ( 
.A(n_1068),
.B(n_1009),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_SL g1144 ( 
.A1(n_1075),
.A2(n_1087),
.B1(n_1067),
.B2(n_1037),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1045),
.B(n_997),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_1068),
.B(n_1019),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1082),
.B(n_937),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1035),
.A2(n_975),
.B(n_955),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_1071),
.B(n_960),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1088),
.B(n_937),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1096),
.A2(n_950),
.B(n_943),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1048),
.B(n_938),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1089),
.A2(n_1090),
.B1(n_1056),
.B2(n_1060),
.Y(n_1153)
);

AOI22xp33_ASAP7_75t_L g1154 ( 
.A1(n_1038),
.A2(n_1010),
.B1(n_938),
.B2(n_1014),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1095),
.A2(n_1080),
.B1(n_1026),
.B2(n_1051),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1074),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1055),
.Y(n_1157)
);

INVxp33_ASAP7_75t_L g1158 ( 
.A(n_1058),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1039),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1040),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1068),
.Y(n_1161)
);

OR2x2_ASAP7_75t_L g1162 ( 
.A(n_1033),
.B(n_960),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1054),
.A2(n_1010),
.B1(n_1017),
.B2(n_1009),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_SL g1164 ( 
.A1(n_1094),
.A2(n_1010),
.B1(n_635),
.B2(n_637),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1073),
.A2(n_964),
.B(n_983),
.C(n_731),
.Y(n_1165)
);

INVx4_ASAP7_75t_L g1166 ( 
.A(n_1081),
.Y(n_1166)
);

AOI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1096),
.A2(n_950),
.B(n_943),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1069),
.B(n_964),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1118),
.B(n_1062),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_1166),
.B(n_1062),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1105),
.B(n_1025),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1166),
.B(n_1094),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1111),
.B(n_1025),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_1097),
.B(n_1092),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1104),
.B(n_1106),
.Y(n_1175)
);

OR2x2_ASAP7_75t_L g1176 ( 
.A(n_1110),
.B(n_1077),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1107),
.B(n_1059),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1115),
.B(n_1123),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1117),
.B(n_1158),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1123),
.B(n_983),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1123),
.B(n_1086),
.Y(n_1181)
);

NAND2xp33_ASAP7_75t_SL g1182 ( 
.A(n_1101),
.B(n_634),
.Y(n_1182)
);

NAND2xp33_ASAP7_75t_R g1183 ( 
.A(n_1119),
.B(n_465),
.Y(n_1183)
);

NAND2xp33_ASAP7_75t_R g1184 ( 
.A(n_1098),
.B(n_468),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_1144),
.B(n_1011),
.Y(n_1185)
);

NAND2xp33_ASAP7_75t_SL g1186 ( 
.A(n_1116),
.B(n_995),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1117),
.B(n_756),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_1144),
.B(n_1114),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_1114),
.B(n_900),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1100),
.B(n_900),
.Y(n_1190)
);

NAND2x1p5_ASAP7_75t_L g1191 ( 
.A(n_1121),
.B(n_903),
.Y(n_1191)
);

NAND2xp33_ASAP7_75t_SL g1192 ( 
.A(n_1113),
.B(n_1091),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1161),
.B(n_1010),
.Y(n_1193)
);

NAND2xp33_ASAP7_75t_SL g1194 ( 
.A(n_1140),
.B(n_903),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1159),
.B(n_1066),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_1146),
.B(n_1120),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1146),
.B(n_906),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1103),
.B(n_1102),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1122),
.B(n_906),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_1122),
.B(n_1128),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1122),
.B(n_906),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1121),
.B(n_903),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1128),
.B(n_906),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1128),
.B(n_903),
.Y(n_1204)
);

NAND2xp33_ASAP7_75t_SL g1205 ( 
.A(n_1125),
.B(n_470),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1137),
.B(n_1164),
.Y(n_1206)
);

NAND2xp33_ASAP7_75t_SL g1207 ( 
.A(n_1131),
.B(n_477),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1137),
.B(n_767),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_SL g1209 ( 
.A(n_1137),
.B(n_767),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1160),
.B(n_752),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1145),
.B(n_767),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1157),
.B(n_752),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_1155),
.B(n_767),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_1155),
.B(n_614),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1127),
.B(n_1138),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_1132),
.B(n_617),
.Y(n_1216)
);

NAND2xp33_ASAP7_75t_SL g1217 ( 
.A(n_1162),
.B(n_480),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1132),
.B(n_1139),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_1139),
.B(n_618),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_1142),
.B(n_621),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_1142),
.B(n_628),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1126),
.B(n_638),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1143),
.B(n_594),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1133),
.B(n_123),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1109),
.B(n_125),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1163),
.B(n_636),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1129),
.B(n_126),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1112),
.B(n_632),
.Y(n_1228)
);

NAND2xp33_ASAP7_75t_SL g1229 ( 
.A(n_1149),
.B(n_481),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1099),
.B(n_0),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1147),
.B(n_482),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1135),
.B(n_631),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1129),
.B(n_127),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1136),
.B(n_627),
.Y(n_1234)
);

NAND2xp33_ASAP7_75t_SL g1235 ( 
.A(n_1130),
.B(n_487),
.Y(n_1235)
);

NAND2xp33_ASAP7_75t_SL g1236 ( 
.A(n_1168),
.B(n_489),
.Y(n_1236)
);

NAND2xp33_ASAP7_75t_SL g1237 ( 
.A(n_1150),
.B(n_491),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1134),
.B(n_626),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1179),
.B(n_1215),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1173),
.B(n_1156),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1202),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1177),
.B(n_1124),
.Y(n_1242)
);

INVx4_ASAP7_75t_L g1243 ( 
.A(n_1227),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1214),
.A2(n_1152),
.B1(n_1154),
.B2(n_1165),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1202),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1195),
.B(n_1151),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1175),
.B(n_1108),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1171),
.B(n_1141),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1230),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_SL g1250 ( 
.A1(n_1225),
.A2(n_543),
.B1(n_608),
.B2(n_597),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1176),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_1182),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1198),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1217),
.A2(n_1153),
.B1(n_597),
.B2(n_608),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1169),
.B(n_1167),
.Y(n_1255)
);

NOR2x1_ASAP7_75t_L g1256 ( 
.A(n_1211),
.B(n_1148),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1196),
.B(n_1),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1178),
.B(n_2),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1210),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1212),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1174),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1172),
.Y(n_1262)
);

INVx4_ASAP7_75t_L g1263 ( 
.A(n_1227),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_1183),
.Y(n_1264)
);

INVxp67_ASAP7_75t_L g1265 ( 
.A(n_1187),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1170),
.Y(n_1266)
);

BUFx8_ASAP7_75t_SL g1267 ( 
.A(n_1233),
.Y(n_1267)
);

CKINVDCx16_ASAP7_75t_R g1268 ( 
.A(n_1184),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1225),
.Y(n_1269)
);

NAND2x1p5_ASAP7_75t_L g1270 ( 
.A(n_1233),
.B(n_128),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1222),
.Y(n_1271)
);

NAND2x1p5_ASAP7_75t_L g1272 ( 
.A(n_1197),
.B(n_129),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1224),
.B(n_1223),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1224),
.B(n_2),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1223),
.B(n_3),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1188),
.B(n_604),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1200),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1185),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1218),
.Y(n_1279)
);

AND2x2_ASAP7_75t_SL g1280 ( 
.A(n_1193),
.B(n_3),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1206),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1193),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1228),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1213),
.B(n_4),
.Y(n_1284)
);

AOI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1186),
.A2(n_499),
.B1(n_496),
.B2(n_498),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1216),
.B(n_4),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1199),
.Y(n_1287)
);

NAND2x1p5_ASAP7_75t_L g1288 ( 
.A(n_1180),
.B(n_131),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_1191),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1190),
.A2(n_503),
.B(n_493),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1205),
.B(n_6),
.Y(n_1291)
);

BUFx8_ASAP7_75t_L g1292 ( 
.A(n_1192),
.Y(n_1292)
);

AND2x4_ASAP7_75t_SL g1293 ( 
.A(n_1235),
.B(n_134),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1201),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1219),
.B(n_6),
.Y(n_1295)
);

AOI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1236),
.A2(n_509),
.B1(n_510),
.B2(n_504),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1226),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1220),
.B(n_7),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1181),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_SL g1300 ( 
.A1(n_1207),
.A2(n_11),
.B1(n_8),
.B2(n_10),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1231),
.B(n_12),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1229),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1203),
.Y(n_1303)
);

AND2x4_ASAP7_75t_SL g1304 ( 
.A(n_1221),
.B(n_136),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1238),
.B(n_12),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1194),
.A2(n_514),
.B(n_511),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1204),
.B(n_1189),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1232),
.B(n_13),
.Y(n_1308)
);

AND3x1_ASAP7_75t_SL g1309 ( 
.A(n_1237),
.B(n_13),
.C(n_14),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1234),
.B(n_1208),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1209),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1179),
.B(n_15),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_1215),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1215),
.Y(n_1314)
);

CKINVDCx16_ASAP7_75t_R g1315 ( 
.A(n_1183),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_1215),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1210),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1177),
.B(n_522),
.Y(n_1318)
);

CKINVDCx12_ASAP7_75t_R g1319 ( 
.A(n_1215),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_1183),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1299),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1253),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1251),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1256),
.A2(n_139),
.B(n_137),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1246),
.B(n_15),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1255),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1313),
.Y(n_1327)
);

NAND2x1p5_ASAP7_75t_L g1328 ( 
.A(n_1243),
.B(n_140),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_1281),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1307),
.A2(n_143),
.B(n_142),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1299),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1307),
.A2(n_145),
.B(n_144),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1261),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1243),
.B(n_146),
.Y(n_1334)
);

BUFx2_ASAP7_75t_L g1335 ( 
.A(n_1263),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1265),
.B(n_16),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1247),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_SL g1338 ( 
.A1(n_1263),
.A2(n_1285),
.B(n_1284),
.Y(n_1338)
);

BUFx2_ASAP7_75t_L g1339 ( 
.A(n_1292),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_1267),
.Y(n_1340)
);

AO21x2_ASAP7_75t_L g1341 ( 
.A1(n_1278),
.A2(n_534),
.B(n_533),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1262),
.Y(n_1342)
);

AO21x2_ASAP7_75t_L g1343 ( 
.A1(n_1242),
.A2(n_544),
.B(n_540),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1284),
.A2(n_148),
.B(n_147),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1266),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_1241),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1241),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1239),
.B(n_16),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1260),
.Y(n_1349)
);

OAI21xp33_ASAP7_75t_SL g1350 ( 
.A1(n_1285),
.A2(n_17),
.B(n_18),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1259),
.Y(n_1351)
);

AO21x2_ASAP7_75t_L g1352 ( 
.A1(n_1249),
.A2(n_550),
.B(n_545),
.Y(n_1352)
);

AO21x2_ASAP7_75t_L g1353 ( 
.A1(n_1248),
.A2(n_1244),
.B(n_1311),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1271),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_1241),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1303),
.Y(n_1356)
);

INVx1_ASAP7_75t_SL g1357 ( 
.A(n_1245),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1292),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1245),
.B(n_149),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1287),
.A2(n_151),
.B(n_150),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1314),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1294),
.A2(n_153),
.B(n_152),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1316),
.B(n_155),
.Y(n_1363)
);

INVx6_ASAP7_75t_L g1364 ( 
.A(n_1289),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1317),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1277),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1279),
.Y(n_1367)
);

BUFx2_ASAP7_75t_SL g1368 ( 
.A(n_1252),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1240),
.Y(n_1369)
);

INVx6_ASAP7_75t_SL g1370 ( 
.A(n_1319),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1269),
.B(n_17),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1282),
.Y(n_1372)
);

INVx1_ASAP7_75t_SL g1373 ( 
.A(n_1273),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_1264),
.Y(n_1374)
);

BUFx2_ASAP7_75t_L g1375 ( 
.A(n_1283),
.Y(n_1375)
);

BUFx5_ASAP7_75t_L g1376 ( 
.A(n_1280),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1289),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1312),
.Y(n_1378)
);

AO21x2_ASAP7_75t_L g1379 ( 
.A1(n_1244),
.A2(n_555),
.B(n_551),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1257),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1276),
.A2(n_1297),
.B(n_1250),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1289),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1258),
.Y(n_1383)
);

BUFx8_ASAP7_75t_L g1384 ( 
.A(n_1275),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1274),
.Y(n_1385)
);

AND2x4_ASAP7_75t_L g1386 ( 
.A(n_1286),
.B(n_157),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1276),
.Y(n_1387)
);

NAND2x1p5_ASAP7_75t_L g1388 ( 
.A(n_1310),
.B(n_158),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1272),
.A2(n_161),
.B(n_160),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1288),
.A2(n_1270),
.B(n_1308),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1301),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_1302),
.Y(n_1392)
);

AO21x2_ASAP7_75t_L g1393 ( 
.A1(n_1318),
.A2(n_559),
.B(n_557),
.Y(n_1393)
);

AOI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1306),
.A2(n_562),
.B(n_560),
.Y(n_1394)
);

OA21x2_ASAP7_75t_L g1395 ( 
.A1(n_1254),
.A2(n_570),
.B(n_564),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1297),
.A2(n_165),
.B(n_162),
.Y(n_1396)
);

INVx3_ASAP7_75t_SL g1397 ( 
.A(n_1320),
.Y(n_1397)
);

OAI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1291),
.A2(n_1296),
.B(n_1290),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1305),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_1295),
.B(n_166),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1367),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1398),
.A2(n_1300),
.B1(n_1296),
.B2(n_1268),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1379),
.A2(n_1300),
.B1(n_1315),
.B2(n_1298),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1366),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1398),
.A2(n_1293),
.B1(n_1309),
.B2(n_1304),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1323),
.Y(n_1406)
);

INVx2_ASAP7_75t_SL g1407 ( 
.A(n_1327),
.Y(n_1407)
);

OAI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1381),
.A2(n_575),
.B1(n_582),
.B2(n_572),
.Y(n_1408)
);

CKINVDCx11_ASAP7_75t_R g1409 ( 
.A(n_1340),
.Y(n_1409)
);

OAI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1381),
.A2(n_585),
.B1(n_586),
.B2(n_584),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1322),
.Y(n_1411)
);

BUFx12f_ASAP7_75t_L g1412 ( 
.A(n_1374),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1325),
.A2(n_598),
.B1(n_600),
.B2(n_592),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_1321),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1379),
.A2(n_624),
.B1(n_606),
.B2(n_610),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1325),
.A2(n_613),
.B1(n_622),
.B2(n_601),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1333),
.Y(n_1417)
);

AOI22xp5_ASAP7_75t_SL g1418 ( 
.A1(n_1340),
.A2(n_1376),
.B1(n_1361),
.B2(n_1368),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1392),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1352),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_1420)
);

CKINVDCx6p67_ASAP7_75t_R g1421 ( 
.A(n_1397),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1342),
.Y(n_1422)
);

INVx1_ASAP7_75t_SL g1423 ( 
.A(n_1397),
.Y(n_1423)
);

INVx1_ASAP7_75t_SL g1424 ( 
.A(n_1392),
.Y(n_1424)
);

INVx6_ASAP7_75t_L g1425 ( 
.A(n_1384),
.Y(n_1425)
);

BUFx8_ASAP7_75t_SL g1426 ( 
.A(n_1339),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_SL g1427 ( 
.A1(n_1376),
.A2(n_1350),
.B1(n_1352),
.B2(n_1395),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1358),
.Y(n_1428)
);

BUFx3_ASAP7_75t_L g1429 ( 
.A(n_1374),
.Y(n_1429)
);

INVx2_ASAP7_75t_SL g1430 ( 
.A(n_1364),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1370),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1345),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1370),
.Y(n_1433)
);

BUFx4f_ASAP7_75t_SL g1434 ( 
.A(n_1384),
.Y(n_1434)
);

INVx6_ASAP7_75t_L g1435 ( 
.A(n_1346),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1376),
.A2(n_22),
.B1(n_19),
.B2(n_20),
.Y(n_1436)
);

INVx6_ASAP7_75t_L g1437 ( 
.A(n_1346),
.Y(n_1437)
);

BUFx8_ASAP7_75t_L g1438 ( 
.A(n_1348),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1321),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_SL g1440 ( 
.A1(n_1376),
.A2(n_26),
.B1(n_23),
.B2(n_24),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1345),
.Y(n_1441)
);

OAI22xp33_ASAP7_75t_SL g1442 ( 
.A1(n_1387),
.A2(n_26),
.B1(n_23),
.B2(n_24),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1376),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_1443)
);

BUFx12f_ASAP7_75t_L g1444 ( 
.A(n_1354),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_SL g1445 ( 
.A1(n_1350),
.A2(n_30),
.B1(n_27),
.B2(n_28),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1356),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1388),
.A2(n_33),
.B1(n_30),
.B2(n_32),
.Y(n_1447)
);

INVx3_ASAP7_75t_SL g1448 ( 
.A(n_1354),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_SL g1449 ( 
.A1(n_1395),
.A2(n_36),
.B1(n_33),
.B2(n_34),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1341),
.A2(n_38),
.B1(n_34),
.B2(n_37),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1356),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1351),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1341),
.A2(n_1399),
.B1(n_1378),
.B2(n_1383),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1369),
.B(n_39),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1375),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_L g1456 ( 
.A(n_1385),
.B(n_1336),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1349),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_SL g1458 ( 
.A1(n_1338),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1365),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_1459)
);

OAI22xp33_ASAP7_75t_SL g1460 ( 
.A1(n_1391),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1380),
.B(n_44),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_SL g1462 ( 
.A1(n_1380),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_1462)
);

AOI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1373),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1329),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_SL g1465 ( 
.A1(n_1353),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_1465)
);

BUFx12f_ASAP7_75t_L g1466 ( 
.A(n_1363),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1373),
.B(n_50),
.Y(n_1467)
);

OAI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1388),
.A2(n_1328),
.B1(n_1329),
.B2(n_1371),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_1346),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1328),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1357),
.B(n_52),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_SL g1472 ( 
.A1(n_1353),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1326),
.Y(n_1473)
);

CKINVDCx6p67_ASAP7_75t_R g1474 ( 
.A(n_1363),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_SL g1475 ( 
.A1(n_1386),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1326),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1372),
.Y(n_1477)
);

AOI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1390),
.A2(n_57),
.B(n_58),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1343),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1343),
.A2(n_62),
.B1(n_59),
.B2(n_61),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1473),
.Y(n_1481)
);

CKINVDCx6p67_ASAP7_75t_R g1482 ( 
.A(n_1409),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1455),
.B(n_1335),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1404),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_1469),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1402),
.A2(n_1371),
.B(n_1334),
.Y(n_1486)
);

AOI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1468),
.A2(n_1334),
.B(n_1396),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1476),
.Y(n_1488)
);

AO31x2_ASAP7_75t_L g1489 ( 
.A1(n_1405),
.A2(n_1337),
.A3(n_1357),
.B(n_1331),
.Y(n_1489)
);

OA21x2_ASAP7_75t_L g1490 ( 
.A1(n_1453),
.A2(n_1332),
.B(n_1330),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1422),
.Y(n_1491)
);

A2O1A1Ixp33_ASAP7_75t_L g1492 ( 
.A1(n_1403),
.A2(n_1386),
.B(n_1400),
.C(n_1389),
.Y(n_1492)
);

OAI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1463),
.A2(n_1331),
.B1(n_1400),
.B2(n_1382),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1423),
.B(n_1393),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1451),
.B(n_1377),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1445),
.A2(n_1359),
.B1(n_1364),
.B2(n_1377),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1432),
.Y(n_1497)
);

BUFx2_ASAP7_75t_R g1498 ( 
.A(n_1426),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1478),
.A2(n_1344),
.B(n_1360),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1441),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1401),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1464),
.B(n_1382),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1446),
.B(n_1347),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1408),
.A2(n_1324),
.B(n_1359),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1411),
.B(n_1347),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1417),
.Y(n_1506)
);

A2O1A1Ixp33_ASAP7_75t_L g1507 ( 
.A1(n_1440),
.A2(n_1362),
.B(n_1393),
.C(n_1355),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1477),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1418),
.B(n_1347),
.Y(n_1509)
);

AOI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1410),
.A2(n_1355),
.B(n_1364),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1456),
.B(n_1457),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1414),
.Y(n_1512)
);

NAND3xp33_ASAP7_75t_L g1513 ( 
.A(n_1465),
.B(n_1355),
.C(n_1394),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1406),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1452),
.Y(n_1515)
);

AOI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1440),
.A2(n_61),
.B(n_63),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1448),
.B(n_63),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1418),
.B(n_64),
.Y(n_1518)
);

OR2x6_ASAP7_75t_L g1519 ( 
.A(n_1466),
.B(n_65),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1424),
.B(n_65),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1419),
.B(n_66),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1461),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1414),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1467),
.A2(n_66),
.B(n_67),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1439),
.B(n_67),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1439),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1454),
.Y(n_1527)
);

INVx1_ASAP7_75t_SL g1528 ( 
.A(n_1428),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_SL g1529 ( 
.A1(n_1442),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_1529)
);

INVx5_ASAP7_75t_SL g1530 ( 
.A(n_1421),
.Y(n_1530)
);

AOI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1415),
.A2(n_69),
.B(n_70),
.Y(n_1531)
);

OAI221xp5_ASAP7_75t_SL g1532 ( 
.A1(n_1463),
.A2(n_1443),
.B1(n_1436),
.B2(n_1475),
.C(n_1420),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1412),
.Y(n_1533)
);

OAI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1472),
.A2(n_71),
.B(n_72),
.Y(n_1534)
);

A2O1A1Ixp33_ASAP7_75t_L g1535 ( 
.A1(n_1427),
.A2(n_75),
.B(n_72),
.C(n_74),
.Y(n_1535)
);

INVx8_ASAP7_75t_L g1536 ( 
.A(n_1444),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1471),
.B(n_75),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1516),
.A2(n_1449),
.B1(n_1450),
.B2(n_1447),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1511),
.B(n_1407),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1534),
.A2(n_1442),
.B1(n_1460),
.B2(n_1479),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1497),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1513),
.A2(n_1460),
.B1(n_1480),
.B2(n_1470),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_SL g1543 ( 
.A1(n_1519),
.A2(n_1434),
.B1(n_1425),
.B2(n_1433),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1483),
.B(n_1429),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1532),
.A2(n_1458),
.B1(n_1462),
.B2(n_1474),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_SL g1546 ( 
.A1(n_1518),
.A2(n_1438),
.B1(n_1425),
.B2(n_1431),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1529),
.A2(n_1459),
.B1(n_1416),
.B2(n_1413),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1482),
.Y(n_1548)
);

AO31x2_ASAP7_75t_L g1549 ( 
.A1(n_1494),
.A2(n_1430),
.A3(n_1437),
.B(n_1435),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_1498),
.B(n_1438),
.Y(n_1550)
);

INVx4_ASAP7_75t_L g1551 ( 
.A(n_1536),
.Y(n_1551)
);

OAI21x1_ASAP7_75t_L g1552 ( 
.A1(n_1487),
.A2(n_1437),
.B(n_1435),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1495),
.B(n_1469),
.Y(n_1553)
);

AOI221xp5_ASAP7_75t_L g1554 ( 
.A1(n_1535),
.A2(n_1469),
.B1(n_79),
.B2(n_76),
.C(n_78),
.Y(n_1554)
);

AOI221xp5_ASAP7_75t_L g1555 ( 
.A1(n_1531),
.A2(n_80),
.B1(n_76),
.B2(n_78),
.C(n_81),
.Y(n_1555)
);

OAI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1486),
.A2(n_84),
.B1(n_80),
.B2(n_81),
.Y(n_1556)
);

A2O1A1Ixp33_ASAP7_75t_L g1557 ( 
.A1(n_1492),
.A2(n_87),
.B(n_85),
.C(n_86),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1523),
.B(n_85),
.Y(n_1558)
);

OAI221xp5_ASAP7_75t_L g1559 ( 
.A1(n_1507),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.C(n_90),
.Y(n_1559)
);

BUFx2_ASAP7_75t_L g1560 ( 
.A(n_1512),
.Y(n_1560)
);

OA21x2_ASAP7_75t_L g1561 ( 
.A1(n_1497),
.A2(n_88),
.B(n_89),
.Y(n_1561)
);

AOI21xp33_ASAP7_75t_SL g1562 ( 
.A1(n_1536),
.A2(n_90),
.B(n_92),
.Y(n_1562)
);

AOI221xp5_ASAP7_75t_L g1563 ( 
.A1(n_1527),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.C(n_95),
.Y(n_1563)
);

OAI221xp5_ASAP7_75t_L g1564 ( 
.A1(n_1527),
.A2(n_96),
.B1(n_93),
.B2(n_94),
.C(n_97),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1490),
.A2(n_1522),
.B1(n_1493),
.B2(n_1496),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1509),
.B(n_98),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1490),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1528),
.B(n_99),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1526),
.B(n_100),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1481),
.B(n_101),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1500),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1504),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_SL g1573 ( 
.A1(n_1537),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_1573)
);

OAI221xp5_ASAP7_75t_L g1574 ( 
.A1(n_1519),
.A2(n_104),
.B1(n_106),
.B2(n_108),
.C(n_109),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1514),
.A2(n_110),
.B1(n_106),
.B2(n_109),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_SL g1576 ( 
.A1(n_1517),
.A2(n_112),
.B1(n_110),
.B2(n_111),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1484),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1500),
.B(n_113),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1491),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_1579)
);

BUFx12f_ASAP7_75t_L g1580 ( 
.A(n_1533),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1525),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1521),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_1520),
.Y(n_1583)
);

BUFx3_ASAP7_75t_L g1584 ( 
.A(n_1580),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1541),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1552),
.B(n_1489),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1561),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1560),
.B(n_1489),
.Y(n_1588)
);

AND2x2_ASAP7_75t_SL g1589 ( 
.A(n_1565),
.B(n_1566),
.Y(n_1589)
);

INVxp67_ASAP7_75t_L g1590 ( 
.A(n_1578),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1561),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1571),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1549),
.B(n_1489),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1549),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1549),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1578),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1570),
.B(n_1481),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1539),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1558),
.Y(n_1599)
);

INVxp67_ASAP7_75t_SL g1600 ( 
.A(n_1583),
.Y(n_1600)
);

NAND2x1_ASAP7_75t_L g1601 ( 
.A(n_1544),
.B(n_1553),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1582),
.B(n_1488),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1569),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1566),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1581),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1567),
.B(n_1503),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1546),
.B(n_1506),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1568),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1581),
.B(n_1506),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1559),
.Y(n_1610)
);

BUFx6f_ASAP7_75t_L g1611 ( 
.A(n_1551),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1564),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1557),
.B(n_1502),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1556),
.Y(n_1614)
);

OAI221xp5_ASAP7_75t_L g1615 ( 
.A1(n_1605),
.A2(n_1540),
.B1(n_1542),
.B2(n_1545),
.C(n_1572),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1596),
.Y(n_1616)
);

OA21x2_ASAP7_75t_L g1617 ( 
.A1(n_1587),
.A2(n_1524),
.B(n_1499),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1585),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1587),
.Y(n_1619)
);

OAI21x1_ASAP7_75t_SL g1620 ( 
.A1(n_1609),
.A2(n_1551),
.B(n_1545),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1591),
.Y(n_1621)
);

OAI211xp5_ASAP7_75t_L g1622 ( 
.A1(n_1605),
.A2(n_1576),
.B(n_1562),
.C(n_1573),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1591),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1597),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1592),
.Y(n_1625)
);

AOI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1612),
.A2(n_1589),
.B(n_1613),
.Y(n_1626)
);

NAND3xp33_ASAP7_75t_L g1627 ( 
.A(n_1612),
.B(n_1554),
.C(n_1555),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1592),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1611),
.Y(n_1629)
);

OR2x2_ASAP7_75t_SL g1630 ( 
.A(n_1611),
.B(n_1543),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1590),
.Y(n_1631)
);

INVxp67_ASAP7_75t_L g1632 ( 
.A(n_1600),
.Y(n_1632)
);

OA21x2_ASAP7_75t_L g1633 ( 
.A1(n_1594),
.A2(n_1510),
.B(n_1538),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1589),
.A2(n_1574),
.B1(n_1563),
.B2(n_1575),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1598),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1611),
.B(n_1548),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1602),
.Y(n_1637)
);

NOR2x1_ASAP7_75t_SL g1638 ( 
.A(n_1588),
.B(n_1485),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1602),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1610),
.A2(n_1550),
.B(n_1547),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1607),
.B(n_1530),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1619),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1631),
.B(n_1614),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1624),
.B(n_1608),
.Y(n_1644)
);

OAI31xp33_ASAP7_75t_L g1645 ( 
.A1(n_1626),
.A2(n_1586),
.A3(n_1593),
.B(n_1606),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1641),
.B(n_1607),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1619),
.Y(n_1647)
);

INVx5_ASAP7_75t_SL g1648 ( 
.A(n_1630),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1616),
.B(n_1599),
.Y(n_1649)
);

BUFx12f_ASAP7_75t_L g1650 ( 
.A(n_1641),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1632),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1629),
.B(n_1611),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1623),
.Y(n_1653)
);

NOR3xp33_ASAP7_75t_L g1654 ( 
.A(n_1622),
.B(n_1547),
.C(n_1584),
.Y(n_1654)
);

INVxp67_ASAP7_75t_L g1655 ( 
.A(n_1627),
.Y(n_1655)
);

INVxp33_ASAP7_75t_L g1656 ( 
.A(n_1636),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1621),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1637),
.B(n_1601),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1639),
.B(n_1530),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1646),
.B(n_1636),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1655),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1651),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1644),
.B(n_1635),
.Y(n_1663)
);

NOR2x1_ASAP7_75t_SL g1664 ( 
.A(n_1650),
.B(n_1635),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1646),
.Y(n_1665)
);

NAND4xp25_ASAP7_75t_L g1666 ( 
.A(n_1654),
.B(n_1615),
.C(n_1640),
.D(n_1634),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1659),
.B(n_1584),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1655),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1651),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1656),
.B(n_1618),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1652),
.B(n_1638),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1653),
.Y(n_1672)
);

NAND4xp75_ASAP7_75t_L g1673 ( 
.A(n_1661),
.B(n_1645),
.C(n_1633),
.D(n_1648),
.Y(n_1673)
);

INVx1_ASAP7_75t_SL g1674 ( 
.A(n_1661),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1667),
.B(n_1656),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1668),
.B(n_1654),
.Y(n_1676)
);

BUFx3_ASAP7_75t_L g1677 ( 
.A(n_1660),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1668),
.B(n_1649),
.Y(n_1678)
);

AOI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1666),
.A2(n_1633),
.B1(n_1621),
.B2(n_1623),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1662),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1669),
.Y(n_1681)
);

XOR2x2_ASAP7_75t_L g1682 ( 
.A(n_1664),
.B(n_1633),
.Y(n_1682)
);

BUFx2_ASAP7_75t_L g1683 ( 
.A(n_1660),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1670),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1675),
.B(n_1665),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1674),
.B(n_1676),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1683),
.B(n_1652),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1677),
.B(n_1648),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1674),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1684),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1678),
.Y(n_1691)
);

NOR2xp67_ASAP7_75t_L g1692 ( 
.A(n_1678),
.B(n_1663),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1680),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1681),
.B(n_1648),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1679),
.B(n_1666),
.Y(n_1695)
);

OAI21xp33_ASAP7_75t_L g1696 ( 
.A1(n_1695),
.A2(n_1682),
.B(n_1672),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1689),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1695),
.A2(n_1673),
.B1(n_1671),
.B2(n_1649),
.Y(n_1698)
);

XOR2x2_ASAP7_75t_L g1699 ( 
.A(n_1686),
.B(n_1643),
.Y(n_1699)
);

OAI21xp33_ASAP7_75t_L g1700 ( 
.A1(n_1685),
.A2(n_1658),
.B(n_1671),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1687),
.B(n_1694),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1686),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1692),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1688),
.A2(n_1620),
.B1(n_1628),
.B2(n_1604),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1690),
.Y(n_1705)
);

OR2x6_ASAP7_75t_L g1706 ( 
.A(n_1693),
.B(n_1642),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1699),
.Y(n_1707)
);

OAI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1698),
.A2(n_1691),
.B1(n_1604),
.B2(n_1657),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1701),
.B(n_1603),
.Y(n_1709)
);

OAI311xp33_ASAP7_75t_L g1710 ( 
.A1(n_1696),
.A2(n_1577),
.A3(n_1579),
.B1(n_1647),
.C1(n_1617),
.Y(n_1710)
);

OAI322xp33_ASAP7_75t_L g1711 ( 
.A1(n_1702),
.A2(n_1625),
.A3(n_1595),
.B1(n_1594),
.B2(n_1617),
.C1(n_1505),
.C2(n_117),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1706),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1706),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1703),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1697),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1709),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1707),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1711),
.B(n_1700),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1712),
.Y(n_1719)
);

NOR2xp67_ASAP7_75t_L g1720 ( 
.A(n_1715),
.B(n_1705),
.Y(n_1720)
);

OAI21xp5_ASAP7_75t_SL g1721 ( 
.A1(n_1714),
.A2(n_1704),
.B(n_1586),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1713),
.B(n_1617),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1711),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1708),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1710),
.B(n_1625),
.Y(n_1725)
);

OAI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1707),
.A2(n_1586),
.B(n_1593),
.Y(n_1726)
);

OAI21xp5_ASAP7_75t_SL g1727 ( 
.A1(n_1707),
.A2(n_1593),
.B(n_1595),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1709),
.B(n_1485),
.Y(n_1728)
);

AOI211xp5_ASAP7_75t_L g1729 ( 
.A1(n_1718),
.A2(n_1485),
.B(n_120),
.C(n_118),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1720),
.B(n_1508),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1716),
.B(n_119),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_1724),
.B(n_1725),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1728),
.B(n_1717),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1719),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1723),
.B(n_119),
.Y(n_1735)
);

INVx2_ASAP7_75t_SL g1736 ( 
.A(n_1722),
.Y(n_1736)
);

OAI221xp5_ASAP7_75t_SL g1737 ( 
.A1(n_1721),
.A2(n_122),
.B1(n_1515),
.B2(n_1501),
.C(n_169),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1725),
.Y(n_1738)
);

AOI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1738),
.A2(n_1727),
.B1(n_1726),
.B2(n_170),
.Y(n_1739)
);

AOI222xp33_ASAP7_75t_L g1740 ( 
.A1(n_1732),
.A2(n_1736),
.B1(n_1735),
.B2(n_1734),
.C1(n_1730),
.C2(n_1733),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1729),
.B(n_167),
.Y(n_1741)
);

NOR3xp33_ASAP7_75t_L g1742 ( 
.A(n_1731),
.B(n_168),
.C(n_172),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1737),
.B(n_173),
.Y(n_1743)
);

OAI222xp33_ASAP7_75t_L g1744 ( 
.A1(n_1738),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.C1(n_177),
.C2(n_180),
.Y(n_1744)
);

AOI222xp33_ASAP7_75t_L g1745 ( 
.A1(n_1738),
.A2(n_181),
.B1(n_183),
.B2(n_187),
.C1(n_188),
.C2(n_189),
.Y(n_1745)
);

INVxp33_ASAP7_75t_L g1746 ( 
.A(n_1742),
.Y(n_1746)
);

AOI221xp5_ASAP7_75t_L g1747 ( 
.A1(n_1739),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.C(n_196),
.Y(n_1747)
);

OAI22x1_ASAP7_75t_L g1748 ( 
.A1(n_1741),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1740),
.Y(n_1749)
);

AOI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1743),
.A2(n_203),
.B1(n_200),
.B2(n_201),
.Y(n_1750)
);

A2O1A1Ixp33_ASAP7_75t_SL g1751 ( 
.A1(n_1744),
.A2(n_208),
.B(n_204),
.C(n_206),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1745),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1740),
.Y(n_1753)
);

A2O1A1Ixp33_ASAP7_75t_SL g1754 ( 
.A1(n_1739),
.A2(n_211),
.B(n_209),
.C(n_210),
.Y(n_1754)
);

AOI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1740),
.A2(n_464),
.B1(n_215),
.B2(n_212),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1740),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1741),
.Y(n_1757)
);

AOI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1749),
.A2(n_221),
.B1(n_214),
.B2(n_217),
.Y(n_1758)
);

AOI21xp33_ASAP7_75t_L g1759 ( 
.A1(n_1754),
.A2(n_222),
.B(n_223),
.Y(n_1759)
);

AOI211xp5_ASAP7_75t_L g1760 ( 
.A1(n_1753),
.A2(n_225),
.B(n_226),
.C(n_228),
.Y(n_1760)
);

OAI221xp5_ASAP7_75t_L g1761 ( 
.A1(n_1756),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.C(n_233),
.Y(n_1761)
);

OAI221xp5_ASAP7_75t_L g1762 ( 
.A1(n_1751),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.C(n_240),
.Y(n_1762)
);

OAI221xp5_ASAP7_75t_L g1763 ( 
.A1(n_1747),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.C(n_246),
.Y(n_1763)
);

O2A1O1Ixp5_ASAP7_75t_SL g1764 ( 
.A1(n_1752),
.A2(n_247),
.B(n_249),
.C(n_250),
.Y(n_1764)
);

OAI211xp5_ASAP7_75t_L g1765 ( 
.A1(n_1755),
.A2(n_1750),
.B(n_1757),
.C(n_1746),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1748),
.B(n_251),
.Y(n_1766)
);

AOI221x1_ASAP7_75t_L g1767 ( 
.A1(n_1749),
.A2(n_252),
.B1(n_253),
.B2(n_258),
.C(n_259),
.Y(n_1767)
);

OAI31xp33_ASAP7_75t_L g1768 ( 
.A1(n_1749),
.A2(n_261),
.A3(n_262),
.B(n_263),
.Y(n_1768)
);

INVx1_ASAP7_75t_SL g1769 ( 
.A(n_1749),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1749),
.B(n_264),
.Y(n_1770)
);

AOI322xp5_ASAP7_75t_L g1771 ( 
.A1(n_1749),
.A2(n_265),
.A3(n_266),
.B1(n_268),
.B2(n_270),
.C1(n_271),
.C2(n_272),
.Y(n_1771)
);

NAND3xp33_ASAP7_75t_SL g1772 ( 
.A(n_1749),
.B(n_273),
.C(n_274),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1769),
.B(n_275),
.Y(n_1773)
);

AOI221xp5_ASAP7_75t_L g1774 ( 
.A1(n_1759),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.C(n_279),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_L g1775 ( 
.A(n_1765),
.B(n_280),
.Y(n_1775)
);

O2A1O1Ixp33_ASAP7_75t_L g1776 ( 
.A1(n_1770),
.A2(n_281),
.B(n_282),
.C(n_283),
.Y(n_1776)
);

OAI221xp5_ASAP7_75t_L g1777 ( 
.A1(n_1762),
.A2(n_284),
.B1(n_287),
.B2(n_289),
.C(n_290),
.Y(n_1777)
);

OAI211xp5_ASAP7_75t_SL g1778 ( 
.A1(n_1768),
.A2(n_292),
.B(n_293),
.C(n_294),
.Y(n_1778)
);

INVxp67_ASAP7_75t_L g1779 ( 
.A(n_1766),
.Y(n_1779)
);

INVx1_ASAP7_75t_SL g1780 ( 
.A(n_1758),
.Y(n_1780)
);

NOR3xp33_ASAP7_75t_SL g1781 ( 
.A(n_1772),
.B(n_295),
.C(n_297),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1767),
.B(n_298),
.Y(n_1782)
);

AOI222xp33_ASAP7_75t_L g1783 ( 
.A1(n_1761),
.A2(n_299),
.B1(n_301),
.B2(n_303),
.C1(n_304),
.C2(n_305),
.Y(n_1783)
);

OAI221xp5_ASAP7_75t_R g1784 ( 
.A1(n_1764),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.C(n_310),
.Y(n_1784)
);

AOI221xp5_ASAP7_75t_L g1785 ( 
.A1(n_1763),
.A2(n_311),
.B1(n_313),
.B2(n_314),
.C(n_315),
.Y(n_1785)
);

OAI211xp5_ASAP7_75t_SL g1786 ( 
.A1(n_1760),
.A2(n_316),
.B(n_318),
.C(n_321),
.Y(n_1786)
);

A2O1A1Ixp33_ASAP7_75t_SL g1787 ( 
.A1(n_1771),
.A2(n_323),
.B(n_324),
.C(n_325),
.Y(n_1787)
);

XOR2xp5_ASAP7_75t_L g1788 ( 
.A(n_1769),
.B(n_326),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1770),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1770),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1769),
.B(n_328),
.Y(n_1791)
);

AOI21xp33_ASAP7_75t_SL g1792 ( 
.A1(n_1762),
.A2(n_329),
.B(n_330),
.Y(n_1792)
);

AOI321xp33_ASAP7_75t_L g1793 ( 
.A1(n_1782),
.A2(n_332),
.A3(n_334),
.B1(n_336),
.B2(n_337),
.C(n_338),
.Y(n_1793)
);

NOR4xp75_ASAP7_75t_L g1794 ( 
.A(n_1777),
.B(n_339),
.C(n_342),
.D(n_343),
.Y(n_1794)
);

HB1xp67_ASAP7_75t_L g1795 ( 
.A(n_1782),
.Y(n_1795)
);

AOI221xp5_ASAP7_75t_L g1796 ( 
.A1(n_1792),
.A2(n_347),
.B1(n_349),
.B2(n_351),
.C(n_352),
.Y(n_1796)
);

AOI222xp33_ASAP7_75t_L g1797 ( 
.A1(n_1779),
.A2(n_355),
.B1(n_356),
.B2(n_357),
.C1(n_358),
.C2(n_360),
.Y(n_1797)
);

OAI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1788),
.A2(n_361),
.B1(n_364),
.B2(n_365),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1773),
.B(n_366),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1791),
.B(n_367),
.Y(n_1800)
);

AOI32xp33_ASAP7_75t_L g1801 ( 
.A1(n_1775),
.A2(n_368),
.A3(n_369),
.B1(n_370),
.B2(n_371),
.Y(n_1801)
);

NOR3xp33_ASAP7_75t_L g1802 ( 
.A(n_1789),
.B(n_373),
.C(n_374),
.Y(n_1802)
);

AOI221xp5_ASAP7_75t_L g1803 ( 
.A1(n_1774),
.A2(n_1780),
.B1(n_1786),
.B2(n_1787),
.C(n_1781),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1795),
.B(n_1790),
.Y(n_1804)
);

OAI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1799),
.A2(n_1785),
.B1(n_1784),
.B2(n_1778),
.Y(n_1805)
);

INVx4_ASAP7_75t_L g1806 ( 
.A(n_1793),
.Y(n_1806)
);

NOR3xp33_ASAP7_75t_L g1807 ( 
.A(n_1800),
.B(n_1776),
.C(n_1783),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1794),
.Y(n_1808)
);

NOR2x1_ASAP7_75t_L g1809 ( 
.A(n_1798),
.B(n_376),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1803),
.A2(n_379),
.B1(n_380),
.B2(n_381),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1802),
.B(n_382),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1804),
.A2(n_1796),
.B(n_1801),
.Y(n_1812)
);

NAND5xp2_ASAP7_75t_L g1813 ( 
.A(n_1807),
.B(n_1797),
.C(n_384),
.D(n_386),
.E(n_387),
.Y(n_1813)
);

NOR3xp33_ASAP7_75t_L g1814 ( 
.A(n_1806),
.B(n_1808),
.C(n_1809),
.Y(n_1814)
);

NOR2x1p5_ASAP7_75t_L g1815 ( 
.A(n_1811),
.B(n_383),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1815),
.Y(n_1816)
);

NOR2x1_ASAP7_75t_L g1817 ( 
.A(n_1812),
.B(n_1805),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1816),
.Y(n_1818)
);

AOI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1817),
.A2(n_1814),
.B1(n_1810),
.B2(n_1813),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1819),
.Y(n_1820)
);

AO22x2_ASAP7_75t_L g1821 ( 
.A1(n_1818),
.A2(n_388),
.B1(n_390),
.B2(n_393),
.Y(n_1821)
);

AOI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1820),
.A2(n_394),
.B1(n_395),
.B2(n_396),
.Y(n_1822)
);

AOI221xp5_ASAP7_75t_L g1823 ( 
.A1(n_1821),
.A2(n_397),
.B1(n_398),
.B2(n_399),
.C(n_400),
.Y(n_1823)
);

AOI31xp33_ASAP7_75t_L g1824 ( 
.A1(n_1823),
.A2(n_401),
.A3(n_405),
.B(n_406),
.Y(n_1824)
);

AOI31xp33_ASAP7_75t_L g1825 ( 
.A1(n_1822),
.A2(n_407),
.A3(n_408),
.B(n_410),
.Y(n_1825)
);

OAI22xp5_ASAP7_75t_SL g1826 ( 
.A1(n_1824),
.A2(n_411),
.B1(n_413),
.B2(n_414),
.Y(n_1826)
);

AOI211xp5_ASAP7_75t_L g1827 ( 
.A1(n_1825),
.A2(n_419),
.B(n_420),
.C(n_421),
.Y(n_1827)
);

AOI221xp5_ASAP7_75t_L g1828 ( 
.A1(n_1826),
.A2(n_423),
.B1(n_424),
.B2(n_425),
.C(n_426),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1827),
.B(n_427),
.Y(n_1829)
);

OR2x6_ASAP7_75t_L g1830 ( 
.A(n_1826),
.B(n_428),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1826),
.B(n_429),
.Y(n_1831)
);

NAND3xp33_ASAP7_75t_L g1832 ( 
.A(n_1829),
.B(n_430),
.C(n_431),
.Y(n_1832)
);

AOI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1830),
.A2(n_434),
.B(n_435),
.Y(n_1833)
);

AOI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1831),
.A2(n_437),
.B1(n_438),
.B2(n_439),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1832),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1833),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1834),
.Y(n_1837)
);

OR2x6_ASAP7_75t_L g1838 ( 
.A(n_1836),
.B(n_1828),
.Y(n_1838)
);

O2A1O1Ixp5_ASAP7_75t_L g1839 ( 
.A1(n_1838),
.A2(n_1835),
.B(n_1837),
.C(n_444),
.Y(n_1839)
);

AOI211xp5_ASAP7_75t_L g1840 ( 
.A1(n_1839),
.A2(n_440),
.B(n_442),
.C(n_445),
.Y(n_1840)
);


endmodule