module fake_jpeg_8898_n_301 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_245;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

HB1xp67_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_41),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_30),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NAND2xp33_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_8),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_31),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_49),
.Y(n_68)
);

CKINVDCx12_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_48),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_27),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_20),
.C(n_34),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_20),
.C(n_34),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_31),
.B1(n_23),
.B2(n_34),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_59),
.B1(n_22),
.B2(n_33),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_55),
.A2(n_26),
.B(n_22),
.C(n_25),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_63),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_31),
.B1(n_23),
.B2(n_20),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_23),
.B1(n_20),
.B2(n_19),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_17),
.B1(n_26),
.B2(n_25),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_32),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_22),
.C(n_15),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_40),
.B1(n_35),
.B2(n_37),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_71),
.A2(n_46),
.B1(n_47),
.B2(n_60),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_77),
.B1(n_84),
.B2(n_55),
.Y(n_96)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_44),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_82),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_47),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_13),
.B(n_16),
.Y(n_118)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_96),
.A2(n_82),
.B1(n_71),
.B2(n_81),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_53),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_84),
.B(n_72),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_101),
.A2(n_21),
.B1(n_43),
.B2(n_22),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_50),
.C(n_49),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_48),
.C(n_65),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_77),
.A2(n_61),
.B1(n_45),
.B2(n_37),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_103),
.A2(n_104),
.B1(n_107),
.B2(n_116),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_86),
.A2(n_61),
.B1(n_45),
.B2(n_43),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_93),
.A2(n_43),
.B1(n_29),
.B2(n_28),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_78),
.A2(n_33),
.B(n_22),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_109),
.B(n_33),
.C(n_73),
.Y(n_138)
);

AND2x4_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_33),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_83),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_68),
.A2(n_43),
.B1(n_29),
.B2(n_28),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_117),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_118),
.B(n_120),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_70),
.B(n_65),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_89),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_140),
.Y(n_152)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_124),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_95),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_131),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_69),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_128),
.B(n_134),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_137),
.C(n_146),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_130),
.B(n_103),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_121),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_71),
.B1(n_81),
.B2(n_92),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_133),
.A2(n_136),
.B1(n_144),
.B2(n_145),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_114),
.B(n_71),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_105),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_135),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_85),
.B1(n_87),
.B2(n_73),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_138),
.A2(n_141),
.B(n_101),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_139),
.A2(n_97),
.B1(n_106),
.B2(n_110),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_29),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_109),
.A2(n_21),
.B1(n_24),
.B2(n_33),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_107),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_112),
.A2(n_29),
.B1(n_28),
.B2(n_21),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_109),
.A2(n_28),
.B1(n_24),
.B2(n_65),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_109),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_57),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_120),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_108),
.A2(n_57),
.B1(n_24),
.B2(n_8),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_149),
.A2(n_138),
.B1(n_141),
.B2(n_129),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_98),
.B(n_117),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_150),
.A2(n_159),
.B(n_171),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_135),
.Y(n_153)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_154),
.A2(n_166),
.B1(n_14),
.B2(n_13),
.Y(n_189)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_169),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_105),
.Y(n_163)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_143),
.A2(n_125),
.B1(n_133),
.B2(n_147),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_164),
.A2(n_176),
.B1(n_125),
.B2(n_144),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_98),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_139),
.C(n_57),
.Y(n_185)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_173),
.Y(n_190)
);

AO21x1_ASAP7_75t_L g171 ( 
.A1(n_134),
.A2(n_116),
.B(n_57),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_172),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_131),
.B(n_100),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_123),
.B(n_106),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_177),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_122),
.B(n_100),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_0),
.B(n_1),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_178),
.A2(n_142),
.B(n_149),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_181),
.A2(n_205),
.B1(n_153),
.B2(n_168),
.Y(n_207)
);

A2O1A1O1Ixp25_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_137),
.B(n_147),
.C(n_132),
.D(n_145),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_177),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_183),
.A2(n_186),
.B(n_10),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_195),
.C(n_200),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_154),
.A2(n_111),
.B(n_1),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_167),
.B(n_14),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_187),
.B(n_178),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_189),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_0),
.C(n_1),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_175),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_175),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_166),
.A2(n_162),
.B1(n_179),
.B2(n_164),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_152),
.B(n_2),
.Y(n_199)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_199),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_2),
.C(n_3),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_152),
.B(n_3),
.C(n_4),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_170),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_209),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_207),
.A2(n_210),
.B1(n_197),
.B2(n_196),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_201),
.A2(n_173),
.B(n_156),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_208),
.A2(n_227),
.B(n_205),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_193),
.A2(n_158),
.B1(n_171),
.B2(n_156),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_188),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_213),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_169),
.Y(n_212)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_192),
.B(n_163),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_161),
.Y(n_214)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_161),
.Y(n_215)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_183),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_199),
.B(n_155),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_220),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_182),
.Y(n_235)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_224),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_155),
.Y(n_222)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

A2O1A1Ixp33_ASAP7_75t_SL g223 ( 
.A1(n_186),
.A2(n_171),
.B(n_165),
.C(n_160),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_223),
.A2(n_193),
.B(n_201),
.Y(n_233)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_185),
.C(n_187),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_244),
.C(n_225),
.Y(n_255)
);

OAI21x1_ASAP7_75t_SL g250 ( 
.A1(n_233),
.A2(n_236),
.B(n_245),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_235),
.B(n_239),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_180),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_238),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_200),
.Y(n_238)
);

XNOR2x1_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_189),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_209),
.A2(n_194),
.B(n_180),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_240),
.A2(n_224),
.B1(n_215),
.B2(n_214),
.Y(n_252)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_243),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_195),
.C(n_184),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_226),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_259),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_219),
.B1(n_194),
.B2(n_181),
.Y(n_251)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_251),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_252),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_228),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_231),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_239),
.A2(n_207),
.B1(n_223),
.B2(n_227),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_254),
.B(n_257),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_244),
.C(n_229),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_234),
.A2(n_223),
.B1(n_219),
.B2(n_228),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_246),
.A2(n_223),
.B1(n_165),
.B2(n_203),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_233),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_236),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_240),
.A2(n_216),
.B1(n_160),
.B2(n_10),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_261),
.A2(n_243),
.B(n_236),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_262),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_265),
.C(n_270),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_230),
.C(n_238),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_250),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_269),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_249),
.C(n_258),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_247),
.C(n_241),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_254),
.B(n_257),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_256),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_260),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_275),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_266),
.A2(n_272),
.B1(n_264),
.B2(n_268),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_280),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_251),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_278),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_265),
.B(n_263),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_256),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_9),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_L g286 ( 
.A1(n_279),
.A2(n_273),
.A3(n_270),
.B1(n_259),
.B2(n_9),
.C1(n_10),
.C2(n_12),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_286),
.B(n_287),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_SL g289 ( 
.A1(n_274),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_289),
.A2(n_5),
.B(n_6),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_283),
.A2(n_12),
.B1(n_9),
.B2(n_7),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_281),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_291),
.B(n_292),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_284),
.B(n_282),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_293),
.A2(n_295),
.B(n_288),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_285),
.A2(n_282),
.B(n_280),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_296),
.B(n_294),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_R g299 ( 
.A(n_298),
.B(n_297),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_289),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_289),
.Y(n_301)
);


endmodule