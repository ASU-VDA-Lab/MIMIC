module fake_jpeg_9761_n_170 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_170);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_38),
.Y(n_40)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

AOI21xp33_ASAP7_75t_L g41 ( 
.A1(n_29),
.A2(n_25),
.B(n_28),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_38),
.B(n_26),
.C(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_30),
.B(n_16),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_17),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_31),
.A2(n_24),
.B1(n_19),
.B2(n_28),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_53),
.B1(n_22),
.B2(n_15),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_14),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_37),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_14),
.Y(n_50)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_0),
.B(n_1),
.Y(n_71)
);

NOR2x1_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_24),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_29),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_31),
.A2(n_19),
.B1(n_22),
.B2(n_27),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_55),
.B(n_56),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_57),
.B(n_60),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_44),
.Y(n_84)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_65),
.Y(n_76)
);

XOR2x1_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_68),
.Y(n_74)
);

OR2x6_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_26),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_54),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_15),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_51),
.B(n_36),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_42),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_49),
.Y(n_70)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_72),
.B(n_84),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_61),
.B(n_58),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_78),
.A2(n_59),
.B1(n_68),
.B2(n_56),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_89),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_44),
.B1(n_38),
.B2(n_33),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_86),
.B1(n_49),
.B2(n_39),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

NOR3xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_87),
.C(n_32),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_57),
.A2(n_33),
.B1(n_51),
.B2(n_48),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_54),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

NOR2x1_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_56),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_92),
.B(n_98),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_55),
.Y(n_94)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_79),
.B(n_78),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_59),
.Y(n_97)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_102),
.Y(n_120)
);

A2O1A1O1Ixp25_ASAP7_75t_L g100 ( 
.A1(n_74),
.A2(n_32),
.B(n_34),
.C(n_35),
.D(n_39),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_96),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_104),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_34),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_34),
.Y(n_105)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_106),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_81),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_113),
.C(n_114),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_75),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_79),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_116),
.B(n_117),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_78),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_85),
.C(n_72),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_95),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_99),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_78),
.B(n_87),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_127),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_100),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_132),
.C(n_133),
.Y(n_144)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_91),
.Y(n_126)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_93),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_128),
.B(n_131),
.Y(n_141)
);

OAI32xp33_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_106),
.A3(n_78),
.B1(n_101),
.B2(n_77),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_77),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_114),
.B(n_8),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_134),
.B(n_12),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_125),
.A2(n_112),
.B(n_111),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_136),
.A2(n_143),
.B(n_11),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_138),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_115),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_118),
.B1(n_117),
.B2(n_42),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_140),
.A2(n_141),
.B1(n_135),
.B2(n_136),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_130),
.B(n_7),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_129),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_146),
.C(n_35),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_130),
.C(n_129),
.Y(n_146)
);

OA21x2_ASAP7_75t_SL g147 ( 
.A1(n_139),
.A2(n_8),
.B(n_11),
.Y(n_147)
);

OAI31xp33_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_149),
.A3(n_2),
.B(n_3),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

FAx1_ASAP7_75t_SL g149 ( 
.A(n_140),
.B(n_35),
.CI(n_2),
.CON(n_149),
.SN(n_149)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_151),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_1),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_155),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_148),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

OAI221xp5_ASAP7_75t_L g160 ( 
.A1(n_157),
.A2(n_149),
.B1(n_3),
.B2(n_152),
.C(n_145),
.Y(n_160)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_146),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_161),
.B(n_163),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_158),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_162),
.B(n_155),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_159),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_168),
.Y(n_169)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_166),
.Y(n_170)
);


endmodule