module real_jpeg_25902_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_347, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_347;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g70 ( 
.A(n_0),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_1),
.A2(n_86),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_1),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_1),
.A2(n_68),
.B1(n_69),
.B2(n_97),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_97),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_97),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_37),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_2),
.A2(n_37),
.B1(n_68),
.B2(n_69),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_2),
.A2(n_37),
.B1(n_96),
.B2(n_299),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_3),
.A2(n_89),
.B(n_91),
.Y(n_88)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_3),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_3),
.B(n_81),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g169 ( 
.A1(n_3),
.A2(n_35),
.B1(n_36),
.B2(n_93),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_3),
.B(n_30),
.C(n_31),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_3),
.B(n_71),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_3),
.A2(n_45),
.B1(n_190),
.B2(n_197),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_6),
.A2(n_68),
.B1(n_69),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_6),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_6),
.A2(n_35),
.B1(n_36),
.B2(n_75),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_75),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_6),
.A2(n_75),
.B1(n_89),
.B2(n_235),
.Y(n_234)
);

INVx8_ASAP7_75t_SL g84 ( 
.A(n_7),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_8),
.A2(n_68),
.B1(n_69),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_8),
.A2(n_73),
.B1(n_96),
.B2(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_73),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_73),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_51),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_9),
.A2(n_51),
.B1(n_68),
.B2(n_69),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_9),
.A2(n_51),
.B1(n_89),
.B2(n_235),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_43),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_10),
.A2(n_43),
.B1(n_68),
.B2(n_69),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_10),
.A2(n_43),
.B1(n_86),
.B2(n_96),
.Y(n_285)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_12),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_12),
.A2(n_60),
.B1(n_68),
.B2(n_69),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_60),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_12),
.A2(n_60),
.B1(n_86),
.B2(n_96),
.Y(n_260)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_13),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_15),
.Y(n_191)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_340),
.C(n_344),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_338),
.B(n_343),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_328),
.B(n_337),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_293),
.A3(n_323),
.B1(n_326),
.B2(n_327),
.C(n_347),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_269),
.B(n_292),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_245),
.B(n_268),
.Y(n_21)
);

O2A1O1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_133),
.B(n_218),
.C(n_244),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_118),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_24),
.B(n_118),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_100),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_56),
.B1(n_98),
.B2(n_99),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_26),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_26),
.B(n_99),
.C(n_100),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_44),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_27),
.B(n_44),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_34),
.B(n_38),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_28),
.B(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_28),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_28),
.B(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_28),
.B(n_93),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_28),
.A2(n_162),
.B(n_310),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_29),
.B(n_203),
.Y(n_202)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_34),
.Y(n_227)
);

AO22x1_ASAP7_75t_L g71 ( 
.A1(n_35),
.A2(n_36),
.B1(n_66),
.B2(n_67),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_35),
.B(n_66),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

OAI32xp33_ASAP7_75t_L g140 ( 
.A1(n_36),
.A2(n_67),
.A3(n_69),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_36),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_38),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_41),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_59),
.B(n_61),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_39),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_39),
.A2(n_150),
.B(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_39),
.A2(n_149),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_39),
.A2(n_148),
.B1(n_149),
.B2(n_170),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_39),
.A2(n_149),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_39),
.A2(n_61),
.B(n_228),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_39),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_49),
.B(n_52),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_45),
.A2(n_52),
.B(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_45),
.A2(n_180),
.B(n_181),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_45),
.A2(n_187),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_45),
.A2(n_144),
.B(n_198),
.Y(n_253)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_46),
.A2(n_47),
.B1(n_50),
.B2(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_46),
.B(n_53),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_46),
.A2(n_186),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_48),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g182 ( 
.A(n_55),
.Y(n_182)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_62),
.C(n_77),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_57),
.A2(n_58),
.B1(n_62),
.B2(n_121),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_59),
.Y(n_162)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_72),
.B1(n_74),
.B2(n_76),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_63),
.A2(n_74),
.B(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_63),
.A2(n_72),
.B1(n_76),
.B2(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_63),
.A2(n_238),
.B(n_239),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_63),
.A2(n_76),
.B1(n_263),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_64),
.A2(n_71),
.B1(n_132),
.B2(n_141),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_64),
.B(n_240),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_64),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_64),
.A2(n_71),
.B(n_110),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_71),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_69),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_68),
.A2(n_83),
.B(n_92),
.C(n_113),
.Y(n_112)
);

HAxp5_ASAP7_75t_SL g141 ( 
.A(n_68),
.B(n_93),
.CON(n_141),
.SN(n_141)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

NAND3xp33_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_82),
.C(n_106),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_71),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_71),
.B(n_240),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_76),
.A2(n_263),
.B(n_264),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_77),
.B(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_80),
.B1(n_88),
.B2(n_94),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_79),
.A2(n_81),
.B1(n_95),
.B2(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_79),
.A2(n_81),
.B1(n_104),
.B2(n_234),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_79),
.A2(n_234),
.B(n_259),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_79),
.A2(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_79),
.B(n_301),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_79),
.A2(n_81),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_79),
.A2(n_284),
.B(n_317),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_79),
.A2(n_81),
.B(n_283),
.Y(n_344)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_85),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_80),
.B(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_80),
.B(n_285),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_80),
.A2(n_298),
.B(n_300),
.Y(n_297)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_L g85 ( 
.A1(n_82),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_89),
.Y(n_235)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_90),
.B(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_93),
.B(n_198),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVx8_ASAP7_75t_L g299 ( 
.A(n_96),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_111),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_107),
.B2(n_108),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_103),
.B(n_107),
.C(n_111),
.Y(n_242)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_109),
.B(n_264),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_110),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_114),
.B1(n_115),
.B2(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_126),
.B(n_127),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.C(n_124),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_119),
.B(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_122),
.B(n_124),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.C(n_130),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_128),
.B1(n_129),
.B2(n_155),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_125),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_127),
.B(n_181),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_213),
.B(n_217),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_164),
.B(n_212),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_151),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_138),
.B(n_151),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_146),
.C(n_147),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_139),
.B(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_143),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_146),
.B(n_147),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_156),
.B2(n_157),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_152),
.B(n_159),
.C(n_163),
.Y(n_214)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_163),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_158),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_161),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_207),
.B(n_211),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_183),
.B(n_206),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_173),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_167),
.B(n_173),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_171),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_179),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_178),
.C(n_179),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_177),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

AOI21xp33_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_193),
.B(n_205),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_192),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_192),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_200),
.B(n_204),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_195),
.B(n_196),
.Y(n_204)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_208),
.B(n_209),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_214),
.B(n_215),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_220),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_242),
.B2(n_243),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_230),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_230),
.C(n_243),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_229),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_229),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_226),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_241),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_236),
.B2(n_237),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_233),
.B(n_236),
.C(n_241),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_239),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_242),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_246),
.B(n_247),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_267),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_254),
.B1(n_265),
.B2(n_266),
.Y(n_248)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_266),
.C(n_267),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_251),
.B(n_252),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_252),
.A2(n_253),
.B1(n_282),
.B2(n_286),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_252),
.A2(n_286),
.B(n_287),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_254),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_258),
.C(n_261),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_261),
.B2(n_262),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_259),
.Y(n_341)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_260),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_270),
.B(n_271),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_290),
.B2(n_291),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_280),
.B1(n_288),
.B2(n_289),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_274),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_274),
.B(n_289),
.C(n_291),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_277),
.B(n_279),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_277),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_278),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_295),
.C(n_311),
.Y(n_294)
);

FAx1_ASAP7_75t_L g325 ( 
.A(n_279),
.B(n_295),
.CI(n_311),
.CON(n_325),
.SN(n_325)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_280),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_287),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_282),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_290),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_312),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_294),
.B(n_312),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_302),
.B2(n_303),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_296),
.A2(n_297),
.B1(n_314),
.B2(n_321),
.Y(n_313)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_305),
.C(n_308),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_297),
.B(n_321),
.C(n_322),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_298),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_300),
.B(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_308),
.B2(n_309),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_308),
.A2(n_309),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_309),
.B(n_315),
.C(n_319),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_322),
.Y(n_312)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_314),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_318),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_324),
.B(n_325),
.Y(n_326)
);

BUFx24_ASAP7_75t_SL g345 ( 
.A(n_325),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_330),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_336),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_332),
.A2(n_333),
.B1(n_334),
.B2(n_335),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_332),
.B(n_335),
.C(n_336),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_333),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_335),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_342),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_340),
.B(n_342),
.Y(n_343)
);


endmodule