module real_jpeg_32728_n_10 (n_8, n_0, n_93, n_95, n_2, n_91, n_9, n_92, n_97, n_6, n_7, n_3, n_99, n_5, n_4, n_98, n_94, n_1, n_96, n_10);

input n_8;
input n_0;
input n_93;
input n_95;
input n_2;
input n_91;
input n_9;
input n_92;
input n_97;
input n_6;
input n_7;
input n_3;
input n_99;
input n_5;
input n_4;
input n_98;
input n_94;
input n_1;
input n_96;

output n_10;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_89;
wire n_16;

AOI221xp5_ASAP7_75t_L g49 ( 
.A1(n_0),
.A2(n_9),
.B1(n_50),
.B2(n_56),
.C(n_57),
.Y(n_49)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g11 ( 
.A1(n_1),
.A2(n_12),
.B1(n_13),
.B2(n_19),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_2),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_2),
.B(n_83),
.Y(n_87)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_4),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_5),
.B(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_6),
.B(n_33),
.Y(n_81)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_7),
.B(n_23),
.Y(n_89)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_9),
.B(n_50),
.C(n_56),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_20),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

NOR2x1_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_15),
.Y(n_13)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_29),
.B(n_88),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_28),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_82),
.B(n_87),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_40),
.B(n_80),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_39),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_96),
.Y(n_56)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_71),
.C(n_72),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_61),
.B(n_70),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_49),
.B1(n_59),
.B2(n_60),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_69),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_69),
.Y(n_70)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2x1_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_91),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_92),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_93),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_94),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_95),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_97),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_98),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_99),
.Y(n_84)
);


endmodule