module fake_jpeg_14173_n_590 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_590);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_590;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_16),
.B(n_17),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_15),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx6f_ASAP7_75t_SL g59 ( 
.A(n_1),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_8),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_62),
.B(n_83),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_18),
.B(n_29),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_63),
.B(n_71),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_64),
.Y(n_166)
);

INVx11_ASAP7_75t_SL g65 ( 
.A(n_34),
.Y(n_65)
);

INVx5_ASAP7_75t_SL g195 ( 
.A(n_65),
.Y(n_195)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_7),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_67),
.B(n_72),
.Y(n_159)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_20),
.B(n_10),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_24),
.B(n_10),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_73),
.B(n_74),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_34),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_75),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_76),
.Y(n_153)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_77),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_78),
.Y(n_161)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_79),
.Y(n_182)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_80),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_81),
.Y(n_179)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_82),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_24),
.B(n_10),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_84),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_86),
.Y(n_146)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_34),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_90),
.B(n_96),
.Y(n_168)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_26),
.B(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_98),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_34),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_94),
.B(n_97),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_26),
.B(n_6),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_95),
.B(n_114),
.Y(n_183)
);

INVx4_ASAP7_75t_SL g96 ( 
.A(n_34),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_43),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_27),
.B(n_58),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_99),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_101),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_50),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_102),
.B(n_106),
.Y(n_160)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_22),
.Y(n_103)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_103),
.Y(n_184)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_25),
.Y(n_104)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_22),
.Y(n_105)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_105),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_29),
.B(n_6),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_25),
.Y(n_107)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_21),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_21),
.Y(n_109)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_109),
.Y(n_170)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_21),
.Y(n_110)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_110),
.Y(n_187)
);

BUFx12_ASAP7_75t_L g111 ( 
.A(n_21),
.Y(n_111)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_27),
.B(n_17),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_13),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_32),
.B(n_6),
.Y(n_114)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_22),
.Y(n_115)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_21),
.Y(n_117)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_117),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_57),
.B(n_4),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_118),
.B(n_0),
.Y(n_171)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_30),
.Y(n_120)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_120),
.Y(n_181)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_46),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_121),
.B(n_123),
.Y(n_174)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_122),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_46),
.B(n_4),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_23),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_124),
.B(n_44),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_63),
.A2(n_23),
.B1(n_30),
.B2(n_53),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_125),
.A2(n_131),
.B1(n_172),
.B2(n_173),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_75),
.A2(n_57),
.B1(n_107),
.B2(n_23),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_128),
.A2(n_176),
.B(n_193),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_71),
.A2(n_37),
.B1(n_32),
.B2(n_41),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_70),
.A2(n_57),
.B1(n_35),
.B2(n_40),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_141),
.A2(n_158),
.B1(n_191),
.B2(n_108),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_142),
.B(n_150),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_118),
.B(n_37),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_145),
.B(n_147),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_117),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_123),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_61),
.A2(n_40),
.B1(n_35),
.B2(n_39),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g169 ( 
.A(n_68),
.B(n_33),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_169),
.B(n_171),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_85),
.A2(n_49),
.B1(n_41),
.B2(n_42),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_92),
.A2(n_49),
.B1(n_42),
.B2(n_53),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_75),
.A2(n_30),
.B1(n_53),
.B2(n_44),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_73),
.B(n_56),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_178),
.B(n_199),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_110),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_82),
.A2(n_56),
.B1(n_54),
.B2(n_51),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_186),
.A2(n_201),
.B1(n_204),
.B2(n_2),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_90),
.B(n_44),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_188),
.B(n_112),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_107),
.B(n_54),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_189),
.B(n_192),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_78),
.A2(n_51),
.B1(n_48),
.B2(n_44),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_88),
.B(n_48),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_66),
.A2(n_44),
.B1(n_33),
.B2(n_11),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_104),
.A2(n_33),
.B1(n_4),
.B2(n_3),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_196),
.A2(n_116),
.B1(n_99),
.B2(n_86),
.Y(n_225)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_89),
.Y(n_198)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_81),
.A2(n_33),
.B1(n_4),
.B2(n_3),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_91),
.Y(n_202)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_202),
.Y(n_247)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_119),
.Y(n_203)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_203),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_122),
.A2(n_33),
.B1(n_11),
.B2(n_14),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_205),
.A2(n_208),
.B1(n_266),
.B2(n_267),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_0),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_206),
.B(n_217),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_141),
.A2(n_101),
.B1(n_105),
.B2(n_120),
.Y(n_208)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_152),
.Y(n_210)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_210),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_211),
.B(n_222),
.Y(n_291)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_139),
.Y(n_212)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_212),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_149),
.B(n_109),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_213),
.B(n_216),
.Y(n_282)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_139),
.Y(n_214)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_214),
.Y(n_298)
);

BUFx12f_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_215),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_168),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_127),
.B(n_0),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_169),
.B(n_87),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_218),
.B(n_270),
.C(n_190),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_84),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_219),
.B(n_220),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_77),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_221),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_138),
.B(n_115),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_159),
.B(n_103),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_224),
.B(n_241),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_225),
.A2(n_258),
.B1(n_153),
.B2(n_166),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_134),
.B(n_0),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_227),
.B(n_246),
.Y(n_308)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_228),
.Y(n_323)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_229),
.Y(n_278)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_155),
.Y(n_230)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_230),
.Y(n_277)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_184),
.Y(n_231)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_231),
.Y(n_301)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_140),
.Y(n_232)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_232),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_168),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_233),
.B(n_248),
.Y(n_280)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_133),
.Y(n_234)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_234),
.Y(n_285)
);

AND2x4_ASAP7_75t_L g236 ( 
.A(n_144),
.B(n_96),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_236),
.B(n_237),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_188),
.Y(n_237)
);

INVx11_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_238),
.Y(n_281)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_156),
.Y(n_239)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_239),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_160),
.B(n_100),
.Y(n_241)
);

OA22x2_ASAP7_75t_L g242 ( 
.A1(n_191),
.A2(n_79),
.B1(n_65),
.B2(n_111),
.Y(n_242)
);

OAI32xp33_ASAP7_75t_L g296 ( 
.A1(n_242),
.A2(n_146),
.A3(n_148),
.B1(n_161),
.B2(n_179),
.Y(n_296)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_164),
.Y(n_243)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_243),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_157),
.B(n_15),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_244),
.B(n_269),
.Y(n_326)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_164),
.Y(n_245)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_245),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_175),
.B(n_1),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_163),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_151),
.B(n_2),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_249),
.B(n_257),
.Y(n_317)
);

INVx13_ASAP7_75t_L g250 ( 
.A(n_199),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_250),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_153),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_251),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_194),
.Y(n_252)
);

INVx8_ASAP7_75t_L g295 ( 
.A(n_252),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_133),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_255),
.Y(n_283)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_181),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_254),
.B(n_256),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_158),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_177),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_136),
.B(n_2),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_165),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_259),
.B(n_260),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_197),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_126),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_261),
.Y(n_288)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_167),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_264),
.Y(n_300)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_170),
.Y(n_264)
);

NOR2x1_ASAP7_75t_L g307 ( 
.A(n_265),
.B(n_148),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_L g266 ( 
.A1(n_176),
.A2(n_111),
.B1(n_64),
.B2(n_76),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_193),
.A2(n_2),
.B1(n_14),
.B2(n_15),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_187),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_268),
.B(n_271),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_143),
.B(n_14),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_162),
.B(n_154),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_137),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_128),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_272),
.B(n_273),
.Y(n_315)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_186),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_274),
.B(n_236),
.Y(n_319)
);

AO22x1_ASAP7_75t_L g276 ( 
.A1(n_185),
.A2(n_154),
.B1(n_146),
.B2(n_196),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_276),
.A2(n_275),
.B(n_265),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_205),
.A2(n_208),
.B1(n_237),
.B2(n_233),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_279),
.A2(n_290),
.B1(n_305),
.B2(n_311),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_284),
.B(n_286),
.Y(n_337)
);

OAI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_240),
.A2(n_185),
.B1(n_190),
.B2(n_130),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_287),
.A2(n_309),
.B1(n_327),
.B2(n_221),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_258),
.A2(n_129),
.B1(n_132),
.B2(n_179),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_296),
.A2(n_316),
.B1(n_318),
.B2(n_321),
.Y(n_345)
);

FAx1_ASAP7_75t_SL g299 ( 
.A(n_217),
.B(n_130),
.CI(n_166),
.CON(n_299),
.SN(n_299)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_299),
.B(n_284),
.Y(n_369)
);

AOI32xp33_ASAP7_75t_L g302 ( 
.A1(n_207),
.A2(n_177),
.A3(n_200),
.B1(n_137),
.B2(n_129),
.Y(n_302)
);

A2O1A1O1Ixp25_ASAP7_75t_L g343 ( 
.A1(n_302),
.A2(n_238),
.B(n_250),
.C(n_234),
.D(n_251),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_218),
.A2(n_132),
.B1(n_161),
.B2(n_135),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_307),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_240),
.A2(n_135),
.B1(n_182),
.B2(n_275),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_207),
.A2(n_182),
.B1(n_267),
.B2(n_266),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_207),
.B(n_226),
.C(n_265),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_313),
.B(n_236),
.C(n_210),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_314),
.B(n_333),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_242),
.A2(n_270),
.B1(n_239),
.B2(n_263),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_242),
.A2(n_270),
.B1(n_261),
.B2(n_276),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_319),
.B(n_289),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_242),
.A2(n_261),
.B1(n_276),
.B2(n_247),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_227),
.B(n_246),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_324),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_257),
.B(n_249),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_235),
.A2(n_223),
.B1(n_206),
.B2(n_271),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_236),
.A2(n_232),
.B1(n_254),
.B2(n_209),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_335),
.B(n_347),
.C(n_349),
.Y(n_380)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_328),
.Y(n_338)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_338),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_339),
.Y(n_392)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_328),
.Y(n_340)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_340),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_291),
.B(n_215),
.Y(n_341)
);

INVxp33_ASAP7_75t_L g397 ( 
.A(n_341),
.Y(n_397)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_277),
.Y(n_342)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_342),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_343),
.A2(n_331),
.B(n_310),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_315),
.A2(n_289),
.B(n_319),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_344),
.A2(n_310),
.B(n_332),
.Y(n_388)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_277),
.Y(n_346)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_346),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_313),
.B(n_230),
.C(n_262),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_294),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_348),
.B(n_354),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_317),
.B(n_324),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_309),
.A2(n_245),
.B1(n_243),
.B2(n_231),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_350),
.A2(n_353),
.B1(n_288),
.B2(n_283),
.Y(n_384)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_312),
.Y(n_351)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_351),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_304),
.A2(n_228),
.B1(n_253),
.B2(n_256),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_280),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_312),
.Y(n_355)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_355),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_291),
.B(n_215),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_356),
.B(n_358),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_325),
.A2(n_252),
.B1(n_214),
.B2(n_212),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_357),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_325),
.B(n_229),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_303),
.Y(n_359)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_359),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_317),
.B(n_322),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_360),
.B(n_361),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_308),
.B(n_306),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_315),
.A2(n_314),
.B(n_289),
.Y(n_362)
);

AOI21xp33_ASAP7_75t_L g389 ( 
.A1(n_362),
.A2(n_364),
.B(n_369),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_327),
.B(n_326),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_363),
.B(n_366),
.Y(n_401)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_303),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_365),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_326),
.B(n_292),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_308),
.B(n_306),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_368),
.B(n_371),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_303),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_372),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_299),
.B(n_305),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_320),
.Y(n_372)
);

AO22x1_ASAP7_75t_SL g373 ( 
.A1(n_304),
.A2(n_296),
.B1(n_302),
.B2(n_311),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_373),
.B(n_374),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_282),
.B(n_307),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_300),
.Y(n_376)
);

CKINVDCx14_ASAP7_75t_R g407 ( 
.A(n_376),
.Y(n_407)
);

INVx5_ASAP7_75t_L g377 ( 
.A(n_285),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_377),
.B(n_378),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_333),
.B(n_288),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_349),
.B(n_299),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_381),
.B(n_360),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_384),
.A2(n_410),
.B1(n_370),
.B2(n_359),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_347),
.B(n_301),
.C(n_330),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_387),
.B(n_400),
.C(n_403),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_388),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_356),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_390),
.B(n_402),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_391),
.B(n_339),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_352),
.A2(n_285),
.B1(n_330),
.B2(n_332),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_394),
.A2(n_405),
.B1(n_408),
.B2(n_350),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_335),
.B(n_301),
.C(n_329),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_378),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_336),
.B(n_281),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_352),
.A2(n_293),
.B1(n_298),
.B2(n_323),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_337),
.A2(n_293),
.B1(n_298),
.B2(n_323),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_371),
.A2(n_297),
.B1(n_281),
.B2(n_278),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_362),
.A2(n_331),
.B(n_334),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_411),
.A2(n_414),
.B(n_367),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_375),
.A2(n_334),
.B(n_295),
.Y(n_414)
);

CKINVDCx14_ASAP7_75t_R g415 ( 
.A(n_375),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_415),
.B(n_375),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_417),
.Y(n_452)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_379),
.Y(n_418)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_418),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_396),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_419),
.B(n_421),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_420),
.B(n_399),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_396),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_381),
.B(n_336),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_422),
.B(n_447),
.Y(n_456)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_379),
.Y(n_423)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_423),
.Y(n_455)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_382),
.Y(n_424)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_424),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_401),
.B(n_366),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_425),
.B(n_428),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_SL g459 ( 
.A(n_426),
.B(n_411),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_416),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_380),
.B(n_368),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_429),
.B(n_440),
.C(n_441),
.Y(n_464)
);

FAx1_ASAP7_75t_SL g430 ( 
.A(n_398),
.B(n_361),
.CI(n_369),
.CON(n_430),
.SN(n_430)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_430),
.A2(n_432),
.B1(n_434),
.B2(n_435),
.Y(n_460)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_382),
.Y(n_431)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_431),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_401),
.B(n_363),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_395),
.A2(n_337),
.B(n_345),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_433),
.A2(n_445),
.B(n_414),
.Y(n_473)
);

CKINVDCx14_ASAP7_75t_R g435 ( 
.A(n_385),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_406),
.B(n_348),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_436),
.A2(n_438),
.B1(n_446),
.B2(n_390),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_392),
.A2(n_337),
.B1(n_373),
.B2(n_343),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_393),
.Y(n_439)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_439),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_380),
.B(n_344),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_400),
.B(n_387),
.C(n_403),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_393),
.Y(n_442)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_442),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_386),
.B(n_372),
.Y(n_443)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_443),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_403),
.B(n_364),
.C(n_374),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_444),
.B(n_383),
.C(n_388),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_406),
.B(n_354),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_386),
.B(n_358),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_449),
.A2(n_410),
.B1(n_384),
.B2(n_402),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_440),
.B(n_398),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_457),
.B(n_462),
.C(n_465),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_458),
.B(n_470),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_459),
.A2(n_473),
.B(n_415),
.Y(n_493)
);

CKINVDCx14_ASAP7_75t_R g500 ( 
.A(n_461),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_429),
.B(n_399),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_463),
.A2(n_434),
.B1(n_421),
.B2(n_437),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_427),
.B(n_389),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_438),
.A2(n_416),
.B1(n_391),
.B2(n_373),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_467),
.A2(n_478),
.B1(n_445),
.B2(n_448),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_445),
.A2(n_448),
.B1(n_449),
.B2(n_419),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_469),
.A2(n_417),
.B1(n_426),
.B2(n_385),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_427),
.B(n_389),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_472),
.B(n_476),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_432),
.A2(n_407),
.B1(n_394),
.B2(n_405),
.Y(n_474)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_474),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_441),
.B(n_383),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_444),
.B(n_420),
.C(n_422),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_477),
.B(n_365),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_433),
.A2(n_373),
.B1(n_353),
.B2(n_408),
.Y(n_478)
);

NAND3xp33_ASAP7_75t_L g479 ( 
.A(n_451),
.B(n_407),
.C(n_443),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_479),
.B(n_455),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_480),
.A2(n_494),
.B1(n_495),
.B2(n_502),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_468),
.B(n_409),
.Y(n_481)
);

NAND3xp33_ASAP7_75t_SL g516 ( 
.A(n_481),
.B(n_486),
.C(n_454),
.Y(n_516)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_466),
.Y(n_482)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_482),
.Y(n_519)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_450),
.Y(n_483)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_483),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_469),
.B(n_383),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_484),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_485),
.A2(n_462),
.B1(n_458),
.B2(n_456),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_409),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_487),
.A2(n_477),
.B1(n_475),
.B2(n_471),
.Y(n_512)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_466),
.Y(n_490)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_490),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_460),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_491),
.B(n_492),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_450),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_493),
.B(n_503),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_463),
.A2(n_430),
.B1(n_447),
.B2(n_439),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_473),
.A2(n_430),
.B1(n_442),
.B2(n_431),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_453),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_496),
.B(n_498),
.Y(n_508)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_453),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_452),
.A2(n_397),
.B(n_423),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_499),
.A2(n_404),
.B(n_340),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_478),
.A2(n_424),
.B1(n_418),
.B2(n_413),
.Y(n_501)
);

INVxp33_ASAP7_75t_L g521 ( 
.A(n_501),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_452),
.A2(n_413),
.B1(n_412),
.B2(n_404),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_500),
.A2(n_467),
.B1(n_470),
.B2(n_457),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_507),
.B(n_510),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_488),
.B(n_464),
.C(n_476),
.Y(n_510)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_511),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_SL g542 ( 
.A1(n_512),
.A2(n_526),
.B(n_513),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_497),
.A2(n_482),
.B1(n_490),
.B2(n_487),
.Y(n_513)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_513),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_495),
.B(n_494),
.Y(n_515)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_515),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_516),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_481),
.B(n_412),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_517),
.B(n_523),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_518),
.A2(n_498),
.B(n_496),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_488),
.B(n_464),
.Y(n_523)
);

CKINVDCx14_ASAP7_75t_R g524 ( 
.A(n_486),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_524),
.B(n_484),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_525),
.A2(n_456),
.B1(n_472),
.B2(n_465),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_502),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_528),
.B(n_529),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_510),
.B(n_504),
.C(n_489),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_514),
.B(n_499),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_532),
.B(n_538),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_515),
.A2(n_493),
.B(n_484),
.Y(n_534)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_534),
.Y(n_548)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_537),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_523),
.B(n_504),
.C(n_489),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_509),
.B(n_485),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_539),
.B(n_542),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_505),
.B(n_377),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_540),
.B(n_512),
.Y(n_556)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_541),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_506),
.B(n_483),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_543),
.B(n_506),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_543),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_545),
.B(n_550),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_535),
.A2(n_536),
.B1(n_533),
.B2(n_522),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_547),
.A2(n_553),
.B1(n_541),
.B2(n_519),
.Y(n_561)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_549),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_530),
.B(n_505),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_530),
.B(n_521),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_552),
.B(n_556),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_543),
.A2(n_525),
.B1(n_519),
.B2(n_522),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_531),
.B(n_509),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_SL g563 ( 
.A(n_557),
.B(n_527),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_551),
.B(n_539),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_558),
.B(n_559),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_544),
.B(n_542),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_561),
.A2(n_562),
.B1(n_563),
.B2(n_549),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_548),
.A2(n_526),
.B1(n_507),
.B2(n_534),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_548),
.B(n_555),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_564),
.B(n_554),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_556),
.A2(n_529),
.B(n_538),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_565),
.B(n_549),
.C(n_520),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_546),
.B(n_528),
.C(n_520),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_568),
.B(n_553),
.C(n_554),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_569),
.B(n_570),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_560),
.B(n_547),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_571),
.B(n_572),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_574),
.B(n_355),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_567),
.B(n_508),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_SL g581 ( 
.A(n_575),
.B(n_338),
.Y(n_581)
);

AO21x1_ASAP7_75t_L g576 ( 
.A1(n_566),
.A2(n_517),
.B(n_508),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_576),
.A2(n_561),
.B1(n_568),
.B2(n_562),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_L g584 ( 
.A1(n_577),
.A2(n_580),
.B(n_582),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_SL g580 ( 
.A1(n_573),
.A2(n_558),
.B(n_518),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_SL g583 ( 
.A(n_581),
.B(n_346),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_583),
.A2(n_585),
.B1(n_342),
.B2(n_351),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_L g585 ( 
.A1(n_578),
.A2(n_570),
.B(n_576),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_584),
.B(n_579),
.C(n_582),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_586),
.B(n_587),
.C(n_297),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_588),
.B(n_295),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_589),
.B(n_278),
.Y(n_590)
);


endmodule