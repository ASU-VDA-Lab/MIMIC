module real_jpeg_28416_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_0),
.B(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_0),
.B(n_28),
.Y(n_27)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_0),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_0),
.A2(n_21),
.B(n_78),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_0),
.B(n_210),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_1),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_1),
.A2(n_26),
.B1(n_33),
.B2(n_35),
.Y(n_86)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_4),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_4),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_4),
.A2(n_33),
.B1(n_35),
.B2(n_51),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_4),
.A2(n_22),
.B1(n_23),
.B2(n_51),
.Y(n_210)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_6),
.A2(n_22),
.B1(n_23),
.B2(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_6),
.A2(n_29),
.B1(n_33),
.B2(n_35),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_6),
.A2(n_29),
.B1(n_49),
.B2(n_50),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_6),
.A2(n_29),
.B1(n_54),
.B2(n_55),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_7),
.A2(n_33),
.B1(n_35),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_7),
.A2(n_41),
.B1(n_54),
.B2(n_55),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_7),
.A2(n_22),
.B1(n_23),
.B2(n_41),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_7),
.B(n_49),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_7),
.A2(n_49),
.B(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_7),
.B(n_93),
.Y(n_165)
);

AOI21xp33_ASAP7_75t_SL g175 ( 
.A1(n_7),
.A2(n_10),
.B(n_33),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g201 ( 
.A1(n_7),
.A2(n_23),
.B(n_38),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_7),
.B(n_71),
.Y(n_205)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_10),
.Y(n_66)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_10),
.A2(n_33),
.B1(n_35),
.B2(n_70),
.Y(n_71)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_11),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_138),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_137),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_111),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_16),
.B(n_111),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_75),
.C(n_88),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_17),
.B(n_75),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_44),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_18),
.B(n_46),
.C(n_62),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_30),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_19),
.B(n_30),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_25),
.B(n_27),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_20),
.B(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_21),
.B(n_78),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_21),
.B(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_22),
.A2(n_23),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_22),
.B(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_25),
.A2(n_81),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_27),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_27),
.B(n_209),
.Y(n_221)
);

INVxp33_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_39),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_31),
.A2(n_86),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_31),
.B(n_192),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_36),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_32),
.B(n_42),
.Y(n_87)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_33),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_33),
.A2(n_37),
.B(n_41),
.C(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_36),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_36),
.B(n_40),
.Y(n_191)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_39),
.B(n_181),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_42),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_40),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_41),
.A2(n_55),
.B(n_66),
.C(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_41),
.B(n_85),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_41),
.B(n_110),
.Y(n_225)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_42),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_42),
.B(n_182),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_62),
.B2(n_63),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_58),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_47),
.B(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_48),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_52),
.B(n_53),
.C(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_53),
.Y(n_61)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_52)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_54),
.B(n_57),
.Y(n_105)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_66),
.B(n_67),
.C(n_71),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_55),
.A2(n_105),
.B1(n_106),
.B2(n_108),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_59),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_60),
.B(n_121),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_72),
.B(n_73),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_65),
.B(n_74),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_65),
.B(n_126),
.Y(n_152)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_71),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_71),
.B(n_102),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_73),
.Y(n_99)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_84),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_84),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_77),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

INVx5_ASAP7_75t_SL g110 ( 
.A(n_79),
.Y(n_110)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_82),
.B(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B(n_87),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_85),
.A2(n_133),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_87),
.B(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_88),
.A2(n_89),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_98),
.C(n_103),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_90),
.A2(n_91),
.B1(n_98),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_93),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_98),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_101),
.B(n_125),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_103),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_109),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_104),
.B(n_109),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_136),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_129),
.B2(n_130),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_122),
.B2(n_123),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_128),
.B(n_151),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_134),
.B2(n_135),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_131),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_131),
.A2(n_134),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_131),
.B(n_174),
.Y(n_193)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

O2A1O1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_168),
.B(n_243),
.C(n_248),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_156),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_140),
.B(n_156),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_153),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_142),
.B(n_143),
.C(n_153),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.C(n_149),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_146),
.A2(n_147),
.B1(n_149),
.B2(n_150),
.Y(n_159)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.C(n_162),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_157),
.A2(n_158),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_162),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.C(n_166),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_166),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_167),
.B(n_215),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_242),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_235),
.B(n_241),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_194),
.B(n_234),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_183),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_172),
.B(n_183),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.C(n_179),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_173),
.B(n_232),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_174),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_232)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_188),
.B2(n_189),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_184),
.B(n_190),
.C(n_193),
.Y(n_236)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_229),
.B(n_233),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_211),
.B(n_228),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_202),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_197),
.B(n_202),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_200),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_208),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_207),
.C(n_208),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_218),
.B(n_227),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_216),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_213),
.B(n_216),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_222),
.B(n_226),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_220),
.B(n_221),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_230),
.B(n_231),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_236),
.B(n_237),
.Y(n_241)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_244),
.B(n_245),
.Y(n_248)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);


endmodule