module fake_ariane_485_n_779 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_14, n_88, n_141, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_779);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_779;

wire n_295;
wire n_556;
wire n_356;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_423;
wire n_347;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_756;
wire n_466;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_143;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_331;
wire n_320;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_206;
wire n_538;
wire n_352;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_543;
wire n_362;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_444;
wire n_355;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_769;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_147;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_580;
wire n_358;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_92),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_7),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

BUFx10_ASAP7_75t_L g145 ( 
.A(n_56),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_42),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_33),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_140),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_139),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_23),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_66),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_62),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_19),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_50),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_127),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_48),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_116),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_124),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_136),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_138),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_65),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_36),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_64),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_70),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_12),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_133),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_101),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_38),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_45),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_6),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_34),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_93),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_73),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_15),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_120),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_16),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_37),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_35),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_128),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_17),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_117),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_63),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_105),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_95),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_4),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_2),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_11),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_80),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_129),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_49),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_54),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_132),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_85),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_134),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_171),
.Y(n_197)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_150),
.B(n_0),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_168),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_142),
.Y(n_207)
);

AND2x4_ASAP7_75t_L g208 ( 
.A(n_165),
.B(n_0),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_1),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

AND2x4_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_1),
.Y(n_211)
);

INVxp33_ASAP7_75t_SL g212 ( 
.A(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_144),
.B(n_2),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_145),
.B(n_3),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_3),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_172),
.B(n_4),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_143),
.Y(n_219)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_145),
.B(n_5),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_175),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_178),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_175),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_153),
.B(n_5),
.Y(n_226)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_192),
.Y(n_229)
);

AND2x4_ASAP7_75t_L g230 ( 
.A(n_146),
.B(n_6),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_193),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_179),
.B(n_7),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_193),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_177),
.Y(n_234)
);

BUFx8_ASAP7_75t_SL g235 ( 
.A(n_187),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_L g236 ( 
.A1(n_212),
.A2(n_187),
.B1(n_181),
.B2(n_149),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_225),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_L g239 ( 
.A1(n_209),
.A2(n_191),
.B1(n_183),
.B2(n_184),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_147),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_197),
.Y(n_242)
);

AND2x4_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_148),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_151),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_225),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_226),
.A2(n_190),
.B1(n_189),
.B2(n_182),
.Y(n_247)
);

AND2x2_ASAP7_75t_SL g248 ( 
.A(n_214),
.B(n_152),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_R g249 ( 
.A1(n_226),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_204),
.B(n_154),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_L g251 ( 
.A1(n_214),
.A2(n_180),
.B1(n_176),
.B2(n_173),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_221),
.A2(n_170),
.B1(n_169),
.B2(n_167),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_222),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_L g255 ( 
.A1(n_222),
.A2(n_166),
.B1(n_164),
.B2(n_163),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_155),
.Y(n_256)
);

AO22x2_ASAP7_75t_L g257 ( 
.A1(n_230),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_257)
);

INVx8_ASAP7_75t_L g258 ( 
.A(n_230),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_199),
.A2(n_161),
.B1(n_160),
.B2(n_159),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_230),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_219),
.B(n_156),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_225),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_230),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_208),
.A2(n_158),
.B1(n_157),
.B2(n_13),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_L g265 ( 
.A1(n_213),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_L g266 ( 
.A1(n_217),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_266)
);

AO22x2_ASAP7_75t_L g267 ( 
.A1(n_208),
.A2(n_14),
.B1(n_17),
.B2(n_18),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_224),
.B(n_18),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_208),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_232),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_208),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_234),
.B(n_27),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_223),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_211),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_274)
);

NAND2xp33_ASAP7_75t_SL g275 ( 
.A(n_211),
.B(n_31),
.Y(n_275)
);

OAI22xp33_ASAP7_75t_L g276 ( 
.A1(n_211),
.A2(n_32),
.B1(n_39),
.B2(n_40),
.Y(n_276)
);

AO22x2_ASAP7_75t_L g277 ( 
.A1(n_211),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_218),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_234),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_L g280 ( 
.A1(n_224),
.A2(n_46),
.B1(n_47),
.B2(n_51),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_216),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_234),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_238),
.Y(n_283)
);

XOR2x2_ASAP7_75t_L g284 ( 
.A(n_248),
.B(n_252),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_279),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_234),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_244),
.B(n_201),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_240),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_282),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_242),
.B(n_235),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_237),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_245),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_246),
.Y(n_294)
);

XNOR2x2_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_201),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_262),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_260),
.B(n_201),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_278),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_261),
.B(n_202),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_254),
.B(n_202),
.Y(n_300)
);

XNOR2x2_ASAP7_75t_L g301 ( 
.A(n_267),
.B(n_202),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_272),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_253),
.B(n_233),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_268),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_243),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_263),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_236),
.B(n_203),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_277),
.B(n_233),
.Y(n_308)
);

OR2x2_ASAP7_75t_SL g309 ( 
.A(n_249),
.B(n_203),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_241),
.B(n_203),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_250),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_251),
.B(n_243),
.Y(n_312)
);

AND2x4_ASAP7_75t_L g313 ( 
.A(n_252),
.B(n_206),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_259),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_259),
.B(n_206),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_264),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_264),
.Y(n_317)
);

NAND2xp33_ASAP7_75t_R g318 ( 
.A(n_277),
.B(n_206),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_258),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_258),
.B(n_231),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_257),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_257),
.B(n_231),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_258),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_275),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_269),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_239),
.B(n_231),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_247),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_269),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_255),
.B(n_233),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_271),
.B(n_218),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_271),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_L g332 ( 
.A(n_274),
.B(n_198),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_270),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g334 ( 
.A(n_265),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_274),
.B(n_196),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_276),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_266),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_281),
.B(n_233),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_281),
.B(n_233),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_280),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_279),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_238),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_274),
.B(n_198),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_237),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_244),
.B(n_196),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_243),
.B(n_198),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_299),
.B(n_200),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_325),
.B(n_200),
.Y(n_348)
);

AND2x4_ASAP7_75t_L g349 ( 
.A(n_313),
.B(n_57),
.Y(n_349)
);

AND2x6_ASAP7_75t_L g350 ( 
.A(n_331),
.B(n_200),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_310),
.B(n_200),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_285),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_286),
.B(n_200),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_289),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_338),
.A2(n_227),
.B(n_220),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_315),
.B(n_210),
.Y(n_356)
);

AND2x2_ASAP7_75t_SL g357 ( 
.A(n_338),
.B(n_210),
.Y(n_357)
);

AND2x4_ASAP7_75t_SL g358 ( 
.A(n_346),
.B(n_228),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_315),
.B(n_210),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_292),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_346),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_344),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_310),
.B(n_210),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_R g364 ( 
.A(n_288),
.B(n_314),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_341),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_293),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_313),
.B(n_210),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_300),
.B(n_215),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_322),
.B(n_215),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_294),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_296),
.Y(n_371)
);

INVxp33_ASAP7_75t_L g372 ( 
.A(n_307),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_341),
.B(n_215),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_298),
.Y(n_374)
);

NOR2xp67_ASAP7_75t_L g375 ( 
.A(n_319),
.B(n_198),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_290),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_320),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_311),
.B(n_215),
.Y(n_378)
);

INVx5_ASAP7_75t_L g379 ( 
.A(n_335),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_323),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_302),
.B(n_215),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_305),
.B(n_328),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_283),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_312),
.B(n_228),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_312),
.B(n_228),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_326),
.B(n_228),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_326),
.B(n_228),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_330),
.B(n_198),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_342),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_337),
.B(n_198),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_297),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_297),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g393 ( 
.A(n_324),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_321),
.B(n_58),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_334),
.B(n_205),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_287),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_287),
.B(n_205),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_306),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_304),
.Y(n_399)
);

NOR2xp67_ASAP7_75t_SL g400 ( 
.A(n_340),
.B(n_205),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_343),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_295),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_345),
.B(n_205),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_301),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_343),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_321),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_333),
.B(n_205),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_329),
.B(n_284),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_345),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_329),
.B(n_205),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_339),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_303),
.B(n_220),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_308),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_408),
.B(n_336),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_364),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_406),
.B(n_327),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_360),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_369),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_369),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_361),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_379),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_396),
.B(n_332),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_396),
.B(n_316),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g424 ( 
.A(n_408),
.B(n_309),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_361),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_406),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_361),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_379),
.Y(n_428)
);

AND2x6_ASAP7_75t_L g429 ( 
.A(n_349),
.B(n_318),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_382),
.B(n_317),
.Y(n_430)
);

BUFx8_ASAP7_75t_SL g431 ( 
.A(n_399),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_361),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_409),
.B(n_318),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_382),
.B(n_291),
.Y(n_434)
);

OR2x6_ASAP7_75t_L g435 ( 
.A(n_402),
.B(n_59),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_349),
.B(n_220),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_372),
.B(n_402),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_409),
.B(n_220),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_402),
.B(n_60),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_365),
.B(n_220),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_349),
.B(n_220),
.Y(n_441)
);

NAND2x1_ASAP7_75t_SL g442 ( 
.A(n_402),
.B(n_67),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_399),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_413),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_411),
.B(n_227),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_360),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_411),
.B(n_404),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_404),
.B(n_227),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_404),
.B(n_68),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_371),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_399),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_379),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_404),
.B(n_69),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_349),
.B(n_394),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_394),
.B(n_71),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_378),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_383),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_371),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_383),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_394),
.B(n_72),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_384),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_394),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_383),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_389),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_412),
.B(n_227),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_371),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_379),
.B(n_227),
.Y(n_467)
);

OR2x6_ASAP7_75t_L g468 ( 
.A(n_398),
.B(n_74),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_365),
.B(n_227),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_371),
.Y(n_470)
);

BUFx12f_ASAP7_75t_L g471 ( 
.A(n_444),
.Y(n_471)
);

INVx6_ASAP7_75t_L g472 ( 
.A(n_450),
.Y(n_472)
);

INVx3_ASAP7_75t_SL g473 ( 
.A(n_415),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_433),
.B(n_391),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_454),
.B(n_379),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_431),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_457),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_417),
.Y(n_478)
);

NAND2xp33_ASAP7_75t_L g479 ( 
.A(n_429),
.B(n_398),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_454),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_L g481 ( 
.A1(n_414),
.A2(n_413),
.B1(n_379),
.B2(n_405),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_423),
.Y(n_482)
);

BUFx8_ASAP7_75t_SL g483 ( 
.A(n_423),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_R g484 ( 
.A(n_436),
.B(n_398),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_450),
.Y(n_485)
);

BUFx2_ASAP7_75t_SL g486 ( 
.A(n_455),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_446),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_459),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_426),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_463),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_429),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_464),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_450),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_458),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_458),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_443),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_458),
.Y(n_497)
);

INVx3_ASAP7_75t_SL g498 ( 
.A(n_455),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_451),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_426),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_466),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_418),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_433),
.B(n_379),
.Y(n_503)
);

BUFx12f_ASAP7_75t_L g504 ( 
.A(n_416),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_416),
.B(n_389),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_466),
.Y(n_506)
);

NAND2x1p5_ASAP7_75t_L g507 ( 
.A(n_460),
.B(n_401),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_466),
.Y(n_508)
);

NAND2x1p5_ASAP7_75t_L g509 ( 
.A(n_460),
.B(n_401),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_420),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_430),
.Y(n_511)
);

INVx8_ASAP7_75t_L g512 ( 
.A(n_429),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_419),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_470),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_470),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_470),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_447),
.B(n_429),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_434),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_SL g519 ( 
.A1(n_486),
.A2(n_441),
.B1(n_436),
.B2(n_439),
.Y(n_519)
);

BUFx4f_ASAP7_75t_SL g520 ( 
.A(n_471),
.Y(n_520)
);

INVx6_ASAP7_75t_L g521 ( 
.A(n_471),
.Y(n_521)
);

INVx11_ASAP7_75t_L g522 ( 
.A(n_504),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_482),
.A2(n_441),
.B1(n_449),
.B2(n_439),
.Y(n_523)
);

INVx1_ASAP7_75t_SL g524 ( 
.A(n_489),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_490),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_502),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_473),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_SL g528 ( 
.A1(n_486),
.A2(n_449),
.B1(n_453),
.B2(n_413),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_502),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_513),
.Y(n_530)
);

CKINVDCx11_ASAP7_75t_R g531 ( 
.A(n_473),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_490),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_504),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_513),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_473),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_511),
.A2(n_437),
.B1(n_453),
.B2(n_435),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_476),
.Y(n_537)
);

INVx6_ASAP7_75t_L g538 ( 
.A(n_472),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_474),
.B(n_461),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_496),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_477),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_477),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_498),
.A2(n_462),
.B1(n_468),
.B2(n_391),
.Y(n_543)
);

INVx6_ASAP7_75t_L g544 ( 
.A(n_472),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_476),
.Y(n_545)
);

CKINVDCx11_ASAP7_75t_R g546 ( 
.A(n_518),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_488),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_503),
.B(n_461),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_488),
.Y(n_549)
);

BUFx8_ASAP7_75t_L g550 ( 
.A(n_489),
.Y(n_550)
);

BUFx12f_ASAP7_75t_L g551 ( 
.A(n_500),
.Y(n_551)
);

NAND2x1p5_ASAP7_75t_L g552 ( 
.A(n_491),
.B(n_421),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_505),
.A2(n_435),
.B1(n_424),
.B2(n_456),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_500),
.B(n_505),
.Y(n_554)
);

INVx5_ASAP7_75t_L g555 ( 
.A(n_512),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_503),
.A2(n_422),
.B(n_438),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_496),
.Y(n_557)
);

BUFx4f_ASAP7_75t_SL g558 ( 
.A(n_505),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_498),
.A2(n_468),
.B1(n_392),
.B2(n_435),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_492),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_492),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_481),
.A2(n_445),
.B1(n_483),
.B2(n_517),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_523),
.A2(n_498),
.B1(n_468),
.B2(n_509),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_519),
.A2(n_507),
.B1(n_509),
.B2(n_380),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_554),
.B(n_378),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_555),
.B(n_493),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_SL g567 ( 
.A1(n_559),
.A2(n_484),
.B1(n_509),
.B2(n_507),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_524),
.B(n_480),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_528),
.A2(n_422),
.B1(n_512),
.B2(n_491),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_551),
.B(n_480),
.Y(n_570)
);

BUFx4f_ASAP7_75t_SL g571 ( 
.A(n_537),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_536),
.A2(n_512),
.B1(n_491),
.B2(n_465),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_524),
.B(n_475),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_SL g574 ( 
.A(n_520),
.B(n_512),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_559),
.A2(n_553),
.B1(n_546),
.B2(n_562),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_538),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_539),
.A2(n_357),
.B1(n_352),
.B2(n_354),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_531),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_543),
.A2(n_405),
.B1(n_401),
.B2(n_556),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_541),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_SL g581 ( 
.A1(n_543),
.A2(n_507),
.B(n_385),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_539),
.A2(n_380),
.B1(n_392),
.B2(n_389),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_525),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_532),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_SL g585 ( 
.A1(n_558),
.A2(n_479),
.B1(n_357),
.B2(n_401),
.Y(n_585)
);

INVx5_ASAP7_75t_L g586 ( 
.A(n_555),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_526),
.Y(n_587)
);

OAI21xp33_ASAP7_75t_L g588 ( 
.A1(n_556),
.A2(n_381),
.B(n_380),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_529),
.B(n_530),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_540),
.Y(n_590)
);

OAI22xp33_ASAP7_75t_L g591 ( 
.A1(n_548),
.A2(n_393),
.B1(n_352),
.B2(n_354),
.Y(n_591)
);

OAI21xp5_ASAP7_75t_SL g592 ( 
.A1(n_533),
.A2(n_548),
.B(n_385),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_545),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_557),
.A2(n_401),
.B1(n_405),
.B2(n_428),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_521),
.Y(n_595)
);

AOI21xp33_ASAP7_75t_L g596 ( 
.A1(n_534),
.A2(n_348),
.B(n_384),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_SL g597 ( 
.A1(n_550),
.A2(n_479),
.B1(n_357),
.B2(n_405),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_555),
.B(n_527),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_535),
.A2(n_393),
.B1(n_432),
.B2(n_420),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_SL g600 ( 
.A1(n_552),
.A2(n_475),
.B(n_412),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_535),
.B(n_367),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_538),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_542),
.B(n_499),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_547),
.B(n_499),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_552),
.A2(n_355),
.B(n_351),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_SL g606 ( 
.A1(n_550),
.A2(n_405),
.B1(n_401),
.B2(n_350),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_L g607 ( 
.A1(n_521),
.A2(n_393),
.B1(n_432),
.B2(n_425),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_549),
.B(n_560),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_561),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_538),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_544),
.B(n_510),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_568),
.B(n_544),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_573),
.B(n_544),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_581),
.A2(n_522),
.B1(n_452),
.B2(n_421),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_565),
.B(n_493),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_592),
.A2(n_452),
.B1(n_428),
.B2(n_352),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_572),
.A2(n_405),
.B1(n_374),
.B2(n_376),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_575),
.A2(n_354),
.B1(n_510),
.B2(n_472),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_597),
.A2(n_374),
.B1(n_376),
.B2(n_478),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_597),
.A2(n_374),
.B1(n_376),
.B2(n_478),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_585),
.A2(n_487),
.B1(n_370),
.B2(n_366),
.Y(n_621)
);

AOI221xp5_ASAP7_75t_SL g622 ( 
.A1(n_601),
.A2(n_381),
.B1(n_353),
.B2(n_366),
.C(n_370),
.Y(n_622)
);

OAI221xp5_ASAP7_75t_L g623 ( 
.A1(n_600),
.A2(n_442),
.B1(n_370),
.B2(n_366),
.C(n_348),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_585),
.A2(n_487),
.B1(n_371),
.B2(n_400),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_579),
.A2(n_569),
.B1(n_563),
.B2(n_567),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_SL g626 ( 
.A1(n_564),
.A2(n_350),
.B1(n_555),
.B2(n_356),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_569),
.A2(n_472),
.B1(n_425),
.B2(n_427),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_574),
.A2(n_400),
.B1(n_395),
.B2(n_350),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_577),
.A2(n_350),
.B1(n_356),
.B2(n_359),
.Y(n_629)
);

NAND3xp33_ASAP7_75t_L g630 ( 
.A(n_580),
.B(n_347),
.C(n_353),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_598),
.B(n_485),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_580),
.B(n_589),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_567),
.A2(n_427),
.B1(n_494),
.B2(n_501),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_602),
.B(n_514),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_577),
.A2(n_501),
.B1(n_494),
.B2(n_506),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_607),
.A2(n_501),
.B1(n_494),
.B2(n_506),
.Y(n_636)
);

OAI22xp33_ASAP7_75t_L g637 ( 
.A1(n_571),
.A2(n_516),
.B1(n_515),
.B2(n_514),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_591),
.A2(n_350),
.B1(n_359),
.B2(n_371),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_SL g639 ( 
.A1(n_582),
.A2(n_350),
.B1(n_448),
.B2(n_355),
.Y(n_639)
);

NOR3xp33_ASAP7_75t_L g640 ( 
.A(n_599),
.B(n_497),
.C(n_351),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_591),
.A2(n_350),
.B1(n_367),
.B2(n_360),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_SL g642 ( 
.A1(n_586),
.A2(n_350),
.B1(n_388),
.B2(n_387),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_598),
.B(n_485),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_596),
.A2(n_362),
.B1(n_387),
.B2(n_386),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_583),
.A2(n_362),
.B1(n_377),
.B2(n_388),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_SL g646 ( 
.A1(n_586),
.A2(n_386),
.B1(n_515),
.B2(n_516),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_606),
.A2(n_497),
.B1(n_508),
.B2(n_495),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_SL g648 ( 
.A1(n_586),
.A2(n_390),
.B1(n_410),
.B2(n_485),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_608),
.B(n_485),
.Y(n_649)
);

OAI221xp5_ASAP7_75t_SL g650 ( 
.A1(n_588),
.A2(n_347),
.B1(n_363),
.B2(n_368),
.C(n_373),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_632),
.B(n_587),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_649),
.B(n_609),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_613),
.B(n_604),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_612),
.Y(n_654)
);

OAI221xp5_ASAP7_75t_SL g655 ( 
.A1(n_623),
.A2(n_603),
.B1(n_606),
.B2(n_611),
.C(n_595),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_615),
.B(n_610),
.Y(n_656)
);

NAND3xp33_ASAP7_75t_SL g657 ( 
.A(n_614),
.B(n_593),
.C(n_578),
.Y(n_657)
);

OAI21xp5_ASAP7_75t_SL g658 ( 
.A1(n_616),
.A2(n_570),
.B(n_576),
.Y(n_658)
);

NAND4xp25_ASAP7_75t_L g659 ( 
.A(n_622),
.B(n_576),
.C(n_605),
.D(n_438),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_634),
.B(n_566),
.Y(n_660)
);

NAND3xp33_ASAP7_75t_L g661 ( 
.A(n_650),
.B(n_594),
.C(n_363),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_SL g662 ( 
.A1(n_625),
.A2(n_566),
.B(n_571),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_SL g663 ( 
.A1(n_626),
.A2(n_508),
.B(n_495),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_639),
.B(n_584),
.Y(n_664)
);

OAI221xp5_ASAP7_75t_L g665 ( 
.A1(n_630),
.A2(n_373),
.B1(n_368),
.B2(n_590),
.C(n_362),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_631),
.B(n_586),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_643),
.B(n_485),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_SL g668 ( 
.A1(n_647),
.A2(n_508),
.B(n_495),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_637),
.B(n_495),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_633),
.B(n_495),
.Y(n_670)
);

NAND3xp33_ASAP7_75t_L g671 ( 
.A(n_640),
.B(n_508),
.C(n_390),
.Y(n_671)
);

NAND2xp33_ASAP7_75t_L g672 ( 
.A(n_638),
.B(n_508),
.Y(n_672)
);

NAND3xp33_ASAP7_75t_L g673 ( 
.A(n_648),
.B(n_377),
.C(n_407),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_638),
.B(n_358),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_636),
.B(n_377),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_629),
.A2(n_407),
.B1(n_410),
.B2(n_358),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_641),
.B(n_358),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_SL g678 ( 
.A1(n_628),
.A2(n_467),
.B(n_469),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_635),
.B(n_469),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_654),
.B(n_624),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_656),
.B(n_641),
.Y(n_681)
);

NOR3xp33_ASAP7_75t_L g682 ( 
.A(n_671),
.B(n_627),
.C(n_618),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_656),
.B(n_619),
.Y(n_683)
);

OAI31xp33_ASAP7_75t_L g684 ( 
.A1(n_655),
.A2(n_629),
.A3(n_620),
.B(n_621),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_669),
.B(n_666),
.Y(n_685)
);

NAND4xp75_ASAP7_75t_L g686 ( 
.A(n_664),
.B(n_375),
.C(n_646),
.D(n_440),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_651),
.B(n_642),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_653),
.B(n_644),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_652),
.B(n_644),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_664),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_672),
.A2(n_617),
.B1(n_645),
.B2(n_375),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_660),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_670),
.B(n_75),
.Y(n_693)
);

NAND3xp33_ASAP7_75t_L g694 ( 
.A(n_662),
.B(n_440),
.C(n_397),
.Y(n_694)
);

NAND3xp33_ASAP7_75t_L g695 ( 
.A(n_659),
.B(n_397),
.C(n_403),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_672),
.A2(n_403),
.B1(n_77),
.B2(n_78),
.Y(n_696)
);

OAI211xp5_ASAP7_75t_SL g697 ( 
.A1(n_658),
.A2(n_76),
.B(n_79),
.C(n_81),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_690),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_692),
.B(n_668),
.Y(n_699)
);

XOR2x2_ASAP7_75t_L g700 ( 
.A(n_686),
.B(n_687),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_685),
.B(n_667),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_685),
.B(n_674),
.Y(n_702)
);

NAND4xp75_ASAP7_75t_L g703 ( 
.A(n_687),
.B(n_674),
.C(n_677),
.D(n_675),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_690),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_681),
.B(n_663),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_680),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_693),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_697),
.B(n_657),
.Y(n_708)
);

XNOR2x1_ASAP7_75t_L g709 ( 
.A(n_700),
.B(n_688),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_705),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_707),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_701),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_701),
.Y(n_713)
);

AOI22x1_ASAP7_75t_L g714 ( 
.A1(n_710),
.A2(n_699),
.B1(n_707),
.B2(n_702),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_710),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_712),
.B(n_705),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_713),
.B(n_702),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_711),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_709),
.A2(n_703),
.B1(n_708),
.B2(n_699),
.Y(n_719)
);

XNOR2x1_ASAP7_75t_L g720 ( 
.A(n_719),
.B(n_700),
.Y(n_720)
);

NOR2x1_ASAP7_75t_SL g721 ( 
.A(n_715),
.B(n_706),
.Y(n_721)
);

OAI322xp33_ASAP7_75t_L g722 ( 
.A1(n_716),
.A2(n_689),
.A3(n_706),
.B1(n_695),
.B2(n_661),
.C1(n_665),
.C2(n_673),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_714),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_723),
.A2(n_717),
.B1(n_718),
.B2(n_682),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_722),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_722),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_726),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_725),
.A2(n_720),
.B1(n_718),
.B2(n_721),
.Y(n_728)
);

OAI22x1_ASAP7_75t_L g729 ( 
.A1(n_724),
.A2(n_693),
.B1(n_704),
.B2(n_698),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_726),
.Y(n_730)
);

OA22x2_ASAP7_75t_L g731 ( 
.A1(n_730),
.A2(n_680),
.B1(n_681),
.B2(n_683),
.Y(n_731)
);

NOR4xp25_ASAP7_75t_L g732 ( 
.A(n_727),
.B(n_696),
.C(n_694),
.D(n_678),
.Y(n_732)
);

AOI221xp5_ASAP7_75t_L g733 ( 
.A1(n_728),
.A2(n_684),
.B1(n_683),
.B2(n_679),
.C(n_691),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_729),
.A2(n_677),
.B1(n_676),
.B2(n_84),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_730),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_728),
.A2(n_676),
.B1(n_83),
.B2(n_86),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_730),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_735),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_737),
.Y(n_739)
);

NOR2x1_ASAP7_75t_L g740 ( 
.A(n_732),
.B(n_82),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_734),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_731),
.Y(n_742)
);

INVxp67_ASAP7_75t_SL g743 ( 
.A(n_736),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_733),
.B(n_90),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_735),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_742),
.Y(n_746)
);

NOR2xp67_ASAP7_75t_L g747 ( 
.A(n_738),
.B(n_91),
.Y(n_747)
);

NAND4xp25_ASAP7_75t_L g748 ( 
.A(n_740),
.B(n_94),
.C(n_96),
.D(n_97),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_739),
.Y(n_749)
);

NOR3xp33_ASAP7_75t_SL g750 ( 
.A(n_745),
.B(n_98),
.C(n_99),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_744),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_743),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_741),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_742),
.Y(n_754)
);

AO22x2_ASAP7_75t_L g755 ( 
.A1(n_754),
.A2(n_100),
.B1(n_102),
.B2(n_103),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_752),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_749),
.B(n_752),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_747),
.B(n_104),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_746),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_751),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_753),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_748),
.A2(n_750),
.B1(n_107),
.B2(n_108),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_756),
.Y(n_763)
);

INVxp67_ASAP7_75t_L g764 ( 
.A(n_757),
.Y(n_764)
);

AO22x2_ASAP7_75t_L g765 ( 
.A1(n_759),
.A2(n_106),
.B1(n_109),
.B2(n_110),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_L g766 ( 
.A1(n_760),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_762),
.A2(n_761),
.B1(n_758),
.B2(n_755),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_755),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_768),
.Y(n_769)
);

INVxp67_ASAP7_75t_SL g770 ( 
.A(n_764),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_763),
.Y(n_771)
);

AO22x1_ASAP7_75t_L g772 ( 
.A1(n_770),
.A2(n_767),
.B1(n_766),
.B2(n_765),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_769),
.A2(n_141),
.B1(n_115),
.B2(n_118),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_771),
.A2(n_114),
.B1(n_119),
.B2(n_121),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_772),
.Y(n_775)
);

OAI22xp33_ASAP7_75t_L g776 ( 
.A1(n_775),
.A2(n_773),
.B1(n_774),
.B2(n_126),
.Y(n_776)
);

INVxp67_ASAP7_75t_SL g777 ( 
.A(n_776),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_777),
.A2(n_122),
.B1(n_125),
.B2(n_130),
.Y(n_778)
);

AOI211xp5_ASAP7_75t_L g779 ( 
.A1(n_778),
.A2(n_131),
.B(n_135),
.C(n_137),
.Y(n_779)
);


endmodule