module real_jpeg_7904_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_213;
wire n_179;
wire n_167;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_0),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_0),
.A2(n_39),
.B1(n_57),
.B2(n_58),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_0),
.A2(n_26),
.B1(n_29),
.B2(n_39),
.Y(n_157)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_2),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_L g155 ( 
.A1(n_2),
.A2(n_54),
.B(n_58),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_2),
.A2(n_52),
.B1(n_61),
.B2(n_154),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_2),
.B(n_65),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_2),
.A2(n_37),
.B(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_2),
.B(n_37),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_2),
.A2(n_81),
.B1(n_82),
.B2(n_230),
.Y(n_232)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_SL g70 ( 
.A(n_7),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_8),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_8),
.A2(n_28),
.B1(n_57),
.B2(n_58),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_8),
.A2(n_28),
.B1(n_37),
.B2(n_40),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_8),
.A2(n_28),
.B1(n_52),
.B2(n_61),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_10),
.A2(n_52),
.B1(n_61),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_10),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_10),
.A2(n_57),
.B1(n_58),
.B2(n_101),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_10),
.A2(n_26),
.B1(n_29),
.B2(n_101),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_10),
.A2(n_37),
.B1(n_40),
.B2(n_101),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_11),
.A2(n_52),
.B1(n_61),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_11),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_11),
.A2(n_57),
.B1(n_58),
.B2(n_150),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_11),
.A2(n_37),
.B1(n_40),
.B2(n_150),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_11),
.A2(n_26),
.B1(n_29),
.B2(n_150),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_12),
.A2(n_37),
.B1(n_40),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_12),
.A2(n_26),
.B1(n_29),
.B2(n_47),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_12),
.A2(n_47),
.B1(n_57),
.B2(n_58),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_13),
.A2(n_52),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_13),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_13),
.A2(n_57),
.B1(n_58),
.B2(n_62),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_13),
.A2(n_26),
.B1(n_29),
.B2(n_62),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_13),
.A2(n_37),
.B1(n_40),
.B2(n_62),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_15),
.A2(n_26),
.B1(n_29),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_15),
.A2(n_34),
.B1(n_52),
.B2(n_61),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_15),
.A2(n_34),
.B1(n_57),
.B2(n_58),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_15),
.A2(n_34),
.B1(n_37),
.B2(n_40),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_133),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_131),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_105),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_19),
.B(n_105),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_78),
.C(n_89),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_20),
.A2(n_21),
.B1(n_78),
.B2(n_160),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_48),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_22),
.B(n_49),
.C(n_77),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_35),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_23),
.B(n_35),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_32),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_24),
.A2(n_82),
.B(n_157),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_25),
.B(n_31),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_26),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_26),
.A2(n_29),
.B1(n_42),
.B2(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_26),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_221)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_29),
.B(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_29),
.B(n_45),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_29),
.B(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_30),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_30),
.A2(n_31),
.B1(n_211),
.B2(n_213),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_33),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_31),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_32),
.A2(n_81),
.B(n_214),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_33),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_41),
.B1(n_44),
.B2(n_46),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_36),
.A2(n_44),
.B(n_95),
.Y(n_94)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_42),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_37),
.A2(n_40),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_37),
.B(n_69),
.Y(n_258)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_40),
.A2(n_74),
.B1(n_253),
.B2(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_41),
.A2(n_46),
.B(n_85),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_41),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_41),
.A2(n_44),
.B1(n_218),
.B2(n_220),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_41),
.A2(n_44),
.B1(n_220),
.B2(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_41),
.A2(n_44),
.B1(n_243),
.B2(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_41),
.A2(n_124),
.B(n_251),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_42),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_43),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_44),
.B(n_87),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_44),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_44),
.B(n_154),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_66),
.B2(n_77),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_60),
.B(n_63),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_51),
.A2(n_56),
.B1(n_60),
.B2(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_51),
.A2(n_113),
.B(n_114),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_51),
.A2(n_56),
.B1(n_100),
.B2(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_51),
.Y(n_177)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B(n_55),
.C(n_56),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_53),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_52),
.A2(n_53),
.B(n_154),
.C(n_155),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_68),
.B(n_69),
.C(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_69),
.Y(n_74)
);

HAxp5_ASAP7_75t_SL g253 ( 
.A(n_58),
.B(n_154),
.CON(n_253),
.SN(n_253)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_64),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_65),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_66),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_71),
.B(n_72),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_76),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_67),
.A2(n_144),
.B1(n_145),
.B2(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_67),
.A2(n_144),
.B1(n_175),
.B2(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_67),
.B(n_154),
.Y(n_241)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_68),
.A2(n_73),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_68),
.B(n_103),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_68),
.A2(n_73),
.B1(n_198),
.B2(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_71),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_73),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_78),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_88),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_80),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_84),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B(n_83),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_81),
.A2(n_92),
.B(n_93),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_81),
.A2(n_82),
.B1(n_92),
.B2(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_81),
.A2(n_82),
.B1(n_212),
.B2(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_81),
.A2(n_83),
.B(n_93),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_82),
.B(n_154),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_84),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_86),
.A2(n_97),
.B(n_126),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_89),
.B(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_98),
.C(n_102),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_91),
.B(n_94),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_98),
.A2(n_99),
.B1(n_102),
.B2(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_102),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_129),
.B2(n_130),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_118),
.B1(n_119),
.B2(n_128),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_116),
.B2(n_117),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_116),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_123),
.B(n_127),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_123),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_129),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_161),
.B(n_284),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_158),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_135),
.B(n_158),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.C(n_140),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_136),
.B(n_139),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_140),
.A2(n_141),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_147),
.C(n_151),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_143),
.B1(n_147),
.B2(n_148),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_145),
.B(n_146),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_156),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_152),
.A2(n_153),
.B1(n_156),
.B2(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_156),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_203),
.Y(n_161)
);

INVxp33_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_184),
.B(n_202),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NOR3xp33_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_204),
.C(n_283),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_181),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_181),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.C(n_171),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.C(n_180),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_174),
.B1(n_180),
.B2(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_180),
.Y(n_190)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_182),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_185),
.B(n_187),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.C(n_193),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_188),
.B(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_191),
.A2(n_193),
.B1(n_194),
.B2(n_281),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_191),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_199),
.C(n_200),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_195),
.A2(n_196),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_269),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_199),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_277),
.B(n_282),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_262),
.B(n_276),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_246),
.B(n_261),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_237),
.B(n_245),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_226),
.B(n_236),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_215),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_210),
.B(n_215),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_221),
.B2(n_225),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_216),
.B(n_225),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_219),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_221),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_231),
.B(n_235),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_228),
.B(n_229),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_238),
.B(n_239),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_247),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_240),
.B(n_247),
.Y(n_261)
);

FAx1_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_242),
.CI(n_244),
.CON(n_240),
.SN(n_240)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_256),
.B2(n_260),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_250),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_252),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_255),
.C(n_260),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_256),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_259),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_259),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_263),
.B(n_264),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_270),
.B2(n_271),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_273),
.C(n_274),
.Y(n_278)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_272),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_273),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_278),
.B(n_279),
.Y(n_282)
);


endmodule