module fake_netlist_6_2798_n_1852 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1852);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1852;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1832;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_50),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_95),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_32),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_31),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_84),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_81),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_74),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_106),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_150),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_16),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_64),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_2),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_23),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_124),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_51),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_143),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_156),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_21),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_12),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_65),
.Y(n_196)
);

BUFx2_ASAP7_75t_SL g197 ( 
.A(n_3),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_166),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_137),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_3),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_175),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_113),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_72),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_104),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_133),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_35),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_169),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_9),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_33),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_45),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_92),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_0),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_112),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_20),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_76),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_37),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_69),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_111),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_116),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_118),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_94),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_171),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_29),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_17),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_105),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_129),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_13),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_135),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_136),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_152),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_57),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_1),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_160),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_134),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_32),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_12),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_109),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_77),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_52),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_34),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_33),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_23),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_170),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_42),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_46),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_54),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_79),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_96),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_119),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_90),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_53),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_11),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_63),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_21),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_8),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_52),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_123),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_103),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_15),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_144),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_7),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_82),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_15),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_44),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_115),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_145),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_89),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_63),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_43),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_38),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_108),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_49),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_100),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_161),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_47),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_51),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_37),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_34),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_146),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_46),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_40),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_14),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_14),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_11),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_27),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_7),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_57),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_75),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_155),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_149),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_164),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_20),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_42),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_173),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_141),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_85),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_13),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_60),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_167),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_38),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_126),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_44),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_6),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_50),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_68),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_153),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_97),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_101),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_172),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_6),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_163),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_99),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_39),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_120),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_10),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_86),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_70),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_47),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_127),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_61),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_48),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_159),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_88),
.Y(n_324)
);

CKINVDCx11_ASAP7_75t_R g325 ( 
.A(n_117),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_55),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_142),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_30),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_98),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_174),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_48),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_54),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_91),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_43),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_87),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_39),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_114),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_45),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_9),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_1),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_16),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_176),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_0),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_30),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_60),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_2),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_107),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_53),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_125),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_67),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_83),
.Y(n_351)
);

BUFx10_ASAP7_75t_L g352 ( 
.A(n_110),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_206),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_277),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_325),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_182),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_238),
.B(n_4),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_206),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_198),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_327),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_277),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_203),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_277),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_277),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_277),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_277),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_199),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_213),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_200),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_202),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_350),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_222),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_200),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_200),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_232),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_232),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_185),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_232),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_261),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_R g380 ( 
.A(n_215),
.B(n_138),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_255),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_255),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_190),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_255),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_260),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_192),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_193),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_260),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_338),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_297),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_201),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_260),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_286),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_204),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_286),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_308),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_286),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_205),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_195),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_338),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_195),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_211),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g403 ( 
.A(n_289),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_196),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_219),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_220),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_226),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_196),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_229),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_350),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_231),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_237),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_234),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_197),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_179),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_218),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_248),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_238),
.B(n_4),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_237),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_242),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_315),
.B(n_178),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_242),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_218),
.Y(n_423)
);

BUFx6f_ASAP7_75t_SL g424 ( 
.A(n_352),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_246),
.Y(n_425)
);

NOR2xp67_ASAP7_75t_L g426 ( 
.A(n_245),
.B(n_5),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_249),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_352),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_246),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_252),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_251),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_258),
.Y(n_432)
);

INVxp33_ASAP7_75t_SL g433 ( 
.A(n_180),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_252),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_218),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_256),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_259),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_267),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_268),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_256),
.Y(n_440)
);

INVx5_ASAP7_75t_L g441 ( 
.A(n_354),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_357),
.A2(n_322),
.B1(n_303),
.B2(n_301),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_361),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_354),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_363),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_421),
.B(n_181),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_361),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_364),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_364),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_360),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_398),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_365),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_415),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_416),
.Y(n_454)
);

AND2x6_ASAP7_75t_L g455 ( 
.A(n_363),
.B(n_225),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_365),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_366),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_366),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_399),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_416),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_423),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_399),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_423),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_401),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_435),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_435),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_369),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_353),
.A2(n_224),
.B1(n_177),
.B2(n_336),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_385),
.B(n_327),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_360),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g471 ( 
.A(n_414),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_369),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_373),
.Y(n_473)
);

OAI21x1_ASAP7_75t_L g474 ( 
.A1(n_418),
.A2(n_275),
.B(n_225),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_389),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_373),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_401),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_374),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_404),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_385),
.B(n_272),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_404),
.Y(n_481)
);

AND2x6_ASAP7_75t_L g482 ( 
.A(n_374),
.B(n_225),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_408),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_375),
.B(n_327),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_400),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_375),
.B(n_333),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_408),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_376),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_412),
.Y(n_489)
);

NOR2x1_ASAP7_75t_L g490 ( 
.A(n_402),
.B(n_333),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_412),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_388),
.B(n_292),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_419),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_388),
.B(n_296),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_376),
.Y(n_495)
);

AND2x6_ASAP7_75t_L g496 ( 
.A(n_378),
.B(n_275),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_419),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_420),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_420),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_392),
.B(n_300),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_378),
.Y(n_501)
);

AND2x2_ASAP7_75t_SL g502 ( 
.A(n_428),
.B(n_275),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_392),
.B(n_302),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_422),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_381),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_381),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_422),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_426),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_382),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_428),
.B(n_352),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_425),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_425),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_353),
.A2(n_273),
.B1(n_247),
.B2(n_216),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_382),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_393),
.B(n_306),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_393),
.B(n_333),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_358),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_446),
.B(n_433),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_446),
.B(n_356),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_444),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_443),
.Y(n_521)
);

BUFx4f_ASAP7_75t_L g522 ( 
.A(n_455),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_444),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_502),
.B(n_377),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_444),
.Y(n_525)
);

INVx4_ASAP7_75t_L g526 ( 
.A(n_461),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_443),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_447),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_445),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_484),
.B(n_342),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_461),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_447),
.Y(n_532)
);

INVx5_ASAP7_75t_L g533 ( 
.A(n_455),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_454),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_445),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_502),
.B(n_383),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_445),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_448),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_442),
.A2(n_362),
.B1(n_403),
.B2(n_368),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_448),
.Y(n_540)
);

NOR2x1p5_ASAP7_75t_L g541 ( 
.A(n_480),
.B(n_355),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_451),
.Y(n_542)
);

AO22x2_ASAP7_75t_L g543 ( 
.A1(n_442),
.A2(n_510),
.B1(n_291),
.B2(n_197),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_449),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_463),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_461),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_449),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_463),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_513),
.A2(n_426),
.B1(n_273),
.B2(n_371),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_463),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_475),
.B(n_358),
.Y(n_551)
);

OR2x6_ASAP7_75t_L g552 ( 
.A(n_490),
.B(n_342),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_450),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_452),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_461),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_475),
.B(n_371),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_465),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_469),
.B(n_395),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_465),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_465),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_502),
.B(n_386),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_469),
.B(n_395),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_452),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_450),
.B(n_387),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_502),
.B(n_391),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_490),
.B(n_394),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_457),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_484),
.A2(n_424),
.B1(n_262),
.B2(n_264),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_457),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_450),
.B(n_405),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_466),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_470),
.B(n_406),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_461),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_466),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_470),
.B(n_407),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_454),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_461),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_466),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_484),
.B(n_342),
.Y(n_579)
);

BUFx2_ASAP7_75t_L g580 ( 
.A(n_517),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_470),
.B(n_409),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_471),
.A2(n_413),
.B1(n_439),
.B2(n_411),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_484),
.B(n_178),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_458),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_458),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_508),
.B(n_417),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_453),
.B(n_431),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_458),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_508),
.B(n_432),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_SL g590 ( 
.A(n_510),
.B(n_424),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_461),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_451),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_453),
.B(n_437),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_471),
.B(n_438),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_480),
.B(n_380),
.Y(n_595)
);

OAI22xp33_ASAP7_75t_L g596 ( 
.A1(n_513),
.A2(n_410),
.B1(n_287),
.B2(n_257),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_492),
.B(n_181),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_471),
.B(n_427),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_484),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_469),
.B(n_397),
.Y(n_600)
);

BUFx10_ASAP7_75t_L g601 ( 
.A(n_485),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_486),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_456),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_492),
.B(n_290),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_494),
.B(n_410),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_494),
.B(n_352),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_516),
.Y(n_607)
);

INVx8_ASAP7_75t_L g608 ( 
.A(n_455),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_517),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_517),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_454),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_454),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_456),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_500),
.B(n_424),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_454),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_456),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_500),
.B(n_290),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_503),
.B(n_515),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_516),
.B(n_397),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_459),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_503),
.B(n_424),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_486),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_456),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_476),
.Y(n_624)
);

AND3x2_ASAP7_75t_L g625 ( 
.A(n_475),
.B(n_291),
.C(n_184),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_516),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_459),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_462),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_476),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_486),
.B(n_384),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_462),
.Y(n_631)
);

NAND3xp33_ASAP7_75t_L g632 ( 
.A(n_515),
.B(n_291),
.C(n_184),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_485),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_486),
.B(n_207),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_486),
.B(n_227),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_476),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_476),
.Y(n_637)
);

BUFx6f_ASAP7_75t_SL g638 ( 
.A(n_455),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_468),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_464),
.Y(n_640)
);

OA22x2_ASAP7_75t_L g641 ( 
.A1(n_474),
.A2(n_294),
.B1(n_278),
.B2(n_270),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_468),
.A2(n_299),
.B1(n_293),
.B2(n_285),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_464),
.Y(n_643)
);

INVx5_ASAP7_75t_L g644 ( 
.A(n_455),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_477),
.Y(n_645)
);

INVx4_ASAP7_75t_SL g646 ( 
.A(n_455),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_478),
.B(n_295),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_478),
.B(n_307),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_477),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_476),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_479),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_476),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_479),
.B(n_359),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_476),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_481),
.B(n_312),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_488),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_474),
.A2(n_294),
.B1(n_262),
.B2(n_264),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_478),
.B(n_481),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_483),
.B(n_317),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_478),
.B(n_318),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_483),
.B(n_384),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_488),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_478),
.B(n_320),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_487),
.Y(n_664)
);

XNOR2xp5_ASAP7_75t_L g665 ( 
.A(n_474),
.B(n_367),
.Y(n_665)
);

NAND2xp33_ASAP7_75t_L g666 ( 
.A(n_455),
.B(n_250),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_487),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_488),
.Y(n_668)
);

INVx4_ASAP7_75t_L g669 ( 
.A(n_514),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_488),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_518),
.B(n_186),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_L g672 ( 
.A1(n_607),
.A2(n_370),
.B1(n_372),
.B2(n_379),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_618),
.B(n_187),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_542),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_607),
.B(n_250),
.Y(n_675)
);

BUFx5_ASAP7_75t_L g676 ( 
.A(n_599),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_521),
.Y(n_677)
);

BUFx5_ASAP7_75t_L g678 ( 
.A(n_599),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_626),
.B(n_183),
.Y(n_679)
);

BUFx2_ASAP7_75t_L g680 ( 
.A(n_580),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_521),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_626),
.B(n_595),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_645),
.B(n_633),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_527),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_630),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_630),
.Y(n_686)
);

INVx1_ASAP7_75t_SL g687 ( 
.A(n_580),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_645),
.B(n_390),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_602),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_519),
.B(n_188),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_667),
.B(n_183),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_558),
.B(n_489),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_594),
.Y(n_693)
);

AND2x6_ASAP7_75t_SL g694 ( 
.A(n_598),
.B(n_265),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_667),
.B(n_597),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_602),
.B(n_250),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_622),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_601),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_622),
.B(n_250),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_633),
.B(n_396),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_604),
.B(n_217),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_640),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_527),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_601),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_587),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_620),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_617),
.B(n_217),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_528),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_576),
.B(n_250),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_620),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_528),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_576),
.B(n_250),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_627),
.Y(n_713)
);

AND2x6_ASAP7_75t_SL g714 ( 
.A(n_653),
.B(n_265),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_532),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_611),
.B(n_221),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_611),
.B(n_280),
.Y(n_717)
);

O2A1O1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_524),
.A2(n_497),
.B(n_512),
.C(n_511),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_536),
.A2(n_310),
.B1(n_330),
.B2(n_349),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_612),
.B(n_221),
.Y(n_720)
);

AND3x1_ASAP7_75t_L g721 ( 
.A(n_549),
.B(n_278),
.C(n_270),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_627),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_586),
.B(n_189),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_534),
.Y(n_724)
);

OAI221xp5_ASAP7_75t_L g725 ( 
.A1(n_549),
.A2(n_311),
.B1(n_339),
.B2(n_328),
.C(n_341),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_522),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_561),
.A2(n_323),
.B1(n_324),
.B2(n_329),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_534),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_592),
.Y(n_729)
);

AO22x2_ASAP7_75t_L g730 ( 
.A1(n_639),
.A2(n_266),
.B1(n_235),
.B2(n_239),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_532),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_612),
.B(n_615),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_615),
.B(n_565),
.Y(n_733)
);

NAND2x1_ASAP7_75t_L g734 ( 
.A(n_534),
.B(n_455),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_538),
.Y(n_735)
);

INVx8_ASAP7_75t_L g736 ( 
.A(n_552),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_614),
.B(n_230),
.Y(n_737)
);

O2A1O1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_605),
.A2(n_498),
.B(n_512),
.C(n_511),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_621),
.B(n_628),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_551),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_628),
.B(n_230),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_631),
.B(n_235),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_631),
.B(n_239),
.Y(n_743)
);

NAND2xp33_ASAP7_75t_L g744 ( 
.A(n_634),
.B(n_335),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_643),
.B(n_244),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_538),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_643),
.B(n_649),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_609),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_641),
.A2(n_288),
.B1(n_284),
.B2(n_281),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_589),
.B(n_191),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_540),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_553),
.B(n_489),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_649),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_581),
.B(n_347),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_539),
.B(n_208),
.C(n_194),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_651),
.B(n_244),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_540),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_651),
.Y(n_758)
);

BUFx8_ASAP7_75t_L g759 ( 
.A(n_551),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_544),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_544),
.Y(n_761)
);

NOR2xp67_ASAP7_75t_L g762 ( 
.A(n_582),
.B(n_491),
.Y(n_762)
);

INVxp67_ASAP7_75t_L g763 ( 
.A(n_556),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_664),
.B(n_263),
.Y(n_764)
);

O2A1O1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_635),
.A2(n_491),
.B(n_493),
.C(n_507),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_564),
.B(n_570),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_664),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_558),
.B(n_263),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_552),
.A2(n_562),
.B1(n_619),
.B2(n_600),
.Y(n_769)
);

OAI221xp5_ASAP7_75t_L g770 ( 
.A1(n_539),
.A2(n_328),
.B1(n_281),
.B2(n_341),
.C(n_344),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_562),
.B(n_266),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_547),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_553),
.B(n_493),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_600),
.B(n_274),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_661),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_661),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_547),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_554),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_619),
.B(n_274),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_554),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_647),
.B(n_309),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_563),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_593),
.B(n_209),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_530),
.B(n_497),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_563),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_567),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_569),
.B(n_310),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_569),
.B(n_313),
.Y(n_788)
);

NOR2x1p5_ASAP7_75t_L g789 ( 
.A(n_610),
.B(n_542),
.Y(n_789)
);

NAND2xp33_ASAP7_75t_L g790 ( 
.A(n_657),
.B(n_351),
.Y(n_790)
);

NOR3xp33_ASAP7_75t_L g791 ( 
.A(n_596),
.B(n_241),
.C(n_243),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_583),
.B(n_313),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_601),
.B(n_498),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_601),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_583),
.B(n_330),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_552),
.A2(n_337),
.B1(n_349),
.B2(n_507),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_566),
.B(n_210),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_545),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_552),
.A2(n_337),
.B1(n_504),
.B2(n_499),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_545),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_552),
.A2(n_590),
.B1(n_543),
.B2(n_530),
.Y(n_801)
);

NAND2xp33_ASAP7_75t_L g802 ( 
.A(n_541),
.B(n_280),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_530),
.B(n_499),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_658),
.B(n_280),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_610),
.B(n_504),
.Y(n_805)
);

INVxp67_ASAP7_75t_SL g806 ( 
.A(n_654),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_530),
.B(n_488),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_579),
.B(n_541),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_522),
.B(n_280),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_579),
.B(n_429),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_641),
.A2(n_284),
.B1(n_288),
.B2(n_311),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_625),
.Y(n_812)
);

AND3x1_ASAP7_75t_L g813 ( 
.A(n_642),
.B(n_332),
.C(n_314),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_568),
.B(n_606),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_572),
.B(n_212),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_575),
.B(n_429),
.Y(n_816)
);

AOI221xp5_ASAP7_75t_L g817 ( 
.A1(n_543),
.A2(n_314),
.B1(n_332),
.B2(n_339),
.C(n_344),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_543),
.A2(n_579),
.B1(n_665),
.B2(n_659),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_543),
.A2(n_455),
.B1(n_482),
.B2(n_496),
.Y(n_819)
);

NOR3xp33_ASAP7_75t_L g820 ( 
.A(n_642),
.B(n_331),
.C(n_326),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_648),
.A2(n_460),
.B(n_509),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_522),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_548),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_579),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_655),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_660),
.B(n_488),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_663),
.B(n_488),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_548),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_550),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_632),
.B(n_514),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_665),
.A2(n_455),
.B1(n_482),
.B2(n_496),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_632),
.B(n_514),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_546),
.B(n_514),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_641),
.A2(n_346),
.B1(n_496),
.B2(n_482),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_669),
.B(n_214),
.Y(n_835)
);

NAND3xp33_ASAP7_75t_L g836 ( 
.A(n_666),
.B(n_340),
.C(n_228),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_638),
.A2(n_496),
.B1(n_482),
.B2(n_506),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_546),
.B(n_514),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_683),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_724),
.A2(n_573),
.B(n_526),
.Y(n_840)
);

OR2x2_ASAP7_75t_L g841 ( 
.A(n_687),
.B(n_430),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_677),
.Y(n_842)
);

BUFx2_ASAP7_75t_L g843 ( 
.A(n_680),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_766),
.B(n_546),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_766),
.B(n_682),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_695),
.B(n_591),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_784),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_671),
.B(n_591),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_726),
.Y(n_849)
);

OAI21xp33_ASAP7_75t_L g850 ( 
.A1(n_671),
.A2(n_233),
.B(n_223),
.Y(n_850)
);

O2A1O1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_733),
.A2(n_584),
.B(n_588),
.C(n_585),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_724),
.A2(n_728),
.B(n_732),
.Y(n_852)
);

BUFx12f_ASAP7_75t_L g853 ( 
.A(n_759),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_681),
.Y(n_854)
);

OAI21xp33_ASAP7_75t_L g855 ( 
.A1(n_690),
.A2(n_240),
.B(n_236),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_726),
.B(n_624),
.Y(n_856)
);

O2A1O1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_733),
.A2(n_584),
.B(n_588),
.C(n_585),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_726),
.Y(n_858)
);

NOR2xp67_ASAP7_75t_L g859 ( 
.A(n_705),
.B(n_693),
.Y(n_859)
);

O2A1O1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_719),
.A2(n_679),
.B(n_770),
.C(n_814),
.Y(n_860)
);

NOR2x1_ASAP7_75t_L g861 ( 
.A(n_789),
.B(n_652),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_818),
.A2(n_670),
.B1(n_652),
.B2(n_656),
.Y(n_862)
);

NAND3xp33_ASAP7_75t_L g863 ( 
.A(n_690),
.B(n_319),
.C(n_253),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_685),
.A2(n_670),
.B1(n_652),
.B2(n_656),
.Y(n_864)
);

BUFx12f_ASAP7_75t_L g865 ( 
.A(n_759),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_739),
.A2(n_624),
.B1(n_636),
.B2(n_668),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_728),
.A2(n_526),
.B(n_573),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_807),
.A2(n_526),
.B(n_573),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_726),
.B(n_629),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_681),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_803),
.A2(n_686),
.B(n_675),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_706),
.B(n_591),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_710),
.B(n_713),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_675),
.A2(n_650),
.B(n_636),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_827),
.A2(n_573),
.B(n_526),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_718),
.A2(n_629),
.B(n_637),
.Y(n_876)
);

A2O1A1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_673),
.A2(n_668),
.B(n_662),
.C(n_650),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_769),
.A2(n_670),
.B1(n_656),
.B2(n_638),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_784),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_722),
.B(n_637),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_822),
.A2(n_608),
.B(n_669),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_822),
.A2(n_608),
.B(n_669),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_822),
.A2(n_608),
.B(n_531),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_723),
.A2(n_638),
.B1(n_662),
.B2(n_608),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_805),
.B(n_434),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_801),
.A2(n_559),
.B1(n_557),
.B2(n_560),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_822),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_740),
.B(n_254),
.Y(n_888)
);

AO21x1_ASAP7_75t_L g889 ( 
.A1(n_737),
.A2(n_809),
.B(n_673),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_753),
.B(n_550),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_758),
.B(n_767),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_676),
.B(n_533),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_816),
.Y(n_893)
);

OAI21xp5_ASAP7_75t_L g894 ( 
.A1(n_709),
.A2(n_613),
.B(n_603),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_780),
.B(n_782),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_786),
.B(n_557),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_684),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_723),
.B(n_559),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_817),
.A2(n_346),
.B1(n_574),
.B2(n_560),
.Y(n_899)
);

AOI21xp33_ASAP7_75t_L g900 ( 
.A1(n_783),
.A2(n_269),
.B(n_271),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_763),
.B(n_276),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_826),
.A2(n_608),
.B(n_531),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_752),
.Y(n_903)
);

NAND2x1p5_ASAP7_75t_L g904 ( 
.A(n_824),
.B(n_533),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_729),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_750),
.B(n_571),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_826),
.A2(n_555),
.B(n_531),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_703),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_750),
.B(n_571),
.Y(n_909)
);

OR2x2_ASAP7_75t_L g910 ( 
.A(n_688),
.B(n_434),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_709),
.A2(n_603),
.B(n_623),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_806),
.A2(n_555),
.B(n_531),
.Y(n_912)
);

NAND2xp33_ASAP7_75t_L g913 ( 
.A(n_676),
.B(n_678),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_773),
.B(n_646),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_712),
.A2(n_613),
.B(n_623),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_702),
.B(n_279),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_747),
.A2(n_555),
.B(n_531),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_810),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_808),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_783),
.A2(n_578),
.B(n_574),
.C(n_616),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_833),
.A2(n_555),
.B(n_577),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_703),
.B(n_578),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_708),
.B(n_711),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_815),
.A2(n_616),
.B(n_520),
.C(n_523),
.Y(n_924)
);

OAI21xp33_ASAP7_75t_L g925 ( 
.A1(n_815),
.A2(n_282),
.B(n_283),
.Y(n_925)
);

NAND3xp33_ASAP7_75t_L g926 ( 
.A(n_797),
.B(n_791),
.C(n_820),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_748),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_838),
.A2(n_555),
.B(n_577),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_708),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_711),
.B(n_520),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_715),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_716),
.A2(n_577),
.B(n_654),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_720),
.A2(n_577),
.B(n_654),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_809),
.A2(n_577),
.B(n_654),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_689),
.A2(n_697),
.B1(n_797),
.B2(n_808),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_692),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_715),
.B(n_731),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_793),
.B(n_298),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_825),
.A2(n_523),
.B1(n_525),
.B2(n_537),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_731),
.B(n_525),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_676),
.B(n_533),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_696),
.A2(n_644),
.B(n_533),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_735),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_735),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_746),
.B(n_529),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_700),
.B(n_775),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_746),
.Y(n_947)
);

BUFx4f_ASAP7_75t_L g948 ( 
.A(n_736),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_751),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_676),
.B(n_678),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_699),
.A2(n_644),
.B(n_533),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_776),
.B(n_304),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_692),
.B(n_646),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_751),
.Y(n_954)
);

O2A1O1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_725),
.A2(n_537),
.B(n_535),
.C(n_529),
.Y(n_955)
);

AOI22x1_ASAP7_75t_L g956 ( 
.A1(n_757),
.A2(n_535),
.B1(n_316),
.B2(n_305),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_762),
.B(n_810),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_765),
.A2(n_321),
.B(n_334),
.C(n_343),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_757),
.B(n_514),
.Y(n_959)
);

INVx2_ASAP7_75t_SL g960 ( 
.A(n_812),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_734),
.A2(n_644),
.B(n_460),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_760),
.B(n_514),
.Y(n_962)
);

NOR2xp67_ASAP7_75t_L g963 ( 
.A(n_674),
.B(n_436),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_749),
.A2(n_482),
.B1(n_496),
.B2(n_345),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_792),
.A2(n_644),
.B(n_460),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_795),
.A2(n_644),
.B(n_460),
.Y(n_966)
);

BUFx12f_ASAP7_75t_L g967 ( 
.A(n_694),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_736),
.Y(n_968)
);

AOI22xp5_ASAP7_75t_L g969 ( 
.A1(n_802),
.A2(n_482),
.B1(n_496),
.B2(n_506),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_790),
.A2(n_473),
.B(n_472),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_760),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_761),
.Y(n_972)
);

NOR3xp33_ASAP7_75t_L g973 ( 
.A(n_672),
.B(n_348),
.C(n_436),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_761),
.B(n_467),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_712),
.A2(n_496),
.B(n_482),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_717),
.A2(n_778),
.B(n_785),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_772),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_738),
.A2(n_440),
.B(n_509),
.C(n_506),
.Y(n_978)
);

AOI22xp33_ASAP7_75t_L g979 ( 
.A1(n_749),
.A2(n_482),
.B1(n_496),
.B2(n_440),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_821),
.A2(n_495),
.B(n_505),
.Y(n_980)
);

INVxp67_ASAP7_75t_L g981 ( 
.A(n_768),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_676),
.B(n_646),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_772),
.A2(n_785),
.B(n_778),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_777),
.A2(n_495),
.B(n_505),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_771),
.A2(n_774),
.B(n_779),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_798),
.Y(n_986)
);

AOI21x1_ASAP7_75t_L g987 ( 
.A1(n_717),
.A2(n_501),
.B(n_467),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_830),
.A2(n_501),
.B(n_467),
.Y(n_988)
);

OAI21x1_ASAP7_75t_L g989 ( 
.A1(n_798),
.A2(n_646),
.B(n_496),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_698),
.B(n_704),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_794),
.B(n_5),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_701),
.A2(n_8),
.B(n_10),
.C(n_17),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_707),
.B(n_496),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_830),
.A2(n_832),
.B(n_744),
.Y(n_994)
);

OAI21x1_ASAP7_75t_L g995 ( 
.A1(n_800),
.A2(n_482),
.B(n_139),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_832),
.A2(n_441),
.B(n_482),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_721),
.B(n_18),
.Y(n_997)
);

AO21x1_ASAP7_75t_L g998 ( 
.A1(n_804),
.A2(n_18),
.B(n_19),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_813),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_676),
.B(n_678),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_781),
.A2(n_441),
.B(n_168),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_799),
.B(n_165),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_755),
.B(n_19),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_754),
.B(n_22),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_691),
.B(n_22),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_741),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_678),
.B(n_441),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_835),
.B(n_441),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_742),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_743),
.A2(n_745),
.B(n_756),
.C(n_764),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_835),
.B(n_441),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_796),
.B(n_162),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_678),
.B(n_441),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_678),
.B(n_831),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_787),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_788),
.B(n_441),
.Y(n_1016)
);

AO21x1_ASAP7_75t_L g1017 ( 
.A1(n_804),
.A2(n_24),
.B(n_25),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_714),
.B(n_26),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_823),
.B(n_829),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_823),
.B(n_27),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_843),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_913),
.A2(n_736),
.B(n_829),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_968),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_1004),
.A2(n_727),
.B(n_819),
.C(n_836),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_845),
.B(n_828),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_968),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_985),
.A2(n_828),
.B(n_834),
.Y(n_1027)
);

O2A1O1Ixp5_ASAP7_75t_L g1028 ( 
.A1(n_889),
.A2(n_730),
.B(n_811),
.C(n_834),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_927),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_981),
.B(n_811),
.Y(n_1030)
);

O2A1O1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_1003),
.A2(n_730),
.B(n_29),
.C(n_31),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_885),
.B(n_903),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_926),
.A2(n_730),
.B1(n_837),
.B2(n_36),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_981),
.B(n_1006),
.Y(n_1034)
);

O2A1O1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_1003),
.A2(n_28),
.B(n_35),
.C(n_36),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_1002),
.A2(n_28),
.B1(n_40),
.B2(n_41),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_1002),
.A2(n_41),
.B1(n_49),
.B2(n_55),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_936),
.B(n_93),
.Y(n_1038)
);

CKINVDCx8_ASAP7_75t_R g1039 ( 
.A(n_968),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_854),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_859),
.B(n_56),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_903),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_893),
.B(n_102),
.Y(n_1043)
);

NAND2x1p5_ASAP7_75t_L g1044 ( 
.A(n_849),
.B(n_858),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_936),
.B(n_80),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_900),
.A2(n_56),
.B(n_58),
.C(n_59),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_1012),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_852),
.A2(n_128),
.B(n_157),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_847),
.B(n_122),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_870),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_950),
.A2(n_121),
.B(n_154),
.Y(n_1051)
);

AOI22x1_ASAP7_75t_L g1052 ( 
.A1(n_994),
.A2(n_78),
.B1(n_151),
.B2(n_148),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_1004),
.A2(n_62),
.B(n_64),
.C(n_65),
.Y(n_1053)
);

BUFx4f_ASAP7_75t_L g1054 ( 
.A(n_853),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_897),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_950),
.A2(n_130),
.B(n_147),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_1000),
.A2(n_1014),
.B(n_867),
.Y(n_1057)
);

OAI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_839),
.A2(n_62),
.B1(n_66),
.B2(n_67),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_905),
.Y(n_1059)
);

AO22x1_ASAP7_75t_L g1060 ( 
.A1(n_1012),
.A2(n_66),
.B1(n_71),
.B2(n_73),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_1000),
.A2(n_131),
.B(n_140),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_973),
.A2(n_158),
.B(n_850),
.C(n_938),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1006),
.B(n_1009),
.Y(n_1063)
);

OAI21xp33_ASAP7_75t_SL g1064 ( 
.A1(n_1014),
.A2(n_891),
.B(n_873),
.Y(n_1064)
);

NOR2xp67_ASAP7_75t_SL g1065 ( 
.A(n_849),
.B(n_858),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_918),
.B(n_953),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1009),
.B(n_938),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_840),
.A2(n_848),
.B(n_875),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_839),
.B(n_895),
.Y(n_1069)
);

BUFx10_ASAP7_75t_L g1070 ( 
.A(n_888),
.Y(n_1070)
);

AOI22xp33_ASAP7_75t_L g1071 ( 
.A1(n_973),
.A2(n_855),
.B1(n_1005),
.B2(n_925),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_844),
.B(n_946),
.Y(n_1072)
);

O2A1O1Ixp33_ASAP7_75t_SL g1073 ( 
.A1(n_958),
.A2(n_877),
.B(n_869),
.C(n_856),
.Y(n_1073)
);

O2A1O1Ixp5_ASAP7_75t_L g1074 ( 
.A1(n_898),
.A2(n_906),
.B(n_909),
.C(n_1011),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_999),
.B(n_888),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_999),
.B(n_901),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_957),
.A2(n_935),
.B1(n_863),
.B2(n_918),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_931),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_SL g1079 ( 
.A1(n_856),
.A2(n_869),
.B(n_982),
.C(n_924),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_901),
.B(n_841),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_SL g1081 ( 
.A1(n_1005),
.A2(n_1010),
.B(n_952),
.C(n_860),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_908),
.B(n_929),
.Y(n_1082)
);

CKINVDCx11_ASAP7_75t_R g1083 ( 
.A(n_865),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_968),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_919),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_847),
.B(n_879),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_944),
.B(n_971),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_919),
.Y(n_1088)
);

O2A1O1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_910),
.A2(n_992),
.B(n_952),
.C(n_1015),
.Y(n_1089)
);

NOR3xp33_ASAP7_75t_SL g1090 ( 
.A(n_1018),
.B(n_916),
.C(n_1020),
.Y(n_1090)
);

AOI21x1_ASAP7_75t_L g1091 ( 
.A1(n_1008),
.A2(n_983),
.B(n_937),
.Y(n_1091)
);

OR2x2_ASAP7_75t_L g1092 ( 
.A(n_960),
.B(n_916),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_879),
.B(n_914),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_977),
.B(n_943),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_914),
.B(n_919),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_953),
.B(n_919),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_947),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_978),
.A2(n_871),
.B(n_846),
.C(n_991),
.Y(n_1098)
);

CKINVDCx14_ASAP7_75t_R g1099 ( 
.A(n_967),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_990),
.B(n_963),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_881),
.A2(n_882),
.B(n_883),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_949),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_902),
.A2(n_868),
.B(n_941),
.Y(n_1103)
);

INVx1_ASAP7_75t_SL g1104 ( 
.A(n_997),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_954),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_861),
.B(n_849),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_972),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_892),
.A2(n_941),
.B(n_923),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_939),
.A2(n_880),
.B(n_920),
.C(n_866),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_892),
.A2(n_917),
.B(n_912),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_986),
.Y(n_1111)
);

O2A1O1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_886),
.A2(n_890),
.B(n_896),
.C(n_872),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_948),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_982),
.A2(n_1007),
.B(n_933),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_849),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_948),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_858),
.B(n_887),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_858),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_899),
.B(n_1019),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1007),
.A2(n_932),
.B(n_928),
.Y(n_1120)
);

AO21x2_ASAP7_75t_L g1121 ( 
.A1(n_876),
.A2(n_976),
.B(n_884),
.Y(n_1121)
);

INVx1_ASAP7_75t_SL g1122 ( 
.A(n_887),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_SL g1123 ( 
.A(n_887),
.B(n_1018),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_921),
.A2(n_907),
.B(n_1013),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_887),
.B(n_862),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_979),
.A2(n_899),
.B1(n_964),
.B2(n_864),
.Y(n_1126)
);

INVx5_ASAP7_75t_L g1127 ( 
.A(n_979),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_964),
.B(n_1017),
.Y(n_1128)
);

NAND2xp33_ASAP7_75t_R g1129 ( 
.A(n_993),
.B(n_940),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_974),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_988),
.A2(n_980),
.B(n_970),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_922),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_904),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_930),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_945),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_934),
.A2(n_962),
.B(n_959),
.Y(n_1136)
);

AO21x2_ASAP7_75t_L g1137 ( 
.A1(n_874),
.A2(n_915),
.B(n_894),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_878),
.B(n_956),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_998),
.A2(n_904),
.B1(n_965),
.B2(n_966),
.Y(n_1139)
);

O2A1O1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_955),
.A2(n_851),
.B(n_857),
.C(n_911),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_989),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_SL g1142 ( 
.A(n_975),
.B(n_1001),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_984),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_987),
.B(n_1016),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_961),
.B(n_942),
.Y(n_1145)
);

AND2x6_ASAP7_75t_L g1146 ( 
.A(n_969),
.B(n_995),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_951),
.B(n_996),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_854),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_854),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_R g1150 ( 
.A(n_905),
.B(n_542),
.Y(n_1150)
);

BUFx8_ASAP7_75t_L g1151 ( 
.A(n_853),
.Y(n_1151)
);

AO21x1_ASAP7_75t_L g1152 ( 
.A1(n_1004),
.A2(n_737),
.B(n_845),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_913),
.A2(n_728),
.B(n_724),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_913),
.A2(n_728),
.B(n_724),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1004),
.A2(n_671),
.B(n_518),
.C(n_766),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_913),
.A2(n_728),
.B(n_724),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_885),
.B(n_683),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_845),
.A2(n_926),
.B1(n_981),
.B2(n_1002),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_845),
.B(n_981),
.Y(n_1159)
);

NAND3xp33_ASAP7_75t_SL g1160 ( 
.A(n_973),
.B(n_518),
.C(n_671),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_845),
.B(n_683),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_842),
.Y(n_1162)
);

INVx2_ASAP7_75t_SL g1163 ( 
.A(n_843),
.Y(n_1163)
);

BUFx8_ASAP7_75t_L g1164 ( 
.A(n_853),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_845),
.B(n_981),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_845),
.B(n_683),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_913),
.A2(n_728),
.B(n_724),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_845),
.B(n_981),
.Y(n_1168)
);

NOR3xp33_ASAP7_75t_SL g1169 ( 
.A(n_1018),
.B(n_610),
.C(n_542),
.Y(n_1169)
);

CKINVDCx14_ASAP7_75t_R g1170 ( 
.A(n_905),
.Y(n_1170)
);

AOI21x1_ASAP7_75t_L g1171 ( 
.A1(n_856),
.A2(n_733),
.B(n_869),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1003),
.A2(n_671),
.B(n_518),
.C(n_900),
.Y(n_1172)
);

AOI221xp5_ASAP7_75t_L g1173 ( 
.A1(n_900),
.A2(n_442),
.B1(n_596),
.B2(n_518),
.C(n_446),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_845),
.B(n_705),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1004),
.A2(n_671),
.B(n_518),
.C(n_766),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_953),
.Y(n_1176)
);

AOI221x1_ASAP7_75t_L g1177 ( 
.A1(n_973),
.A2(n_543),
.B1(n_926),
.B2(n_1004),
.C(n_737),
.Y(n_1177)
);

AO32x2_ASAP7_75t_L g1178 ( 
.A1(n_1033),
.A2(n_1158),
.A3(n_1037),
.B1(n_1036),
.B2(n_1047),
.Y(n_1178)
);

AOI221xp5_ASAP7_75t_L g1179 ( 
.A1(n_1173),
.A2(n_1172),
.B1(n_1155),
.B2(n_1175),
.C(n_1080),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1111),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1153),
.A2(n_1156),
.B(n_1154),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1101),
.A2(n_1110),
.B(n_1114),
.Y(n_1182)
);

AOI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1138),
.A2(n_1091),
.B(n_1057),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_1039),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1066),
.B(n_1113),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1160),
.A2(n_1081),
.B(n_1075),
.C(n_1076),
.Y(n_1186)
);

NAND3xp33_ASAP7_75t_L g1187 ( 
.A(n_1071),
.B(n_1174),
.C(n_1089),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1062),
.A2(n_1024),
.B(n_1064),
.C(n_1067),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1103),
.A2(n_1120),
.B(n_1124),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1136),
.A2(n_1068),
.B(n_1131),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1158),
.A2(n_1090),
.B(n_1077),
.C(n_1041),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1127),
.A2(n_1168),
.B1(n_1159),
.B2(n_1165),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1157),
.B(n_1161),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1131),
.A2(n_1108),
.B(n_1167),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1022),
.A2(n_1171),
.B(n_1141),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1074),
.A2(n_1112),
.B(n_1121),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1141),
.A2(n_1145),
.B(n_1147),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1104),
.B(n_1034),
.Y(n_1198)
);

O2A1O1Ixp33_ASAP7_75t_SL g1199 ( 
.A1(n_1045),
.A2(n_1043),
.B(n_1049),
.C(n_1033),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1053),
.A2(n_1035),
.B(n_1036),
.C(n_1037),
.Y(n_1200)
);

INVx6_ASAP7_75t_L g1201 ( 
.A(n_1021),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_SL g1202 ( 
.A1(n_1031),
.A2(n_1061),
.B(n_1056),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1166),
.B(n_1032),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_1104),
.B(n_1034),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1127),
.A2(n_1030),
.B1(n_1125),
.B2(n_1072),
.Y(n_1205)
);

NOR2x1_ASAP7_75t_R g1206 ( 
.A(n_1083),
.B(n_1116),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1100),
.A2(n_1098),
.B(n_1127),
.C(n_1030),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1121),
.A2(n_1025),
.B(n_1140),
.Y(n_1208)
);

NAND2x1p5_ASAP7_75t_L g1209 ( 
.A(n_1029),
.B(n_1065),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1109),
.A2(n_1127),
.B(n_1027),
.Y(n_1210)
);

AO31x2_ASAP7_75t_L g1211 ( 
.A1(n_1177),
.A2(n_1144),
.A3(n_1126),
.B(n_1048),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1162),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1163),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1069),
.B(n_1063),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1150),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1096),
.B(n_1176),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1063),
.B(n_1134),
.Y(n_1217)
);

AO21x1_ASAP7_75t_L g1218 ( 
.A1(n_1046),
.A2(n_1128),
.B(n_1142),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1073),
.A2(n_1142),
.B(n_1119),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1079),
.A2(n_1126),
.B(n_1137),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1047),
.A2(n_1123),
.B1(n_1058),
.B2(n_1092),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1137),
.A2(n_1130),
.B(n_1132),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1135),
.A2(n_1143),
.B(n_1082),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1087),
.Y(n_1224)
);

O2A1O1Ixp33_ASAP7_75t_SL g1225 ( 
.A1(n_1086),
.A2(n_1087),
.B(n_1094),
.C(n_1093),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1070),
.B(n_1123),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_1059),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1139),
.A2(n_1052),
.B(n_1051),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1097),
.Y(n_1229)
);

OAI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1042),
.A2(n_1054),
.B1(n_1176),
.B2(n_1102),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1070),
.B(n_1107),
.Y(n_1231)
);

OAI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1028),
.A2(n_1146),
.B(n_1148),
.Y(n_1232)
);

AO32x2_ASAP7_75t_L g1233 ( 
.A1(n_1129),
.A2(n_1060),
.A3(n_1146),
.B1(n_1169),
.B2(n_1044),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1040),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1095),
.A2(n_1117),
.B(n_1044),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1050),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1170),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1055),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1038),
.A2(n_1105),
.B(n_1149),
.C(n_1078),
.Y(n_1239)
);

NAND3x1_ASAP7_75t_L g1240 ( 
.A(n_1151),
.B(n_1164),
.C(n_1054),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1146),
.A2(n_1133),
.B(n_1122),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1038),
.B(n_1106),
.Y(n_1242)
);

NAND2x1p5_ASAP7_75t_L g1243 ( 
.A(n_1023),
.B(n_1026),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1106),
.B(n_1088),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1023),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1146),
.A2(n_1133),
.B(n_1122),
.Y(n_1246)
);

AO31x2_ASAP7_75t_L g1247 ( 
.A1(n_1133),
.A2(n_1115),
.A3(n_1085),
.B(n_1088),
.Y(n_1247)
);

NAND2x1p5_ASAP7_75t_L g1248 ( 
.A(n_1026),
.B(n_1084),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_1085),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1085),
.B(n_1088),
.Y(n_1250)
);

AO31x2_ASAP7_75t_L g1251 ( 
.A1(n_1115),
.A2(n_1118),
.A3(n_1084),
.B(n_1026),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1084),
.B(n_1115),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1151),
.A2(n_1164),
.B(n_1099),
.Y(n_1253)
);

AO31x2_ASAP7_75t_L g1254 ( 
.A1(n_1177),
.A2(n_1152),
.A3(n_889),
.B(n_1144),
.Y(n_1254)
);

OA21x2_ASAP7_75t_L g1255 ( 
.A1(n_1177),
.A2(n_1074),
.B(n_1131),
.Y(n_1255)
);

OAI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1155),
.A2(n_1175),
.B(n_1172),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1174),
.B(n_845),
.Y(n_1257)
);

INVxp67_ASAP7_75t_SL g1258 ( 
.A(n_1065),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1101),
.A2(n_1110),
.B(n_1114),
.Y(n_1259)
);

NAND3xp33_ASAP7_75t_L g1260 ( 
.A(n_1155),
.B(n_1175),
.C(n_1172),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1111),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1155),
.A2(n_1175),
.B1(n_845),
.B2(n_1172),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1080),
.B(n_1172),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1174),
.B(n_845),
.Y(n_1264)
);

BUFx10_ASAP7_75t_L g1265 ( 
.A(n_1041),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1111),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1174),
.B(n_705),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1111),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1177),
.A2(n_1152),
.A3(n_889),
.B(n_1144),
.Y(n_1269)
);

NAND3xp33_ASAP7_75t_L g1270 ( 
.A(n_1155),
.B(n_1175),
.C(n_1172),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1080),
.B(n_1172),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1153),
.A2(n_913),
.B(n_728),
.Y(n_1272)
);

BUFx12f_ASAP7_75t_L g1273 ( 
.A(n_1083),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1174),
.B(n_845),
.Y(n_1274)
);

CKINVDCx11_ASAP7_75t_R g1275 ( 
.A(n_1083),
.Y(n_1275)
);

INVx3_ASAP7_75t_L g1276 ( 
.A(n_1133),
.Y(n_1276)
);

A2O1A1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1172),
.A2(n_1175),
.B(n_1155),
.C(n_1173),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1155),
.A2(n_1175),
.B(n_1172),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1111),
.Y(n_1279)
);

BUFx12f_ASAP7_75t_L g1280 ( 
.A(n_1083),
.Y(n_1280)
);

INVx4_ASAP7_75t_SL g1281 ( 
.A(n_1023),
.Y(n_1281)
);

A2O1A1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1172),
.A2(n_1175),
.B(n_1155),
.C(n_1173),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1155),
.A2(n_1175),
.B(n_1172),
.Y(n_1283)
);

CKINVDCx8_ASAP7_75t_R g1284 ( 
.A(n_1029),
.Y(n_1284)
);

AO31x2_ASAP7_75t_L g1285 ( 
.A1(n_1177),
.A2(n_1152),
.A3(n_889),
.B(n_1144),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1101),
.A2(n_1110),
.B(n_1114),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1080),
.B(n_1172),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1021),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1174),
.B(n_845),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1155),
.A2(n_1175),
.B(n_1172),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1150),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1174),
.B(n_705),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1080),
.B(n_1172),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1153),
.A2(n_913),
.B(n_728),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1066),
.B(n_1113),
.Y(n_1295)
);

BUFx10_ASAP7_75t_L g1296 ( 
.A(n_1041),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_SL g1297 ( 
.A(n_1080),
.B(n_1172),
.Y(n_1297)
);

NAND2x1p5_ASAP7_75t_L g1298 ( 
.A(n_1021),
.B(n_1029),
.Y(n_1298)
);

AOI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1138),
.A2(n_1091),
.B(n_1057),
.Y(n_1299)
);

OA21x2_ASAP7_75t_L g1300 ( 
.A1(n_1177),
.A2(n_1074),
.B(n_1131),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1174),
.B(n_845),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1080),
.B(n_1172),
.Y(n_1302)
);

O2A1O1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1155),
.A2(n_1175),
.B(n_1172),
.C(n_1160),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1101),
.A2(n_1110),
.B(n_1114),
.Y(n_1304)
);

NAND3x1_ASAP7_75t_L g1305 ( 
.A(n_1173),
.B(n_1018),
.C(n_820),
.Y(n_1305)
);

AO31x2_ASAP7_75t_L g1306 ( 
.A1(n_1177),
.A2(n_1152),
.A3(n_889),
.B(n_1144),
.Y(n_1306)
);

A2O1A1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1172),
.A2(n_1175),
.B(n_1155),
.C(n_1173),
.Y(n_1307)
);

NOR2xp67_ASAP7_75t_L g1308 ( 
.A(n_1176),
.B(n_981),
.Y(n_1308)
);

NAND3xp33_ASAP7_75t_SL g1309 ( 
.A(n_1173),
.B(n_1172),
.C(n_1155),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1155),
.A2(n_1175),
.B(n_1172),
.Y(n_1310)
);

INVx4_ASAP7_75t_L g1311 ( 
.A(n_1023),
.Y(n_1311)
);

O2A1O1Ixp33_ASAP7_75t_SL g1312 ( 
.A1(n_1155),
.A2(n_1175),
.B(n_1081),
.C(n_1172),
.Y(n_1312)
);

A2O1A1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1172),
.A2(n_1175),
.B(n_1155),
.C(n_1173),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1066),
.B(n_1113),
.Y(n_1314)
);

A2O1A1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1172),
.A2(n_1175),
.B(n_1155),
.C(n_1173),
.Y(n_1315)
);

AOI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1138),
.A2(n_1091),
.B(n_1057),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1174),
.B(n_845),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1153),
.A2(n_913),
.B(n_728),
.Y(n_1318)
);

AOI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1173),
.A2(n_1160),
.B1(n_671),
.B2(n_1155),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1157),
.B(n_683),
.Y(n_1320)
);

O2A1O1Ixp33_ASAP7_75t_SL g1321 ( 
.A1(n_1155),
.A2(n_1175),
.B(n_1081),
.C(n_1172),
.Y(n_1321)
);

INVx2_ASAP7_75t_SL g1322 ( 
.A(n_1021),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1101),
.A2(n_1110),
.B(n_1114),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1174),
.B(n_845),
.Y(n_1324)
);

AOI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1173),
.A2(n_1160),
.B1(n_671),
.B2(n_1155),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1039),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1066),
.B(n_1113),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_1021),
.Y(n_1328)
);

BUFx2_ASAP7_75t_L g1329 ( 
.A(n_1288),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1305),
.A2(n_1309),
.B1(n_1319),
.B2(n_1325),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1267),
.A2(n_1292),
.B1(n_1257),
.B2(n_1289),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1264),
.B(n_1274),
.Y(n_1332)
);

BUFx12f_ASAP7_75t_L g1333 ( 
.A(n_1275),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1179),
.A2(n_1187),
.B1(n_1293),
.B2(n_1297),
.Y(n_1334)
);

INVx2_ASAP7_75t_SL g1335 ( 
.A(n_1201),
.Y(n_1335)
);

NAND2x1p5_ASAP7_75t_L g1336 ( 
.A(n_1226),
.B(n_1241),
.Y(n_1336)
);

BUFx4f_ASAP7_75t_SL g1337 ( 
.A(n_1273),
.Y(n_1337)
);

INVx2_ASAP7_75t_SL g1338 ( 
.A(n_1201),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1187),
.A2(n_1302),
.B1(n_1271),
.B2(n_1287),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1301),
.A2(n_1324),
.B1(n_1317),
.B2(n_1319),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1284),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1320),
.B(n_1242),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1298),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1263),
.A2(n_1270),
.B1(n_1260),
.B2(n_1325),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1213),
.Y(n_1345)
);

OAI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1221),
.A2(n_1260),
.B1(n_1270),
.B2(n_1210),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1256),
.A2(n_1290),
.B1(n_1310),
.B2(n_1283),
.Y(n_1347)
);

CKINVDCx11_ASAP7_75t_R g1348 ( 
.A(n_1280),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1212),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1221),
.A2(n_1191),
.B1(n_1198),
.B2(n_1204),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1184),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1256),
.A2(n_1278),
.B1(n_1283),
.B2(n_1290),
.Y(n_1352)
);

CKINVDCx20_ASAP7_75t_R g1353 ( 
.A(n_1215),
.Y(n_1353)
);

CKINVDCx20_ASAP7_75t_R g1354 ( 
.A(n_1291),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_1237),
.Y(n_1355)
);

INVxp67_ASAP7_75t_SL g1356 ( 
.A(n_1224),
.Y(n_1356)
);

INVx6_ASAP7_75t_L g1357 ( 
.A(n_1184),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1277),
.A2(n_1282),
.B1(n_1313),
.B2(n_1315),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1328),
.Y(n_1359)
);

INVx6_ASAP7_75t_L g1360 ( 
.A(n_1184),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1261),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1216),
.B(n_1185),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1266),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1268),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1279),
.Y(n_1365)
);

CKINVDCx20_ASAP7_75t_R g1366 ( 
.A(n_1322),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1278),
.A2(n_1310),
.B1(n_1262),
.B2(n_1218),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_SL g1368 ( 
.A1(n_1326),
.A2(n_1227),
.B1(n_1231),
.B2(n_1214),
.Y(n_1368)
);

INVxp67_ASAP7_75t_SL g1369 ( 
.A(n_1222),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1205),
.A2(n_1192),
.B1(n_1193),
.B2(n_1203),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1232),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1265),
.A2(n_1296),
.B1(n_1202),
.B2(n_1208),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1307),
.A2(n_1308),
.B1(n_1207),
.B2(n_1217),
.Y(n_1373)
);

INVx5_ASAP7_75t_L g1374 ( 
.A(n_1245),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1265),
.A2(n_1296),
.B1(n_1220),
.B2(n_1219),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1308),
.A2(n_1186),
.B1(n_1188),
.B2(n_1239),
.Y(n_1376)
);

AOI22xp5_ASAP7_75t_SL g1377 ( 
.A1(n_1185),
.A2(n_1327),
.B1(n_1295),
.B2(n_1314),
.Y(n_1377)
);

CKINVDCx11_ASAP7_75t_R g1378 ( 
.A(n_1326),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1229),
.Y(n_1379)
);

CKINVDCx6p67_ASAP7_75t_R g1380 ( 
.A(n_1326),
.Y(n_1380)
);

OAI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1178),
.A2(n_1236),
.B1(n_1238),
.B2(n_1234),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_SL g1382 ( 
.A1(n_1209),
.A2(n_1327),
.B1(n_1314),
.B2(n_1295),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_SL g1383 ( 
.A1(n_1178),
.A2(n_1200),
.B1(n_1303),
.B2(n_1321),
.Y(n_1383)
);

CKINVDCx11_ASAP7_75t_R g1384 ( 
.A(n_1240),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1223),
.A2(n_1178),
.B1(n_1230),
.B2(n_1255),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1255),
.A2(n_1300),
.B1(n_1232),
.B2(n_1196),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1247),
.Y(n_1387)
);

BUFx10_ASAP7_75t_L g1388 ( 
.A(n_1244),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_SL g1389 ( 
.A1(n_1312),
.A2(n_1300),
.B1(n_1253),
.B2(n_1258),
.Y(n_1389)
);

INVx3_ASAP7_75t_SL g1390 ( 
.A(n_1281),
.Y(n_1390)
);

CKINVDCx11_ASAP7_75t_R g1391 ( 
.A(n_1281),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_1243),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1199),
.A2(n_1225),
.B(n_1228),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1247),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1249),
.A2(n_1276),
.B1(n_1235),
.B2(n_1194),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1233),
.A2(n_1190),
.B1(n_1246),
.B2(n_1272),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1276),
.A2(n_1250),
.B1(n_1197),
.B2(n_1311),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1252),
.A2(n_1248),
.B1(n_1311),
.B2(n_1294),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_SL g1399 ( 
.A1(n_1206),
.A2(n_1233),
.B1(n_1181),
.B2(n_1318),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1183),
.A2(n_1316),
.B1(n_1299),
.B2(n_1233),
.Y(n_1400)
);

AOI22xp5_ASAP7_75t_SL g1401 ( 
.A1(n_1206),
.A2(n_1211),
.B1(n_1251),
.B2(n_1306),
.Y(n_1401)
);

OAI21xp5_ASAP7_75t_SL g1402 ( 
.A1(n_1211),
.A2(n_1269),
.B(n_1306),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_SL g1403 ( 
.A1(n_1211),
.A2(n_1189),
.B1(n_1182),
.B2(n_1304),
.Y(n_1403)
);

CKINVDCx14_ASAP7_75t_R g1404 ( 
.A(n_1254),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1259),
.A2(n_1286),
.B1(n_1323),
.B2(n_1195),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1254),
.Y(n_1406)
);

CKINVDCx11_ASAP7_75t_R g1407 ( 
.A(n_1269),
.Y(n_1407)
);

INVx5_ASAP7_75t_L g1408 ( 
.A(n_1285),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1285),
.A2(n_1155),
.B1(n_1175),
.B2(n_1267),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1285),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1180),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1180),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1309),
.A2(n_1173),
.B1(n_1160),
.B2(n_1179),
.Y(n_1413)
);

INVx8_ASAP7_75t_L g1414 ( 
.A(n_1184),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1288),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1210),
.A2(n_913),
.B(n_1153),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_SL g1417 ( 
.A1(n_1267),
.A2(n_1292),
.B1(n_1075),
.B2(n_1076),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1180),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1267),
.A2(n_1155),
.B1(n_1175),
.B2(n_1292),
.Y(n_1419)
);

INVx6_ASAP7_75t_L g1420 ( 
.A(n_1184),
.Y(n_1420)
);

BUFx12f_ASAP7_75t_L g1421 ( 
.A(n_1275),
.Y(n_1421)
);

BUFx3_ASAP7_75t_L g1422 ( 
.A(n_1201),
.Y(n_1422)
);

BUFx10_ASAP7_75t_L g1423 ( 
.A(n_1201),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_SL g1424 ( 
.A1(n_1187),
.A2(n_1036),
.B1(n_1037),
.B2(n_1047),
.Y(n_1424)
);

BUFx2_ASAP7_75t_SL g1425 ( 
.A(n_1284),
.Y(n_1425)
);

CKINVDCx20_ASAP7_75t_R g1426 ( 
.A(n_1275),
.Y(n_1426)
);

BUFx4f_ASAP7_75t_SL g1427 ( 
.A(n_1273),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1201),
.Y(n_1428)
);

INVx8_ASAP7_75t_L g1429 ( 
.A(n_1184),
.Y(n_1429)
);

BUFx10_ASAP7_75t_L g1430 ( 
.A(n_1201),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1201),
.Y(n_1431)
);

CKINVDCx11_ASAP7_75t_R g1432 ( 
.A(n_1275),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1201),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1288),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1267),
.A2(n_1155),
.B1(n_1175),
.B2(n_1292),
.Y(n_1435)
);

CKINVDCx20_ASAP7_75t_R g1436 ( 
.A(n_1275),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1267),
.A2(n_1155),
.B1(n_1175),
.B2(n_1292),
.Y(n_1437)
);

INVx6_ASAP7_75t_L g1438 ( 
.A(n_1184),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1309),
.A2(n_1173),
.B1(n_1160),
.B2(n_1179),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_SL g1440 ( 
.A1(n_1187),
.A2(n_1036),
.B1(n_1037),
.B2(n_1047),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1257),
.B(n_1264),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1288),
.Y(n_1442)
);

INVx6_ASAP7_75t_L g1443 ( 
.A(n_1184),
.Y(n_1443)
);

BUFx8_ASAP7_75t_SL g1444 ( 
.A(n_1273),
.Y(n_1444)
);

CKINVDCx11_ASAP7_75t_R g1445 ( 
.A(n_1275),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1257),
.B(n_1264),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1267),
.A2(n_1155),
.B1(n_1175),
.B2(n_1292),
.Y(n_1447)
);

INVx1_ASAP7_75t_SL g1448 ( 
.A(n_1288),
.Y(n_1448)
);

OAI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1319),
.A2(n_1325),
.B1(n_1036),
.B2(n_1037),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1180),
.Y(n_1450)
);

AOI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1305),
.A2(n_1160),
.B1(n_1173),
.B2(n_518),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1416),
.A2(n_1393),
.B(n_1405),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1406),
.Y(n_1453)
);

OAI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1451),
.A2(n_1439),
.B(n_1413),
.Y(n_1454)
);

INVx3_ASAP7_75t_L g1455 ( 
.A(n_1336),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_L g1456 ( 
.A(n_1417),
.B(n_1331),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1340),
.B(n_1332),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1410),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1387),
.Y(n_1459)
);

INVx3_ASAP7_75t_L g1460 ( 
.A(n_1336),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1394),
.Y(n_1461)
);

INVx2_ASAP7_75t_SL g1462 ( 
.A(n_1388),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1404),
.B(n_1371),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1371),
.B(n_1347),
.Y(n_1464)
);

CKINVDCx20_ASAP7_75t_R g1465 ( 
.A(n_1426),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1408),
.Y(n_1466)
);

CKINVDCx20_ASAP7_75t_R g1467 ( 
.A(n_1436),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1347),
.B(n_1352),
.Y(n_1468)
);

OA21x2_ASAP7_75t_L g1469 ( 
.A1(n_1386),
.A2(n_1402),
.B(n_1367),
.Y(n_1469)
);

AO21x2_ASAP7_75t_L g1470 ( 
.A1(n_1400),
.A2(n_1346),
.B(n_1369),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1369),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1352),
.B(n_1330),
.Y(n_1472)
);

OA21x2_ASAP7_75t_L g1473 ( 
.A1(n_1386),
.A2(n_1367),
.B(n_1385),
.Y(n_1473)
);

AOI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1358),
.A2(n_1346),
.B(n_1373),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1356),
.Y(n_1475)
);

CKINVDCx20_ASAP7_75t_R g1476 ( 
.A(n_1432),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1356),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1441),
.B(n_1446),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1381),
.Y(n_1479)
);

INVx2_ASAP7_75t_SL g1480 ( 
.A(n_1388),
.Y(n_1480)
);

OR2x6_ASAP7_75t_L g1481 ( 
.A(n_1376),
.B(n_1409),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1383),
.B(n_1401),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1395),
.A2(n_1372),
.B(n_1398),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1382),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1334),
.B(n_1413),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1349),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1383),
.B(n_1344),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1343),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1361),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1363),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1364),
.Y(n_1491)
);

BUFx2_ASAP7_75t_L g1492 ( 
.A(n_1365),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1411),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1412),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1418),
.Y(n_1495)
);

INVx3_ASAP7_75t_L g1496 ( 
.A(n_1450),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1379),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1395),
.A2(n_1372),
.B(n_1375),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_1448),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1407),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1399),
.Y(n_1501)
);

INVxp33_ASAP7_75t_L g1502 ( 
.A(n_1342),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1329),
.Y(n_1503)
);

INVx4_ASAP7_75t_L g1504 ( 
.A(n_1374),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1415),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1377),
.B(n_1397),
.Y(n_1506)
);

INVx1_ASAP7_75t_SL g1507 ( 
.A(n_1359),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1403),
.Y(n_1508)
);

BUFx4f_ASAP7_75t_SL g1509 ( 
.A(n_1333),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1375),
.A2(n_1397),
.B(n_1344),
.Y(n_1510)
);

INVxp33_ASAP7_75t_L g1511 ( 
.A(n_1434),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1403),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1385),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1396),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1374),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1334),
.Y(n_1516)
);

BUFx4f_ASAP7_75t_SL g1517 ( 
.A(n_1421),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1350),
.Y(n_1518)
);

OR2x6_ASAP7_75t_L g1519 ( 
.A(n_1368),
.B(n_1447),
.Y(n_1519)
);

OAI21xp33_ASAP7_75t_SL g1520 ( 
.A1(n_1439),
.A2(n_1339),
.B(n_1419),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1442),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1370),
.B(n_1389),
.Y(n_1522)
);

NAND3xp33_ASAP7_75t_SL g1523 ( 
.A(n_1435),
.B(n_1437),
.C(n_1440),
.Y(n_1523)
);

O2A1O1Ixp33_ASAP7_75t_SL g1524 ( 
.A1(n_1449),
.A2(n_1335),
.B(n_1338),
.C(n_1424),
.Y(n_1524)
);

INVx2_ASAP7_75t_SL g1525 ( 
.A(n_1374),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1389),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1449),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1345),
.Y(n_1528)
);

OAI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1362),
.A2(n_1355),
.B(n_1366),
.Y(n_1529)
);

INVx1_ASAP7_75t_SL g1530 ( 
.A(n_1425),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1502),
.B(n_1341),
.Y(n_1531)
);

CKINVDCx16_ASAP7_75t_R g1532 ( 
.A(n_1465),
.Y(n_1532)
);

O2A1O1Ixp33_ASAP7_75t_L g1533 ( 
.A1(n_1454),
.A2(n_1390),
.B(n_1351),
.C(n_1392),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1463),
.B(n_1514),
.Y(n_1534)
);

A2O1A1Ixp33_ASAP7_75t_L g1535 ( 
.A1(n_1474),
.A2(n_1429),
.B(n_1414),
.C(n_1431),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1507),
.B(n_1422),
.Y(n_1536)
);

O2A1O1Ixp33_ASAP7_75t_L g1537 ( 
.A1(n_1520),
.A2(n_1390),
.B(n_1433),
.C(n_1428),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1456),
.A2(n_1380),
.B1(n_1443),
.B2(n_1438),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1492),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1467),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1497),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1457),
.B(n_1414),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1514),
.B(n_1443),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1494),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1497),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1478),
.B(n_1354),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1511),
.B(n_1353),
.Y(n_1547)
);

NAND2xp33_ASAP7_75t_R g1548 ( 
.A(n_1503),
.B(n_1445),
.Y(n_1548)
);

O2A1O1Ixp33_ASAP7_75t_L g1549 ( 
.A1(n_1520),
.A2(n_1384),
.B(n_1391),
.C(n_1378),
.Y(n_1549)
);

OAI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1523),
.A2(n_1485),
.B(n_1481),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1500),
.B(n_1420),
.Y(n_1551)
);

AOI221xp5_ASAP7_75t_L g1552 ( 
.A1(n_1524),
.A2(n_1429),
.B1(n_1438),
.B2(n_1357),
.C(n_1360),
.Y(n_1552)
);

A2O1A1Ixp33_ASAP7_75t_L g1553 ( 
.A1(n_1487),
.A2(n_1438),
.B(n_1357),
.C(n_1360),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1455),
.B(n_1360),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1500),
.B(n_1423),
.Y(n_1555)
);

AO21x1_ASAP7_75t_L g1556 ( 
.A1(n_1487),
.A2(n_1337),
.B(n_1427),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1500),
.B(n_1423),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1455),
.B(n_1430),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1464),
.B(n_1430),
.Y(n_1559)
);

NAND2xp33_ASAP7_75t_L g1560 ( 
.A(n_1472),
.B(n_1427),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1519),
.A2(n_1348),
.B1(n_1444),
.B2(n_1481),
.Y(n_1561)
);

NOR2x1_ASAP7_75t_SL g1562 ( 
.A(n_1481),
.B(n_1519),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1460),
.B(n_1496),
.Y(n_1563)
);

AND2x2_ASAP7_75t_SL g1564 ( 
.A(n_1482),
.B(n_1469),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1469),
.B(n_1496),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1469),
.B(n_1496),
.Y(n_1566)
);

A2O1A1Ixp33_ASAP7_75t_L g1567 ( 
.A1(n_1522),
.A2(n_1510),
.B(n_1518),
.C(n_1482),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_SL g1568 ( 
.A(n_1476),
.B(n_1509),
.Y(n_1568)
);

A2O1A1Ixp33_ASAP7_75t_L g1569 ( 
.A1(n_1522),
.A2(n_1510),
.B(n_1518),
.C(n_1472),
.Y(n_1569)
);

NAND3xp33_ASAP7_75t_L g1570 ( 
.A(n_1519),
.B(n_1516),
.C(n_1518),
.Y(n_1570)
);

AO32x2_ASAP7_75t_L g1571 ( 
.A1(n_1462),
.A2(n_1480),
.A3(n_1525),
.B1(n_1515),
.B2(n_1479),
.Y(n_1571)
);

NAND3xp33_ASAP7_75t_L g1572 ( 
.A(n_1519),
.B(n_1501),
.C(n_1527),
.Y(n_1572)
);

O2A1O1Ixp33_ASAP7_75t_SL g1573 ( 
.A1(n_1527),
.A2(n_1462),
.B(n_1480),
.C(n_1501),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1469),
.B(n_1513),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1508),
.B(n_1512),
.Y(n_1575)
);

AND2x2_ASAP7_75t_SL g1576 ( 
.A(n_1473),
.B(n_1506),
.Y(n_1576)
);

AND2x4_ASAP7_75t_SL g1577 ( 
.A(n_1505),
.B(n_1504),
.Y(n_1577)
);

O2A1O1Ixp33_ASAP7_75t_L g1578 ( 
.A1(n_1519),
.A2(n_1468),
.B(n_1528),
.C(n_1499),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1486),
.B(n_1489),
.Y(n_1579)
);

NAND4xp25_ASAP7_75t_L g1580 ( 
.A(n_1503),
.B(n_1521),
.C(n_1489),
.D(n_1491),
.Y(n_1580)
);

OA21x2_ASAP7_75t_L g1581 ( 
.A1(n_1452),
.A2(n_1498),
.B(n_1483),
.Y(n_1581)
);

AOI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1470),
.A2(n_1471),
.B(n_1477),
.Y(n_1582)
);

NAND2x1p5_ASAP7_75t_L g1583 ( 
.A(n_1471),
.B(n_1475),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1490),
.B(n_1491),
.Y(n_1584)
);

OAI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1484),
.A2(n_1530),
.B1(n_1468),
.B2(n_1506),
.Y(n_1585)
);

OAI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1483),
.A2(n_1498),
.B(n_1452),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1493),
.B(n_1495),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1541),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1565),
.B(n_1566),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1550),
.A2(n_1506),
.B1(n_1484),
.B2(n_1526),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1565),
.B(n_1458),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1563),
.B(n_1466),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1574),
.B(n_1458),
.Y(n_1593)
);

INVxp67_ASAP7_75t_L g1594 ( 
.A(n_1544),
.Y(n_1594)
);

BUFx6f_ASAP7_75t_L g1595 ( 
.A(n_1581),
.Y(n_1595)
);

OAI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1572),
.A2(n_1570),
.B1(n_1484),
.B2(n_1585),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1545),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1576),
.B(n_1459),
.Y(n_1598)
);

OAI221xp5_ASAP7_75t_L g1599 ( 
.A1(n_1549),
.A2(n_1526),
.B1(n_1529),
.B2(n_1521),
.C(n_1473),
.Y(n_1599)
);

INVxp67_ASAP7_75t_SL g1600 ( 
.A(n_1582),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1584),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1564),
.B(n_1461),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1564),
.B(n_1461),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1534),
.B(n_1473),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1539),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1581),
.B(n_1461),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1581),
.B(n_1586),
.Y(n_1607)
);

BUFx12f_ASAP7_75t_L g1608 ( 
.A(n_1540),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1575),
.B(n_1470),
.Y(n_1609)
);

AOI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1561),
.A2(n_1506),
.B1(n_1473),
.B2(n_1470),
.Y(n_1610)
);

BUFx3_ASAP7_75t_L g1611 ( 
.A(n_1577),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1609),
.B(n_1583),
.Y(n_1612)
);

AO22x1_ASAP7_75t_L g1613 ( 
.A1(n_1600),
.A2(n_1558),
.B1(n_1559),
.B2(n_1554),
.Y(n_1613)
);

NOR3xp33_ASAP7_75t_SL g1614 ( 
.A(n_1596),
.B(n_1548),
.C(n_1540),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1597),
.Y(n_1615)
);

OAI31xp33_ASAP7_75t_L g1616 ( 
.A1(n_1599),
.A2(n_1567),
.A3(n_1569),
.B(n_1537),
.Y(n_1616)
);

OAI211xp5_ASAP7_75t_L g1617 ( 
.A1(n_1610),
.A2(n_1578),
.B(n_1567),
.C(n_1533),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1606),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1609),
.B(n_1583),
.Y(n_1619)
);

INVx1_ASAP7_75t_SL g1620 ( 
.A(n_1595),
.Y(n_1620)
);

AND2x2_ASAP7_75t_SL g1621 ( 
.A(n_1610),
.B(n_1560),
.Y(n_1621)
);

NAND2x1p5_ASAP7_75t_L g1622 ( 
.A(n_1595),
.B(n_1607),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1589),
.B(n_1571),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1600),
.B(n_1579),
.Y(n_1624)
);

AO21x2_ASAP7_75t_L g1625 ( 
.A1(n_1607),
.A2(n_1569),
.B(n_1453),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1599),
.B(n_1580),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1589),
.B(n_1571),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1591),
.B(n_1571),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1595),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1595),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1594),
.B(n_1551),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1591),
.B(n_1571),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1595),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1595),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1593),
.B(n_1587),
.Y(n_1635)
);

AOI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1590),
.A2(n_1560),
.B1(n_1573),
.B2(n_1553),
.C(n_1535),
.Y(n_1636)
);

INVx3_ASAP7_75t_L g1637 ( 
.A(n_1592),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1608),
.A2(n_1556),
.B1(n_1559),
.B2(n_1542),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1588),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1588),
.Y(n_1640)
);

INVx3_ASAP7_75t_L g1641 ( 
.A(n_1637),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1623),
.B(n_1601),
.Y(n_1642)
);

INVx4_ASAP7_75t_L g1643 ( 
.A(n_1621),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1640),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1618),
.Y(n_1645)
);

INVx1_ASAP7_75t_SL g1646 ( 
.A(n_1624),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1626),
.B(n_1608),
.Y(n_1647)
);

NAND2xp33_ASAP7_75t_SL g1648 ( 
.A(n_1614),
.B(n_1602),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1618),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1622),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1640),
.Y(n_1651)
);

INVx2_ASAP7_75t_SL g1652 ( 
.A(n_1629),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1639),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1618),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1627),
.B(n_1604),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1624),
.B(n_1594),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1639),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1639),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1640),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1624),
.B(n_1605),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1627),
.B(n_1602),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1635),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1612),
.B(n_1619),
.Y(n_1663)
);

NOR2x1_ASAP7_75t_L g1664 ( 
.A(n_1617),
.B(n_1611),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1628),
.B(n_1603),
.Y(n_1665)
);

AND2x4_ASAP7_75t_L g1666 ( 
.A(n_1637),
.B(n_1598),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1635),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1615),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1635),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1628),
.B(n_1603),
.Y(n_1670)
);

INVx2_ASAP7_75t_SL g1671 ( 
.A(n_1653),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1653),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1663),
.B(n_1612),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1652),
.Y(n_1674)
);

AOI21xp33_ASAP7_75t_SL g1675 ( 
.A1(n_1647),
.A2(n_1532),
.B(n_1626),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1652),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1644),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1661),
.B(n_1628),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1644),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1661),
.B(n_1628),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1661),
.B(n_1632),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1644),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1665),
.B(n_1632),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1664),
.B(n_1631),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1652),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1664),
.B(n_1631),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1656),
.B(n_1612),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1651),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1642),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1665),
.B(n_1632),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1651),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1651),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1659),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1665),
.B(n_1632),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1663),
.B(n_1612),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1642),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1659),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1642),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1657),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1657),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1658),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1658),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1647),
.B(n_1517),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1668),
.Y(n_1704)
);

NOR2x1_ASAP7_75t_L g1705 ( 
.A(n_1643),
.B(n_1617),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1668),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1668),
.Y(n_1707)
);

OAI21xp33_ASAP7_75t_L g1708 ( 
.A1(n_1656),
.A2(n_1614),
.B(n_1617),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1662),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1662),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1667),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1646),
.B(n_1619),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1667),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1678),
.B(n_1643),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1693),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1671),
.Y(n_1716)
);

INVxp67_ASAP7_75t_L g1717 ( 
.A(n_1705),
.Y(n_1717)
);

NAND2x1_ASAP7_75t_L g1718 ( 
.A(n_1705),
.B(n_1643),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1708),
.B(n_1646),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1687),
.B(n_1660),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1671),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1684),
.B(n_1686),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1678),
.B(n_1643),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1680),
.B(n_1643),
.Y(n_1724)
);

NOR2xp67_ASAP7_75t_SL g1725 ( 
.A(n_1675),
.B(n_1608),
.Y(n_1725)
);

AOI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1703),
.A2(n_1648),
.B1(n_1621),
.B2(n_1614),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1680),
.B(n_1681),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1673),
.B(n_1660),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1677),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1675),
.B(n_1619),
.Y(n_1730)
);

NAND2x1p5_ASAP7_75t_L g1731 ( 
.A(n_1672),
.B(n_1621),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1677),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1681),
.B(n_1670),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1683),
.B(n_1690),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1673),
.B(n_1568),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1695),
.B(n_1619),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1693),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1683),
.B(n_1670),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1697),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1697),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1679),
.Y(n_1741)
);

INVx1_ASAP7_75t_SL g1742 ( 
.A(n_1712),
.Y(n_1742)
);

INVx2_ASAP7_75t_SL g1743 ( 
.A(n_1672),
.Y(n_1743)
);

INVx1_ASAP7_75t_SL g1744 ( 
.A(n_1712),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1679),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1690),
.B(n_1670),
.Y(n_1746)
);

AO21x1_ASAP7_75t_L g1747 ( 
.A1(n_1699),
.A2(n_1648),
.B(n_1616),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1695),
.A2(n_1621),
.B1(n_1636),
.B2(n_1625),
.Y(n_1748)
);

NOR3xp33_ASAP7_75t_L g1749 ( 
.A(n_1699),
.B(n_1538),
.C(n_1636),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_SL g1750 ( 
.A(n_1694),
.B(n_1621),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1717),
.B(n_1694),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1729),
.Y(n_1752)
);

OAI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1726),
.A2(n_1638),
.B1(n_1636),
.B2(n_1689),
.Y(n_1753)
);

NAND2xp33_ASAP7_75t_L g1754 ( 
.A(n_1749),
.B(n_1638),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_SL g1755 ( 
.A1(n_1731),
.A2(n_1625),
.B1(n_1562),
.B2(n_1650),
.Y(n_1755)
);

INVxp67_ASAP7_75t_L g1756 ( 
.A(n_1735),
.Y(n_1756)
);

AOI222xp33_ASAP7_75t_L g1757 ( 
.A1(n_1719),
.A2(n_1650),
.B1(n_1698),
.B2(n_1689),
.C1(n_1696),
.C2(n_1701),
.Y(n_1757)
);

AOI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1747),
.A2(n_1625),
.B1(n_1613),
.B2(n_1650),
.Y(n_1758)
);

NOR3xp33_ASAP7_75t_SL g1759 ( 
.A(n_1722),
.B(n_1616),
.C(n_1536),
.Y(n_1759)
);

OAI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1748),
.A2(n_1698),
.B1(n_1696),
.B2(n_1669),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1742),
.B(n_1744),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1714),
.B(n_1655),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1734),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1729),
.Y(n_1764)
);

AOI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1747),
.A2(n_1616),
.B(n_1625),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1720),
.B(n_1669),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1732),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1716),
.B(n_1700),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1732),
.Y(n_1769)
);

OAI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1718),
.A2(n_1701),
.B(n_1700),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1741),
.Y(n_1771)
);

AOI222xp33_ASAP7_75t_L g1772 ( 
.A1(n_1750),
.A2(n_1702),
.B1(n_1613),
.B2(n_1710),
.C1(n_1709),
.C2(n_1713),
.Y(n_1772)
);

OAI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1718),
.A2(n_1702),
.B(n_1622),
.Y(n_1773)
);

AOI22xp33_ASAP7_75t_L g1774 ( 
.A1(n_1725),
.A2(n_1625),
.B1(n_1531),
.B2(n_1546),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1745),
.Y(n_1775)
);

OAI22xp33_ASAP7_75t_SL g1776 ( 
.A1(n_1731),
.A2(n_1622),
.B1(n_1711),
.B2(n_1710),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1763),
.B(n_1716),
.Y(n_1777)
);

AOI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1765),
.A2(n_1731),
.B(n_1730),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1752),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1764),
.Y(n_1780)
);

XNOR2x2_ASAP7_75t_L g1781 ( 
.A(n_1758),
.B(n_1721),
.Y(n_1781)
);

OAI32xp33_ASAP7_75t_L g1782 ( 
.A1(n_1753),
.A2(n_1721),
.A3(n_1728),
.B1(n_1724),
.B2(n_1714),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1763),
.B(n_1725),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1767),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1756),
.B(n_1723),
.Y(n_1785)
);

AOI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1754),
.A2(n_1625),
.B1(n_1743),
.B2(n_1723),
.Y(n_1786)
);

AOI221xp5_ASAP7_75t_L g1787 ( 
.A1(n_1754),
.A2(n_1743),
.B1(n_1724),
.B2(n_1740),
.C(n_1739),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1769),
.Y(n_1788)
);

HB1xp67_ASAP7_75t_L g1789 ( 
.A(n_1761),
.Y(n_1789)
);

AOI222xp33_ASAP7_75t_L g1790 ( 
.A1(n_1774),
.A2(n_1715),
.B1(n_1737),
.B2(n_1736),
.C1(n_1727),
.C2(n_1734),
.Y(n_1790)
);

AND2x4_ASAP7_75t_SL g1791 ( 
.A(n_1759),
.B(n_1555),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1771),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1775),
.Y(n_1793)
);

AO21x1_ASAP7_75t_L g1794 ( 
.A1(n_1770),
.A2(n_1734),
.B(n_1688),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1751),
.B(n_1728),
.Y(n_1795)
);

AO22x2_ASAP7_75t_L g1796 ( 
.A1(n_1760),
.A2(n_1674),
.B1(n_1676),
.B2(n_1685),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1777),
.Y(n_1797)
);

OAI322xp33_ASAP7_75t_SL g1798 ( 
.A1(n_1785),
.A2(n_1768),
.A3(n_1759),
.B1(n_1772),
.B2(n_1757),
.C1(n_1713),
.C2(n_1711),
.Y(n_1798)
);

OAI31xp33_ASAP7_75t_L g1799 ( 
.A1(n_1791),
.A2(n_1778),
.A3(n_1774),
.B(n_1781),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1789),
.B(n_1762),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1794),
.A2(n_1776),
.B(n_1773),
.Y(n_1801)
);

AOI222xp33_ASAP7_75t_L g1802 ( 
.A1(n_1787),
.A2(n_1727),
.B1(n_1746),
.B2(n_1738),
.C1(n_1733),
.C2(n_1709),
.Y(n_1802)
);

OAI211xp5_ASAP7_75t_SL g1803 ( 
.A1(n_1790),
.A2(n_1755),
.B(n_1766),
.C(n_1720),
.Y(n_1803)
);

AO22x1_ASAP7_75t_L g1804 ( 
.A1(n_1783),
.A2(n_1746),
.B1(n_1738),
.B2(n_1733),
.Y(n_1804)
);

INVxp67_ASAP7_75t_L g1805 ( 
.A(n_1795),
.Y(n_1805)
);

AOI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1790),
.A2(n_1625),
.B1(n_1613),
.B2(n_1543),
.Y(n_1806)
);

NOR2x1_ASAP7_75t_L g1807 ( 
.A(n_1779),
.B(n_1682),
.Y(n_1807)
);

INVxp67_ASAP7_75t_SL g1808 ( 
.A(n_1786),
.Y(n_1808)
);

XNOR2xp5_ASAP7_75t_L g1809 ( 
.A(n_1800),
.B(n_1792),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1807),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1805),
.B(n_1793),
.Y(n_1811)
);

INVxp67_ASAP7_75t_L g1812 ( 
.A(n_1808),
.Y(n_1812)
);

NOR3xp33_ASAP7_75t_L g1813 ( 
.A(n_1797),
.B(n_1782),
.C(n_1780),
.Y(n_1813)
);

NAND4xp25_ASAP7_75t_L g1814 ( 
.A(n_1799),
.B(n_1786),
.C(n_1788),
.D(n_1784),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1804),
.Y(n_1815)
);

OA22x2_ASAP7_75t_L g1816 ( 
.A1(n_1806),
.A2(n_1691),
.B1(n_1688),
.B2(n_1682),
.Y(n_1816)
);

NOR2x1_ASAP7_75t_L g1817 ( 
.A(n_1801),
.B(n_1691),
.Y(n_1817)
);

INVxp67_ASAP7_75t_L g1818 ( 
.A(n_1802),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1815),
.B(n_1796),
.Y(n_1819)
);

AOI211xp5_ASAP7_75t_L g1820 ( 
.A1(n_1814),
.A2(n_1803),
.B(n_1798),
.C(n_1796),
.Y(n_1820)
);

AOI221xp5_ASAP7_75t_L g1821 ( 
.A1(n_1814),
.A2(n_1692),
.B1(n_1706),
.B2(n_1704),
.C(n_1707),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1810),
.Y(n_1822)
);

AOI211xp5_ASAP7_75t_L g1823 ( 
.A1(n_1812),
.A2(n_1557),
.B(n_1547),
.C(n_1552),
.Y(n_1823)
);

OAI211xp5_ASAP7_75t_L g1824 ( 
.A1(n_1817),
.A2(n_1676),
.B(n_1674),
.C(n_1685),
.Y(n_1824)
);

AOI31xp33_ASAP7_75t_L g1825 ( 
.A1(n_1820),
.A2(n_1809),
.A3(n_1818),
.B(n_1811),
.Y(n_1825)
);

NAND4xp75_ASAP7_75t_L g1826 ( 
.A(n_1819),
.B(n_1813),
.C(n_1816),
.D(n_1692),
.Y(n_1826)
);

INVx2_ASAP7_75t_SL g1827 ( 
.A(n_1822),
.Y(n_1827)
);

OAI211xp5_ASAP7_75t_SL g1828 ( 
.A1(n_1821),
.A2(n_1535),
.B(n_1706),
.C(n_1704),
.Y(n_1828)
);

AOI221xp5_ASAP7_75t_L g1829 ( 
.A1(n_1824),
.A2(n_1707),
.B1(n_1620),
.B2(n_1630),
.C(n_1633),
.Y(n_1829)
);

OAI221xp5_ASAP7_75t_L g1830 ( 
.A1(n_1823),
.A2(n_1622),
.B1(n_1641),
.B2(n_1553),
.C(n_1620),
.Y(n_1830)
);

A2O1A1Ixp33_ASAP7_75t_L g1831 ( 
.A1(n_1820),
.A2(n_1629),
.B(n_1633),
.C(n_1630),
.Y(n_1831)
);

NOR2x1_ASAP7_75t_L g1832 ( 
.A(n_1826),
.B(n_1641),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1827),
.B(n_1831),
.Y(n_1833)
);

NAND2xp33_ASAP7_75t_L g1834 ( 
.A(n_1825),
.B(n_1829),
.Y(n_1834)
);

NAND4xp75_ASAP7_75t_L g1835 ( 
.A(n_1828),
.B(n_1629),
.C(n_1634),
.D(n_1630),
.Y(n_1835)
);

NOR2x1_ASAP7_75t_L g1836 ( 
.A(n_1830),
.B(n_1641),
.Y(n_1836)
);

AOI32xp33_ASAP7_75t_L g1837 ( 
.A1(n_1834),
.A2(n_1641),
.A3(n_1620),
.B1(n_1666),
.B2(n_1633),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1833),
.B(n_1629),
.Y(n_1838)
);

AOI22x1_ASAP7_75t_L g1839 ( 
.A1(n_1832),
.A2(n_1622),
.B1(n_1649),
.B2(n_1645),
.Y(n_1839)
);

AOI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1838),
.A2(n_1836),
.B1(n_1835),
.B2(n_1634),
.Y(n_1840)
);

OAI22x1_ASAP7_75t_L g1841 ( 
.A1(n_1840),
.A2(n_1839),
.B1(n_1837),
.B2(n_1641),
.Y(n_1841)
);

INVx3_ASAP7_75t_SL g1842 ( 
.A(n_1841),
.Y(n_1842)
);

OAI21x1_ASAP7_75t_L g1843 ( 
.A1(n_1841),
.A2(n_1649),
.B(n_1645),
.Y(n_1843)
);

HB1xp67_ASAP7_75t_L g1844 ( 
.A(n_1843),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1842),
.Y(n_1845)
);

OAI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1845),
.A2(n_1649),
.B(n_1645),
.Y(n_1846)
);

AO22x2_ASAP7_75t_L g1847 ( 
.A1(n_1844),
.A2(n_1649),
.B1(n_1654),
.B2(n_1645),
.Y(n_1847)
);

AOI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1846),
.A2(n_1654),
.B1(n_1629),
.B2(n_1633),
.Y(n_1848)
);

AOI21xp33_ASAP7_75t_L g1849 ( 
.A1(n_1848),
.A2(n_1847),
.B(n_1633),
.Y(n_1849)
);

OAI22xp33_ASAP7_75t_L g1850 ( 
.A1(n_1849),
.A2(n_1654),
.B1(n_1630),
.B2(n_1634),
.Y(n_1850)
);

OAI221xp5_ASAP7_75t_R g1851 ( 
.A1(n_1850),
.A2(n_1654),
.B1(n_1622),
.B2(n_1634),
.C(n_1630),
.Y(n_1851)
);

AOI211xp5_ASAP7_75t_L g1852 ( 
.A1(n_1851),
.A2(n_1488),
.B(n_1634),
.C(n_1573),
.Y(n_1852)
);


endmodule