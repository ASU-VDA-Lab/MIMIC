module fake_jpeg_30796_n_312 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_312);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_31),
.Y(n_62)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_51),
.B(n_52),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_38),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_45),
.Y(n_54)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_55),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_35),
.B1(n_30),
.B2(n_32),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_56),
.A2(n_65),
.B1(n_25),
.B2(n_21),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_49),
.A2(n_32),
.B1(n_24),
.B2(n_31),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_57),
.A2(n_25),
.B1(n_21),
.B2(n_27),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_45),
.B(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_67),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_32),
.B(n_29),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_61),
.B(n_36),
.C(n_19),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_79),
.Y(n_94)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_63),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_30),
.B1(n_37),
.B2(n_22),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_43),
.B(n_34),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_73),
.Y(n_103)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_40),
.B(n_33),
.Y(n_73)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_46),
.A2(n_50),
.B1(n_47),
.B2(n_30),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_83),
.B1(n_26),
.B2(n_25),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_27),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_81),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_40),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_41),
.B(n_33),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_82),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_41),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_41),
.B(n_24),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_30),
.B1(n_31),
.B2(n_24),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_36),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_89),
.Y(n_113)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

AND2x4_ASAP7_75t_SL g89 ( 
.A(n_50),
.B(n_29),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_93),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_95),
.A2(n_107),
.B1(n_112),
.B2(n_116),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_96),
.A2(n_109),
.B1(n_122),
.B2(n_79),
.Y(n_144)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_26),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_120),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_51),
.A2(n_23),
.B1(n_29),
.B2(n_22),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_71),
.A2(n_37),
.B1(n_22),
.B2(n_23),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_110),
.A2(n_117),
.B1(n_87),
.B2(n_84),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_56),
.A2(n_36),
.B1(n_23),
.B2(n_37),
.Y(n_112)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_55),
.A2(n_29),
.B1(n_27),
.B2(n_26),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_88),
.A2(n_36),
.B1(n_21),
.B2(n_19),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_118),
.A2(n_124),
.B(n_69),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_36),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_89),
.A2(n_19),
.B1(n_10),
.B2(n_3),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_121),
.A2(n_123),
.B1(n_17),
.B2(n_16),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_61),
.A2(n_11),
.B1(n_17),
.B2(n_4),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_89),
.A2(n_19),
.B1(n_11),
.B2(n_4),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_83),
.A2(n_19),
.B1(n_10),
.B2(n_4),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_125),
.B(n_127),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_92),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_92),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_129),
.B(n_138),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_58),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_132),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_59),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_102),
.A2(n_70),
.B(n_67),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_142),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_81),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_135),
.B(n_139),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_141),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_103),
.B(n_94),
.C(n_102),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_70),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_101),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_94),
.B(n_76),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_152),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_144),
.A2(n_146),
.B1(n_147),
.B2(n_121),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_149),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_96),
.A2(n_76),
.B1(n_86),
.B2(n_79),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_122),
.A2(n_118),
.B1(n_124),
.B2(n_103),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_98),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_113),
.A2(n_87),
.B(n_75),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_109),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_98),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_151),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_SL g152 ( 
.A(n_97),
.B(n_77),
.C(n_64),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_66),
.C(n_53),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_123),
.C(n_112),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_105),
.B(n_66),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_95),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_113),
.A2(n_84),
.B(n_2),
.C(n_1),
.Y(n_157)
);

NAND5xp2_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_104),
.C(n_2),
.D(n_6),
.E(n_7),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_158),
.A2(n_166),
.B1(n_183),
.B2(n_189),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_178),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_135),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_170),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_144),
.A2(n_129),
.B1(n_127),
.B2(n_147),
.Y(n_166)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

INVx2_ASAP7_75t_R g169 ( 
.A(n_134),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_169),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_156),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_155),
.Y(n_200)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_180),
.B(n_182),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_99),
.C(n_111),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_185),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_132),
.B(n_91),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_130),
.A2(n_152),
.B1(n_146),
.B2(n_125),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_128),
.B(n_100),
.C(n_90),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_12),
.B(n_5),
.Y(n_204)
);

MAJx2_ASAP7_75t_L g188 ( 
.A(n_131),
.B(n_119),
.C(n_104),
.Y(n_188)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_133),
.C(n_142),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_130),
.A2(n_93),
.B1(n_68),
.B2(n_74),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_139),
.B(n_90),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_190),
.B(n_136),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_160),
.A2(n_138),
.B1(n_141),
.B2(n_143),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_170),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_160),
.A2(n_138),
.B1(n_157),
.B2(n_148),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_169),
.A2(n_153),
.B1(n_140),
.B2(n_157),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_200),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_201),
.B(n_160),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_171),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_168),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_204),
.A2(n_186),
.B(n_173),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_183),
.A2(n_153),
.B1(n_140),
.B2(n_115),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_205),
.A2(n_213),
.B1(n_217),
.B2(n_161),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_133),
.Y(n_206)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_166),
.B(n_151),
.Y(n_208)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_208),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_162),
.B(n_149),
.Y(n_209)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_173),
.B(n_15),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_212),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_179),
.A2(n_74),
.B1(n_53),
.B2(n_136),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_187),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_177),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_179),
.A2(n_64),
.B1(n_119),
.B2(n_114),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_172),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_223),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_219),
.A2(n_191),
.B1(n_195),
.B2(n_217),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_188),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_224),
.B(n_225),
.Y(n_254)
);

OA22x2_ASAP7_75t_L g248 ( 
.A1(n_227),
.A2(n_229),
.B1(n_212),
.B2(n_210),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_159),
.B1(n_178),
.B2(n_158),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_164),
.C(n_185),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_236),
.C(n_237),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_193),
.B(n_182),
.Y(n_231)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_231),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_194),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_207),
.Y(n_252)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_174),
.Y(n_234)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_235),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_174),
.C(n_190),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_196),
.B(n_163),
.C(n_180),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_159),
.C(n_189),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_202),
.C(n_207),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_239),
.Y(n_245)
);

NOR4xp25_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_214),
.C(n_211),
.D(n_195),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_246),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_243),
.A2(n_247),
.B1(n_227),
.B2(n_248),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_197),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_244),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_222),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_219),
.A2(n_191),
.B1(n_213),
.B2(n_204),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_237),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_253),
.Y(n_265)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_252),
.Y(n_259)
);

OAI21xp33_ASAP7_75t_L g253 ( 
.A1(n_226),
.A2(n_215),
.B(n_192),
.Y(n_253)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_257),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_221),
.B1(n_238),
.B2(n_218),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_261),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_248),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_247),
.A2(n_225),
.B1(n_234),
.B2(n_236),
.Y(n_263)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_263),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_220),
.Y(n_264)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_264),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_230),
.C(n_223),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_267),
.C(n_268),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_224),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_228),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_243),
.A2(n_256),
.B1(n_245),
.B2(n_244),
.Y(n_271)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_271),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_215),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_250),
.C(n_254),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_281),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_276),
.A2(n_270),
.B1(n_258),
.B2(n_260),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_265),
.Y(n_285)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_262),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_269),
.A2(n_248),
.B(n_241),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_282),
.A2(n_203),
.B(n_5),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_256),
.C(n_257),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_268),
.C(n_265),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_284),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_285),
.B(n_286),
.Y(n_296)
);

AOI322xp5_ASAP7_75t_SL g287 ( 
.A1(n_274),
.A2(n_263),
.A3(n_266),
.B1(n_267),
.B2(n_241),
.C1(n_251),
.C2(n_192),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_287),
.B(n_283),
.Y(n_297)
);

NAND4xp25_ASAP7_75t_SL g288 ( 
.A(n_282),
.B(n_167),
.C(n_203),
.D(n_6),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_15),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_16),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_84),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_278),
.C(n_280),
.Y(n_298)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_292),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_294),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_277),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_298),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_295),
.A2(n_273),
.B1(n_284),
.B2(n_288),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_8),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_296),
.A2(n_279),
.B(n_286),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_302),
.A2(n_289),
.B(n_84),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_295),
.B1(n_285),
.B2(n_290),
.Y(n_304)
);

O2A1O1Ixp33_ASAP7_75t_SL g308 ( 
.A1(n_304),
.A2(n_305),
.B(n_306),
.C(n_301),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_306),
.A2(n_303),
.B(n_300),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_307),
.B(n_308),
.Y(n_309)
);

AOI322xp5_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_8),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_14),
.C2(n_10),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_310),
.A2(n_14),
.B1(n_13),
.B2(n_2),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_13),
.Y(n_312)
);


endmodule