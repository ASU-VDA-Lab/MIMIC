module fake_ibex_863_n_1217 (n_151, n_147, n_85, n_167, n_128, n_208, n_234, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_8, n_118, n_224, n_183, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_14, n_0, n_239, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_80, n_172, n_215, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_92, n_144, n_170, n_213, n_101, n_190, n_113, n_138, n_230, n_96, n_185, n_68, n_117, n_214, n_238, n_79, n_81, n_35, n_159, n_202, n_231, n_158, n_211, n_218, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_19, n_228, n_1217);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_208;
input n_234;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_8;
input n_118;
input n_224;
input n_183;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_14;
input n_0;
input n_239;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_80;
input n_172;
input n_215;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_213;
input n_101;
input n_190;
input n_113;
input n_138;
input n_230;
input n_96;
input n_185;
input n_68;
input n_117;
input n_214;
input n_238;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_218;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_19;
input n_228;

output n_1217;

wire n_1084;
wire n_599;
wire n_778;
wire n_822;
wire n_1042;
wire n_507;
wire n_743;
wire n_1060;
wire n_540;
wire n_754;
wire n_395;
wire n_1104;
wire n_1148;
wire n_992;
wire n_1011;
wire n_756;
wire n_529;
wire n_389;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_1090;
wire n_1110;
wire n_946;
wire n_1196;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_1182;
wire n_926;
wire n_1097;
wire n_1079;
wire n_1031;
wire n_1143;
wire n_328;
wire n_372;
wire n_341;
wire n_293;
wire n_418;
wire n_256;
wire n_510;
wire n_845;
wire n_947;
wire n_981;
wire n_972;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_1067;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_1080;
wire n_1162;
wire n_1199;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_1125;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_432;
wire n_1034;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_412;
wire n_457;
wire n_357;
wire n_494;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_1018;
wire n_1044;
wire n_1106;
wire n_1129;
wire n_449;
wire n_1131;
wire n_547;
wire n_1134;
wire n_727;
wire n_1138;
wire n_1077;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_1174;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_1147;
wire n_542;
wire n_900;
wire n_376;
wire n_1098;
wire n_377;
wire n_584;
wire n_1189;
wire n_531;
wire n_647;
wire n_1187;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_698;
wire n_375;
wire n_317;
wire n_340;
wire n_280;
wire n_708;
wire n_901;
wire n_1096;
wire n_667;
wire n_884;
wire n_1061;
wire n_682;
wire n_850;
wire n_1166;
wire n_1181;
wire n_1140;
wire n_326;
wire n_327;
wire n_879;
wire n_1056;
wire n_723;
wire n_270;
wire n_1144;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_1010;
wire n_1203;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_470;
wire n_276;
wire n_339;
wire n_770;
wire n_965;
wire n_348;
wire n_1109;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_243;
wire n_497;
wire n_287;
wire n_711;
wire n_671;
wire n_876;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_989;
wire n_373;
wire n_1051;
wire n_854;
wire n_1008;
wire n_1193;
wire n_458;
wire n_244;
wire n_1053;
wire n_1112;
wire n_1207;
wire n_343;
wire n_310;
wire n_714;
wire n_1076;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_1172;
wire n_1099;
wire n_598;
wire n_825;
wire n_740;
wire n_1169;
wire n_386;
wire n_549;
wire n_1210;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_1201;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_1055;
wire n_673;
wire n_798;
wire n_732;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_1103;
wire n_1161;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_1177;
wire n_1057;
wire n_1068;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_1184;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_1195;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_1141;
wire n_523;
wire n_694;
wire n_787;
wire n_1075;
wire n_1136;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_1197;
wire n_574;
wire n_1168;
wire n_289;
wire n_716;
wire n_865;
wire n_1130;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_1179;
wire n_1192;
wire n_933;
wire n_1081;
wire n_1153;
wire n_279;
wire n_1037;
wire n_374;
wire n_538;
wire n_464;
wire n_669;
wire n_838;
wire n_987;
wire n_1155;
wire n_750;
wire n_1021;
wire n_746;
wire n_1188;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_1117;
wire n_1191;
wire n_1101;
wire n_518;
wire n_367;
wire n_1052;
wire n_852;
wire n_789;
wire n_1133;
wire n_880;
wire n_654;
wire n_1083;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_1178;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_1211;
wire n_570;
wire n_1116;
wire n_623;
wire n_585;
wire n_1030;
wire n_1094;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_1214;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_487;
wire n_769;
wire n_1137;
wire n_1082;
wire n_660;
wire n_1213;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_980;
wire n_454;
wire n_1070;
wire n_1074;
wire n_777;
wire n_1200;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_1120;
wire n_576;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_1180;
wire n_619;
wire n_1089;
wire n_536;
wire n_1124;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_246;
wire n_442;
wire n_1064;
wire n_1071;
wire n_922;
wire n_1171;
wire n_438;
wire n_851;
wire n_993;
wire n_1028;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_1183;
wire n_253;
wire n_1204;
wire n_300;
wire n_1151;
wire n_1135;
wire n_1146;
wire n_973;
wire n_358;
wire n_771;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_999;
wire n_1092;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_1066;
wire n_245;
wire n_589;
wire n_571;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1062;
wire n_1142;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_1215;
wire n_335;
wire n_413;
wire n_1072;
wire n_263;
wire n_1173;
wire n_1069;
wire n_573;
wire n_1208;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_949;
wire n_1007;
wire n_1126;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_699;
wire n_1063;
wire n_351;
wire n_456;
wire n_368;
wire n_834;
wire n_257;
wire n_1115;
wire n_935;
wire n_869;
wire n_998;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_1054;
wire n_672;
wire n_1100;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_553;
wire n_554;
wire n_1078;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_1170;
wire n_605;
wire n_539;
wire n_392;
wire n_354;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_1049;
wire n_1086;
wire n_763;
wire n_1158;
wire n_745;
wire n_329;
wire n_1149;
wire n_447;
wire n_1176;
wire n_940;
wire n_444;
wire n_562;
wire n_564;
wire n_506;
wire n_868;
wire n_546;
wire n_788;
wire n_1202;
wire n_795;
wire n_1065;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_1160;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_1026;
wire n_1216;
wire n_397;
wire n_283;
wire n_366;
wire n_803;
wire n_894;
wire n_1033;
wire n_1118;
wire n_692;
wire n_627;
wire n_990;
wire n_1198;
wire n_709;
wire n_322;
wire n_499;
wire n_888;
wire n_1087;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_1114;
wire n_409;
wire n_1093;
wire n_582;
wire n_978;
wire n_818;
wire n_1167;
wire n_653;
wire n_1205;
wire n_579;
wire n_899;
wire n_843;
wire n_1019;
wire n_1059;
wire n_902;
wire n_332;
wire n_799;
wire n_1190;
wire n_517;
wire n_744;
wire n_817;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_1107;
wire n_381;
wire n_1073;
wire n_1108;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_1209;
wire n_1111;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_285;
wire n_247;
wire n_379;
wire n_320;
wire n_1128;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_268;
wire n_440;
wire n_858;
wire n_385;
wire n_342;
wire n_414;
wire n_430;
wire n_807;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_1145;
wire n_977;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_1113;
wire n_820;
wire n_805;
wire n_670;
wire n_728;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_1164;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_1175;
wire n_485;
wire n_1139;
wire n_870;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_1212;
wire n_461;
wire n_575;
wire n_313;
wire n_1159;
wire n_1119;
wire n_903;
wire n_1154;
wire n_519;
wire n_345;
wire n_408;
wire n_1085;
wire n_361;
wire n_1095;
wire n_455;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_1091;
wire n_885;
wire n_513;
wire n_588;
wire n_877;
wire n_1121;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_1088;
wire n_896;
wire n_528;
wire n_1005;
wire n_1102;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_1150;
wire n_462;
wire n_1194;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_1165;
wire n_1185;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_897;
wire n_889;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_1122;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_890;
wire n_874;
wire n_921;
wire n_912;
wire n_1105;
wire n_1058;
wire n_1163;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_1123;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_1000;
wire n_984;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_298;
wire n_587;
wire n_1035;
wire n_760;
wire n_1038;
wire n_1157;
wire n_751;
wire n_806;
wire n_1127;
wire n_932;
wire n_1186;
wire n_657;
wire n_764;
wire n_1156;
wire n_1206;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;
wire n_1050;

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_157),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_103),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_115),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_104),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_30),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_100),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_234),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_160),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_131),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_44),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_110),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_164),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_35),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_31),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_91),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_206),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_156),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_28),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_117),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_34),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_158),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_129),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_184),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_230),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_211),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_6),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_4),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_216),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_142),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_215),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_105),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_237),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_155),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_68),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_219),
.B(n_212),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_52),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_165),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_207),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_166),
.Y(n_280)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_203),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_144),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_32),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_217),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_9),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_188),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_114),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_183),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_221),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_61),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_138),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_154),
.B(n_139),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_223),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_193),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_84),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_66),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_65),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_204),
.Y(n_298)
);

BUFx5_ASAP7_75t_L g299 ( 
.A(n_224),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_92),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_52),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_76),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_185),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_36),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_7),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_152),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_32),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_95),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_218),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_53),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_83),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_44),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_21),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_48),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_23),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_111),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_47),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_10),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_18),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_153),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_21),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_43),
.Y(n_322)
);

BUFx2_ASAP7_75t_SL g323 ( 
.A(n_75),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_145),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_151),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_36),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_50),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_123),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_181),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_176),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_228),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_54),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_101),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_64),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_27),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_97),
.Y(n_336)
);

BUFx8_ASAP7_75t_SL g337 ( 
.A(n_14),
.Y(n_337)
);

BUFx5_ASAP7_75t_L g338 ( 
.A(n_135),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_182),
.B(n_63),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_56),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_72),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_133),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_225),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_20),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_202),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_106),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_82),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_65),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_194),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_128),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_130),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_175),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_227),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_47),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_229),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_24),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_174),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_57),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_186),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_231),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_220),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_118),
.Y(n_362)
);

BUFx10_ASAP7_75t_L g363 ( 
.A(n_180),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_39),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_98),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_85),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_9),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_179),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_40),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_240),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_121),
.Y(n_371)
);

BUFx8_ASAP7_75t_SL g372 ( 
.A(n_161),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_132),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_62),
.Y(n_374)
);

NOR2xp67_ASAP7_75t_L g375 ( 
.A(n_64),
.B(n_80),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_79),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_205),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_102),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_120),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_49),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_136),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_18),
.Y(n_382)
);

CKINVDCx14_ASAP7_75t_R g383 ( 
.A(n_69),
.Y(n_383)
);

CKINVDCx14_ASAP7_75t_R g384 ( 
.A(n_82),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_236),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_0),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_99),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_214),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_86),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_25),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_170),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_172),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_50),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_213),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_67),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_168),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_77),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_81),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_226),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_177),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_163),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_89),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_11),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_232),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_247),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_372),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_303),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_378),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_267),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_352),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_300),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_245),
.B(n_274),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_281),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_315),
.B(n_0),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_281),
.Y(n_415)
);

NOR2x1_ASAP7_75t_L g416 ( 
.A(n_391),
.B(n_93),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_300),
.Y(n_417)
);

BUFx12f_ASAP7_75t_L g418 ( 
.A(n_363),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_281),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_383),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_372),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_367),
.B(n_1),
.Y(n_422)
);

BUFx8_ASAP7_75t_L g423 ( 
.A(n_392),
.Y(n_423)
);

BUFx8_ASAP7_75t_L g424 ( 
.A(n_335),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_383),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_378),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_386),
.Y(n_427)
);

OA21x2_ASAP7_75t_L g428 ( 
.A1(n_253),
.A2(n_96),
.B(n_94),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_378),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_281),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_281),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_384),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_281),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_369),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_382),
.Y(n_435)
);

OA21x2_ASAP7_75t_L g436 ( 
.A1(n_253),
.A2(n_271),
.B(n_257),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_382),
.B(n_2),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_397),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_397),
.B(n_4),
.Y(n_439)
);

BUFx8_ASAP7_75t_L g440 ( 
.A(n_390),
.Y(n_440)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_363),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_264),
.B(n_5),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_254),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_363),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_322),
.B(n_5),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_299),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_261),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_246),
.Y(n_448)
);

INVx5_ASAP7_75t_L g449 ( 
.A(n_264),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_337),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_350),
.B(n_8),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_275),
.Y(n_452)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_273),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_283),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_295),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_246),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_299),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_328),
.B(n_11),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_252),
.B(n_107),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_340),
.B(n_12),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_299),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_341),
.B(n_12),
.Y(n_462)
);

OAI22x1_ASAP7_75t_R g463 ( 
.A1(n_255),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_246),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_304),
.Y(n_465)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_330),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_296),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_302),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_299),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_307),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_304),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_310),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_312),
.B(n_13),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_299),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_318),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_332),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_344),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_255),
.Y(n_478)
);

OA21x2_ASAP7_75t_L g479 ( 
.A1(n_257),
.A2(n_109),
.B(n_108),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_290),
.Y(n_480)
);

INVx5_ASAP7_75t_L g481 ( 
.A(n_330),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_299),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_241),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_347),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_290),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_338),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_358),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_338),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_271),
.B(n_16),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_338),
.Y(n_490)
);

BUFx8_ASAP7_75t_L g491 ( 
.A(n_338),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_364),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_343),
.B(n_19),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_437),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_408),
.Y(n_495)
);

NAND2xp33_ASAP7_75t_L g496 ( 
.A(n_425),
.B(n_338),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_411),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_437),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_439),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_409),
.A2(n_407),
.B1(n_410),
.B2(n_405),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_425),
.A2(n_242),
.B1(n_248),
.B2(n_241),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_439),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_491),
.B(n_278),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_436),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_441),
.B(n_251),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_406),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_422),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_422),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_491),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_441),
.B(n_256),
.Y(n_510)
);

OR2x6_ASAP7_75t_L g511 ( 
.A(n_418),
.B(n_323),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_417),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_432),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_422),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_418),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_R g516 ( 
.A(n_406),
.B(n_242),
.Y(n_516)
);

CKINVDCx14_ASAP7_75t_R g517 ( 
.A(n_421),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_413),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_444),
.B(n_259),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_442),
.B(n_458),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_493),
.B(n_293),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_427),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_444),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_412),
.A2(n_248),
.B1(n_288),
.B2(n_262),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_415),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_458),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_419),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_443),
.B(n_308),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_419),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_421),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_451),
.B(n_268),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_453),
.B(n_277),
.Y(n_532)
);

AND2x6_ASAP7_75t_L g533 ( 
.A(n_416),
.B(n_343),
.Y(n_533)
);

OAI22xp33_ASAP7_75t_L g534 ( 
.A1(n_420),
.A2(n_301),
.B1(n_305),
.B2(n_297),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_480),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_450),
.Y(n_536)
);

NAND2xp33_ASAP7_75t_L g537 ( 
.A(n_430),
.B(n_338),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_423),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_447),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_452),
.Y(n_540)
);

OAI22xp33_ASAP7_75t_L g541 ( 
.A1(n_445),
.A2(n_301),
.B1(n_305),
.B2(n_297),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_431),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_449),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_454),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_455),
.Y(n_545)
);

NOR2x1p5_ASAP7_75t_L g546 ( 
.A(n_450),
.B(n_380),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_467),
.B(n_308),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_468),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_433),
.Y(n_549)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_453),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_470),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_472),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_475),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_476),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_477),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_451),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_423),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_433),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_484),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_446),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_408),
.Y(n_561)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_487),
.B(n_334),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_446),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_492),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_423),
.A2(n_294),
.B1(n_345),
.B2(n_298),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_466),
.B(n_435),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_466),
.B(n_285),
.Y(n_567)
);

INVxp33_ASAP7_75t_L g568 ( 
.A(n_414),
.Y(n_568)
);

OAI22xp33_ASAP7_75t_L g569 ( 
.A1(n_478),
.A2(n_366),
.B1(n_314),
.B2(n_389),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_424),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_449),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_438),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_483),
.Y(n_573)
);

INVx5_ASAP7_75t_L g574 ( 
.A(n_449),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_473),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_457),
.Y(n_576)
);

OR2x6_ASAP7_75t_L g577 ( 
.A(n_485),
.B(n_375),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_481),
.B(n_457),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_481),
.B(n_361),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_SL g580 ( 
.A(n_424),
.B(n_298),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_483),
.B(n_311),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_461),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_461),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_428),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_469),
.B(n_388),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_469),
.Y(n_586)
);

OAI22xp33_ASAP7_75t_L g587 ( 
.A1(n_460),
.A2(n_314),
.B1(n_366),
.B2(n_393),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_474),
.B(n_388),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_489),
.A2(n_398),
.B1(n_402),
.B2(n_395),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_474),
.B(n_482),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_486),
.B(n_313),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_462),
.B(n_317),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_486),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_488),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_490),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_440),
.Y(n_596)
);

OAI22xp33_ASAP7_75t_SL g597 ( 
.A1(n_463),
.A2(n_319),
.B1(n_326),
.B2(n_321),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_490),
.B(n_338),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_489),
.B(n_243),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_480),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_456),
.B(n_249),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_456),
.Y(n_602)
);

INVx5_ASAP7_75t_L g603 ( 
.A(n_426),
.Y(n_603)
);

INVx8_ASAP7_75t_L g604 ( 
.A(n_456),
.Y(n_604)
);

INVx4_ASAP7_75t_SL g605 ( 
.A(n_429),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_448),
.B(n_327),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_428),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_448),
.B(n_250),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_428),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_464),
.Y(n_610)
);

AND3x2_ASAP7_75t_L g611 ( 
.A(n_459),
.B(n_362),
.C(n_309),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_464),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_479),
.A2(n_345),
.B1(n_359),
.B2(n_353),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_465),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_497),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_500),
.A2(n_359),
.B1(n_371),
.B2(n_353),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_575),
.B(n_258),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_566),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_520),
.A2(n_479),
.B(n_276),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_568),
.B(n_348),
.Y(n_620)
);

O2A1O1Ixp33_ASAP7_75t_L g621 ( 
.A1(n_613),
.A2(n_403),
.B(n_339),
.C(n_260),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_509),
.B(n_263),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_562),
.B(n_354),
.Y(n_623)
);

NOR3xp33_ASAP7_75t_L g624 ( 
.A(n_597),
.B(n_374),
.C(n_356),
.Y(n_624)
);

CKINVDCx11_ASAP7_75t_R g625 ( 
.A(n_535),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_SL g626 ( 
.A(n_538),
.B(n_371),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_505),
.B(n_265),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_512),
.B(n_376),
.Y(n_628)
);

OR2x2_ASAP7_75t_SL g629 ( 
.A(n_515),
.B(n_379),
.Y(n_629)
);

OAI221xp5_ASAP7_75t_L g630 ( 
.A1(n_589),
.A2(n_556),
.B1(n_599),
.B2(n_544),
.C(n_545),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_592),
.B(n_279),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_539),
.B(n_282),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_SL g633 ( 
.A1(n_580),
.A2(n_381),
.B1(n_385),
.B2(n_379),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_540),
.B(n_287),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_548),
.B(n_306),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_498),
.A2(n_266),
.B1(n_270),
.B2(n_269),
.Y(n_636)
);

AO21x1_ASAP7_75t_L g637 ( 
.A1(n_584),
.A2(n_280),
.B(n_272),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_551),
.B(n_316),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_510),
.B(n_244),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_494),
.A2(n_286),
.B1(n_289),
.B2(n_284),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_507),
.B(n_325),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_531),
.A2(n_514),
.B1(n_508),
.B2(n_499),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_511),
.B(n_557),
.Y(n_643)
);

AND2x6_ASAP7_75t_SL g644 ( 
.A(n_577),
.B(n_291),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_513),
.B(n_336),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_508),
.B(n_526),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_552),
.B(n_342),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_553),
.B(n_351),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_554),
.B(n_555),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_523),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_559),
.B(n_365),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_516),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_511),
.B(n_355),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_519),
.B(n_502),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_564),
.B(n_387),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_521),
.B(n_532),
.Y(n_656)
);

BUFx6f_ASAP7_75t_SL g657 ( 
.A(n_511),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_604),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_567),
.B(n_399),
.Y(n_659)
);

AOI221xp5_ASAP7_75t_L g660 ( 
.A1(n_587),
.A2(n_370),
.B1(n_320),
.B2(n_324),
.C(n_404),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_599),
.B(n_329),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_503),
.B(n_331),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_591),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_581),
.B(n_333),
.Y(n_664)
);

NOR3xp33_ASAP7_75t_L g665 ( 
.A(n_587),
.B(n_349),
.C(n_346),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_533),
.B(n_357),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_504),
.A2(n_377),
.B1(n_368),
.B2(n_360),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_572),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_533),
.B(n_373),
.Y(n_669)
);

NOR3xp33_ASAP7_75t_L g670 ( 
.A(n_534),
.B(n_396),
.C(n_394),
.Y(n_670)
);

INVx4_ASAP7_75t_L g671 ( 
.A(n_604),
.Y(n_671)
);

OAI22xp33_ASAP7_75t_L g672 ( 
.A1(n_577),
.A2(n_400),
.B1(n_401),
.B2(n_292),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_570),
.Y(n_673)
);

BUFx6f_ASAP7_75t_SL g674 ( 
.A(n_577),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_522),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_606),
.Y(n_676)
);

NAND2xp33_ASAP7_75t_L g677 ( 
.A(n_607),
.B(n_590),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_550),
.B(n_471),
.Y(n_678)
);

NOR2xp67_ASAP7_75t_L g679 ( 
.A(n_570),
.B(n_22),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_550),
.B(n_471),
.Y(n_680)
);

INVx8_ASAP7_75t_L g681 ( 
.A(n_596),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_593),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_528),
.B(n_22),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_528),
.A2(n_547),
.B1(n_609),
.B2(n_584),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_496),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_685)
);

OAI21xp5_ASAP7_75t_L g686 ( 
.A1(n_584),
.A2(n_113),
.B(n_112),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_547),
.B(n_116),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_609),
.B(n_119),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_601),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_608),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_594),
.B(n_29),
.Y(n_691)
);

NAND2x1p5_ASAP7_75t_L g692 ( 
.A(n_546),
.B(n_31),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_611),
.Y(n_693)
);

INVx4_ASAP7_75t_L g694 ( 
.A(n_574),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_595),
.B(n_33),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_608),
.Y(n_696)
);

INVxp67_ASAP7_75t_L g697 ( 
.A(n_585),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_585),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_588),
.A2(n_534),
.B1(n_517),
.B2(n_569),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_607),
.A2(n_537),
.B(n_598),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_588),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_518),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_530),
.B(n_122),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_525),
.B(n_124),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_527),
.B(n_125),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_579),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_529),
.B(n_126),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_542),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_543),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_542),
.B(n_127),
.Y(n_710)
);

NOR3xp33_ASAP7_75t_L g711 ( 
.A(n_541),
.B(n_45),
.C(n_46),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_501),
.B(n_46),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_549),
.B(n_134),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_558),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_517),
.B(n_137),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_560),
.A2(n_582),
.B1(n_563),
.B2(n_586),
.Y(n_716)
);

OR2x6_ASAP7_75t_L g717 ( 
.A(n_600),
.B(n_569),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_506),
.B(n_140),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_536),
.B(n_565),
.Y(n_719)
);

O2A1O1Ixp5_ASAP7_75t_L g720 ( 
.A1(n_576),
.A2(n_169),
.B(n_239),
.C(n_238),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_582),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_541),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_583),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_583),
.B(n_141),
.Y(n_724)
);

O2A1O1Ixp5_ASAP7_75t_L g725 ( 
.A1(n_586),
.A2(n_171),
.B(n_235),
.C(n_233),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_610),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_615),
.B(n_535),
.Y(n_727)
);

O2A1O1Ixp5_ASAP7_75t_L g728 ( 
.A1(n_637),
.A2(n_578),
.B(n_543),
.C(n_602),
.Y(n_728)
);

OR2x6_ASAP7_75t_SL g729 ( 
.A(n_673),
.B(n_610),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_623),
.B(n_612),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_663),
.B(n_571),
.Y(n_731)
);

OAI21xp33_ASAP7_75t_L g732 ( 
.A1(n_654),
.A2(n_699),
.B(n_626),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_620),
.B(n_67),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_681),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_658),
.Y(n_735)
);

CKINVDCx20_ASAP7_75t_R g736 ( 
.A(n_625),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_616),
.B(n_70),
.Y(n_737)
);

O2A1O1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_670),
.A2(n_630),
.B(n_621),
.C(n_672),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_628),
.B(n_71),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_681),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_643),
.B(n_72),
.Y(n_741)
);

NAND3xp33_ASAP7_75t_SL g742 ( 
.A(n_652),
.B(n_73),
.C(n_74),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_642),
.B(n_73),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_664),
.A2(n_672),
.B1(n_643),
.B2(n_660),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_711),
.A2(n_603),
.B1(n_614),
.B2(n_561),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_649),
.B(n_661),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_631),
.B(n_645),
.Y(n_747)
);

OAI21xp5_ASAP7_75t_L g748 ( 
.A1(n_688),
.A2(n_603),
.B(n_605),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_668),
.B(n_74),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_711),
.A2(n_712),
.B1(n_618),
.B2(n_667),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_646),
.A2(n_495),
.B(n_614),
.Y(n_751)
);

NAND3xp33_ASAP7_75t_L g752 ( 
.A(n_688),
.B(n_624),
.C(n_719),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_668),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_L g754 ( 
.A1(n_698),
.A2(n_701),
.B1(n_640),
.B2(n_689),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_633),
.B(n_76),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_640),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_671),
.B(n_78),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_675),
.B(n_80),
.Y(n_758)
);

AOI33xp33_ASAP7_75t_L g759 ( 
.A1(n_636),
.A2(n_81),
.A3(n_85),
.B1(n_86),
.B2(n_87),
.B3(n_88),
.Y(n_759)
);

OAI21xp5_ASAP7_75t_L g760 ( 
.A1(n_720),
.A2(n_725),
.B(n_716),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_627),
.B(n_89),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_627),
.B(n_636),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_662),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_763)
);

AOI21xp33_ASAP7_75t_L g764 ( 
.A1(n_639),
.A2(n_90),
.B(n_143),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_717),
.B(n_146),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_706),
.A2(n_147),
.B(n_148),
.Y(n_766)
);

AOI21x1_ASAP7_75t_L g767 ( 
.A1(n_678),
.A2(n_149),
.B(n_150),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_717),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_717),
.Y(n_769)
);

NAND3xp33_ASAP7_75t_L g770 ( 
.A(n_624),
.B(n_159),
.C(n_162),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_653),
.B(n_167),
.Y(n_771)
);

INVx11_ASAP7_75t_L g772 ( 
.A(n_657),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_676),
.Y(n_773)
);

CKINVDCx11_ASAP7_75t_R g774 ( 
.A(n_644),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_693),
.B(n_641),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_694),
.Y(n_776)
);

AOI21xp33_ASAP7_75t_L g777 ( 
.A1(n_666),
.A2(n_173),
.B(n_178),
.Y(n_777)
);

AND2x6_ASAP7_75t_L g778 ( 
.A(n_685),
.B(n_187),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_SL g779 ( 
.A1(n_674),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_779)
);

O2A1O1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_683),
.A2(n_192),
.B(n_195),
.C(n_196),
.Y(n_780)
);

NAND2x1p5_ASAP7_75t_L g781 ( 
.A(n_650),
.B(n_197),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_722),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_655),
.B(n_210),
.Y(n_783)
);

AOI21x1_ASAP7_75t_L g784 ( 
.A1(n_680),
.A2(n_198),
.B(n_199),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_692),
.B(n_200),
.Y(n_785)
);

OAI21xp5_ASAP7_75t_L g786 ( 
.A1(n_720),
.A2(n_201),
.B(n_208),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_622),
.B(n_209),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_659),
.A2(n_651),
.B(n_648),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_632),
.B(n_634),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_709),
.Y(n_790)
);

AND2x2_ASAP7_75t_SL g791 ( 
.A(n_702),
.B(n_708),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_635),
.A2(n_647),
.B(n_638),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_690),
.A2(n_696),
.B1(n_721),
.B2(n_669),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_702),
.A2(n_708),
.B1(n_714),
.B2(n_723),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_714),
.A2(n_629),
.B1(n_695),
.B2(n_691),
.Y(n_795)
);

AND2x2_ASAP7_75t_SL g796 ( 
.A(n_715),
.B(n_718),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_692),
.B(n_726),
.Y(n_797)
);

INVx6_ASAP7_75t_L g798 ( 
.A(n_679),
.Y(n_798)
);

NOR2x1p5_ASAP7_75t_SL g799 ( 
.A(n_682),
.B(n_725),
.Y(n_799)
);

BUFx4f_ASAP7_75t_L g800 ( 
.A(n_703),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_710),
.A2(n_713),
.B(n_724),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_705),
.B(n_707),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_699),
.A2(n_613),
.B1(n_556),
.B2(n_665),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_658),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_667),
.A2(n_697),
.B1(n_684),
.B2(n_613),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_663),
.B(n_575),
.Y(n_806)
);

NOR3xp33_ASAP7_75t_L g807 ( 
.A(n_633),
.B(n_478),
.C(n_597),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_663),
.B(n_575),
.Y(n_808)
);

INVxp67_ASAP7_75t_SL g809 ( 
.A(n_616),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_R g810 ( 
.A(n_625),
.B(n_570),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_619),
.A2(n_677),
.B(n_700),
.Y(n_811)
);

NOR3xp33_ASAP7_75t_L g812 ( 
.A(n_633),
.B(n_478),
.C(n_597),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_619),
.A2(n_677),
.B(n_700),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_619),
.A2(n_677),
.B(n_700),
.Y(n_814)
);

A2O1A1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_654),
.A2(n_656),
.B(n_617),
.C(n_661),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_623),
.B(n_568),
.Y(n_816)
);

O2A1O1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_665),
.A2(n_500),
.B(n_670),
.C(n_630),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_663),
.B(n_575),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_R g819 ( 
.A(n_625),
.B(n_570),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_R g820 ( 
.A(n_625),
.B(n_570),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_663),
.B(n_575),
.Y(n_821)
);

O2A1O1Ixp5_ASAP7_75t_SL g822 ( 
.A1(n_795),
.A2(n_764),
.B(n_786),
.C(n_777),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_809),
.B(n_744),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_727),
.B(n_816),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_821),
.B(n_808),
.Y(n_825)
);

INVx4_ASAP7_75t_L g826 ( 
.A(n_772),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_746),
.A2(n_815),
.B1(n_803),
.B2(n_805),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_818),
.B(n_750),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_773),
.B(n_817),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_738),
.B(n_754),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_754),
.B(n_762),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_740),
.Y(n_832)
);

BUFx12f_ASAP7_75t_L g833 ( 
.A(n_774),
.Y(n_833)
);

OA22x2_ASAP7_75t_L g834 ( 
.A1(n_782),
.A2(n_768),
.B1(n_769),
.B2(n_795),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_792),
.A2(n_789),
.B(n_801),
.Y(n_835)
);

BUFx6f_ASAP7_75t_SL g836 ( 
.A(n_734),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_758),
.Y(n_837)
);

BUFx4_ASAP7_75t_SL g838 ( 
.A(n_736),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_757),
.B(n_735),
.Y(n_839)
);

INVx5_ASAP7_75t_L g840 ( 
.A(n_776),
.Y(n_840)
);

BUFx5_ASAP7_75t_L g841 ( 
.A(n_753),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_805),
.A2(n_791),
.B1(n_794),
.B2(n_752),
.Y(n_842)
);

O2A1O1Ixp5_ASAP7_75t_L g843 ( 
.A1(n_748),
.A2(n_761),
.B(n_800),
.C(n_783),
.Y(n_843)
);

AOI21x1_ASAP7_75t_L g844 ( 
.A1(n_767),
.A2(n_784),
.B(n_751),
.Y(n_844)
);

INVx1_ASAP7_75t_SL g845 ( 
.A(n_731),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_804),
.B(n_739),
.Y(n_846)
);

BUFx12f_ASAP7_75t_L g847 ( 
.A(n_737),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_733),
.B(n_797),
.Y(n_848)
);

AOI211x1_ASAP7_75t_L g849 ( 
.A1(n_756),
.A2(n_770),
.B(n_742),
.C(n_743),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_755),
.B(n_807),
.Y(n_850)
);

AO21x1_ASAP7_75t_L g851 ( 
.A1(n_781),
.A2(n_780),
.B(n_766),
.Y(n_851)
);

CKINVDCx11_ASAP7_75t_R g852 ( 
.A(n_729),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_741),
.B(n_730),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_796),
.A2(n_793),
.B1(n_765),
.B2(n_749),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_776),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_812),
.B(n_775),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_810),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_759),
.B(n_787),
.Y(n_858)
);

NOR2x1_ASAP7_75t_L g859 ( 
.A(n_785),
.B(n_771),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_819),
.B(n_820),
.Y(n_860)
);

OAI21xp5_ASAP7_75t_SL g861 ( 
.A1(n_763),
.A2(n_779),
.B(n_781),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_778),
.B(n_799),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_798),
.B(n_790),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_806),
.B(n_818),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_806),
.B(n_808),
.Y(n_865)
);

AO31x2_ASAP7_75t_L g866 ( 
.A1(n_811),
.A2(n_637),
.A3(n_814),
.B(n_813),
.Y(n_866)
);

BUFx5_ASAP7_75t_L g867 ( 
.A(n_753),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_760),
.A2(n_684),
.B(n_815),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_746),
.A2(n_619),
.B(n_788),
.Y(n_869)
);

AO31x2_ASAP7_75t_L g870 ( 
.A1(n_811),
.A2(n_637),
.A3(n_814),
.B(n_813),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_746),
.A2(n_619),
.B(n_788),
.Y(n_871)
);

INVx4_ASAP7_75t_L g872 ( 
.A(n_772),
.Y(n_872)
);

BUFx2_ASAP7_75t_L g873 ( 
.A(n_740),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_746),
.A2(n_619),
.B(n_788),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_810),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_760),
.A2(n_684),
.B(n_815),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_740),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_806),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_806),
.B(n_808),
.Y(n_879)
);

INVx3_ASAP7_75t_SL g880 ( 
.A(n_740),
.Y(n_880)
);

INVx1_ASAP7_75t_SL g881 ( 
.A(n_806),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_760),
.A2(n_684),
.B(n_815),
.Y(n_882)
);

AOI31xp67_ASAP7_75t_L g883 ( 
.A1(n_802),
.A2(n_687),
.A3(n_705),
.B(n_704),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_760),
.A2(n_684),
.B(n_815),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_815),
.A2(n_732),
.B(n_788),
.C(n_747),
.Y(n_885)
);

BUFx10_ASAP7_75t_L g886 ( 
.A(n_757),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_SL g887 ( 
.A1(n_744),
.A2(n_803),
.B(n_746),
.Y(n_887)
);

BUFx2_ASAP7_75t_L g888 ( 
.A(n_740),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_809),
.B(n_573),
.Y(n_889)
);

INVx5_ASAP7_75t_L g890 ( 
.A(n_757),
.Y(n_890)
);

AO31x2_ASAP7_75t_L g891 ( 
.A1(n_811),
.A2(n_637),
.A3(n_814),
.B(n_813),
.Y(n_891)
);

BUFx2_ASAP7_75t_SL g892 ( 
.A(n_740),
.Y(n_892)
);

AO31x2_ASAP7_75t_L g893 ( 
.A1(n_811),
.A2(n_637),
.A3(n_814),
.B(n_813),
.Y(n_893)
);

O2A1O1Ixp5_ASAP7_75t_L g894 ( 
.A1(n_760),
.A2(n_637),
.B(n_728),
.C(n_811),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_760),
.A2(n_684),
.B(n_815),
.Y(n_895)
);

NOR2xp67_ASAP7_75t_L g896 ( 
.A(n_806),
.B(n_808),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_760),
.A2(n_684),
.B(n_815),
.Y(n_897)
);

OAI22x1_ASAP7_75t_L g898 ( 
.A1(n_803),
.A2(n_616),
.B1(n_565),
.B2(n_524),
.Y(n_898)
);

OAI21x1_ASAP7_75t_L g899 ( 
.A1(n_811),
.A2(n_814),
.B(n_813),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_806),
.B(n_818),
.Y(n_900)
);

OAI21x1_ASAP7_75t_L g901 ( 
.A1(n_811),
.A2(n_814),
.B(n_813),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_811),
.A2(n_814),
.B(n_813),
.Y(n_902)
);

INVx1_ASAP7_75t_SL g903 ( 
.A(n_806),
.Y(n_903)
);

AO31x2_ASAP7_75t_L g904 ( 
.A1(n_811),
.A2(n_637),
.A3(n_814),
.B(n_813),
.Y(n_904)
);

OR2x2_ASAP7_75t_L g905 ( 
.A(n_806),
.B(n_478),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_806),
.B(n_808),
.Y(n_906)
);

NAND3x1_ASAP7_75t_L g907 ( 
.A(n_807),
.B(n_812),
.C(n_670),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_806),
.B(n_818),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_806),
.B(n_818),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_806),
.B(n_818),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_SL g911 ( 
.A(n_757),
.B(n_613),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_806),
.B(n_808),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_760),
.A2(n_684),
.B(n_815),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_740),
.Y(n_914)
);

A2O1A1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_815),
.A2(n_732),
.B(n_788),
.C(n_747),
.Y(n_915)
);

OAI21x1_ASAP7_75t_SL g916 ( 
.A1(n_746),
.A2(n_686),
.B(n_792),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_815),
.A2(n_732),
.B(n_788),
.C(n_747),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_740),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_815),
.A2(n_732),
.B(n_788),
.C(n_747),
.Y(n_919)
);

OA21x2_ASAP7_75t_L g920 ( 
.A1(n_760),
.A2(n_786),
.B(n_686),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_806),
.B(n_818),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_776),
.Y(n_922)
);

NAND3xp33_ASAP7_75t_L g923 ( 
.A(n_745),
.B(n_752),
.C(n_815),
.Y(n_923)
);

INVxp67_ASAP7_75t_L g924 ( 
.A(n_806),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_806),
.Y(n_925)
);

INVx4_ASAP7_75t_L g926 ( 
.A(n_772),
.Y(n_926)
);

BUFx8_ASAP7_75t_L g927 ( 
.A(n_734),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_760),
.A2(n_684),
.B(n_815),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_776),
.Y(n_929)
);

O2A1O1Ixp5_ASAP7_75t_SL g930 ( 
.A1(n_795),
.A2(n_435),
.B(n_434),
.C(n_764),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_809),
.B(n_573),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_806),
.B(n_808),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_806),
.B(n_818),
.Y(n_933)
);

O2A1O1Ixp5_ASAP7_75t_L g934 ( 
.A1(n_760),
.A2(n_637),
.B(n_728),
.C(n_811),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_835),
.A2(n_915),
.B(n_885),
.Y(n_935)
);

AO31x2_ASAP7_75t_L g936 ( 
.A1(n_842),
.A2(n_827),
.A3(n_919),
.B(n_917),
.Y(n_936)
);

BUFx2_ASAP7_75t_R g937 ( 
.A(n_875),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_927),
.Y(n_938)
);

NOR2xp67_ASAP7_75t_L g939 ( 
.A(n_826),
.B(n_872),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_896),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_924),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_925),
.B(n_865),
.Y(n_942)
);

INVxp33_ASAP7_75t_SL g943 ( 
.A(n_838),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_896),
.B(n_906),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_854),
.B(n_862),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_822),
.A2(n_934),
.B(n_894),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_881),
.A2(n_903),
.B1(n_932),
.B2(n_931),
.Y(n_947)
);

OA21x2_ASAP7_75t_L g948 ( 
.A1(n_899),
.A2(n_902),
.B(n_901),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_905),
.B(n_825),
.Y(n_949)
);

NAND2x1p5_ASAP7_75t_L g950 ( 
.A(n_890),
.B(n_840),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_855),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_868),
.A2(n_882),
.B(n_876),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_869),
.A2(n_874),
.B(n_871),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_927),
.Y(n_954)
);

AOI21x1_ASAP7_75t_L g955 ( 
.A1(n_862),
.A2(n_844),
.B(n_851),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_887),
.B(n_827),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_864),
.B(n_900),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_857),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_823),
.B(n_908),
.Y(n_959)
);

NAND2x1p5_ASAP7_75t_L g960 ( 
.A(n_890),
.B(n_840),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_845),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_909),
.Y(n_962)
);

AO21x2_ASAP7_75t_L g963 ( 
.A1(n_882),
.A2(n_895),
.B(n_884),
.Y(n_963)
);

INVxp33_ASAP7_75t_SL g964 ( 
.A(n_852),
.Y(n_964)
);

AO21x2_ASAP7_75t_L g965 ( 
.A1(n_884),
.A2(n_897),
.B(n_895),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_910),
.B(n_921),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_933),
.B(n_824),
.Y(n_967)
);

AOI21xp33_ASAP7_75t_SL g968 ( 
.A1(n_834),
.A2(n_880),
.B(n_898),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_850),
.B(n_828),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_879),
.B(n_912),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_829),
.B(n_830),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_831),
.B(n_842),
.Y(n_972)
);

BUFx2_ASAP7_75t_SL g973 ( 
.A(n_836),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_845),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_897),
.A2(n_913),
.B(n_928),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_892),
.B(n_832),
.Y(n_976)
);

OR2x6_ASAP7_75t_L g977 ( 
.A(n_826),
.B(n_872),
.Y(n_977)
);

INVx6_ASAP7_75t_L g978 ( 
.A(n_926),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_913),
.A2(n_928),
.B(n_923),
.Y(n_979)
);

BUFx6f_ASAP7_75t_SL g980 ( 
.A(n_926),
.Y(n_980)
);

OAI21x1_ASAP7_75t_SL g981 ( 
.A1(n_861),
.A2(n_916),
.B(n_858),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_853),
.B(n_848),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_833),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_886),
.B(n_856),
.Y(n_984)
);

OAI21x1_ASAP7_75t_L g985 ( 
.A1(n_930),
.A2(n_843),
.B(n_920),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_886),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_847),
.B(n_839),
.Y(n_987)
);

CKINVDCx6p67_ASAP7_75t_R g988 ( 
.A(n_836),
.Y(n_988)
);

BUFx2_ASAP7_75t_L g989 ( 
.A(n_914),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_837),
.B(n_911),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_907),
.A2(n_859),
.B(n_883),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_846),
.B(n_849),
.Y(n_992)
);

AOI21x1_ASAP7_75t_L g993 ( 
.A1(n_866),
.A2(n_904),
.B(n_893),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_863),
.Y(n_994)
);

AO31x2_ASAP7_75t_L g995 ( 
.A1(n_866),
.A2(n_893),
.A3(n_904),
.B(n_870),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_866),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_870),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_918),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_922),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_891),
.Y(n_1000)
);

BUFx5_ASAP7_75t_L g1001 ( 
.A(n_841),
.Y(n_1001)
);

AOI21xp33_ASAP7_75t_L g1002 ( 
.A1(n_929),
.A2(n_860),
.B(n_873),
.Y(n_1002)
);

CKINVDCx6p67_ASAP7_75t_R g1003 ( 
.A(n_877),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_841),
.A2(n_867),
.B(n_888),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_924),
.B(n_925),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_878),
.B(n_924),
.Y(n_1006)
);

NAND3xp33_ASAP7_75t_L g1007 ( 
.A(n_889),
.B(n_931),
.C(n_849),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_835),
.A2(n_915),
.B(n_885),
.Y(n_1008)
);

INVx4_ASAP7_75t_L g1009 ( 
.A(n_840),
.Y(n_1009)
);

BUFx12f_ASAP7_75t_L g1010 ( 
.A(n_983),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_967),
.B(n_957),
.Y(n_1011)
);

INVx5_ASAP7_75t_SL g1012 ( 
.A(n_988),
.Y(n_1012)
);

INVxp67_ASAP7_75t_L g1013 ( 
.A(n_1005),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_948),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_948),
.Y(n_1015)
);

OA21x2_ASAP7_75t_L g1016 ( 
.A1(n_953),
.A2(n_946),
.B(n_935),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_959),
.B(n_949),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_944),
.B(n_957),
.Y(n_1018)
);

BUFx2_ASAP7_75t_L g1019 ( 
.A(n_1001),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_944),
.B(n_966),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_966),
.B(n_959),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_961),
.Y(n_1022)
);

BUFx10_ASAP7_75t_L g1023 ( 
.A(n_980),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_950),
.Y(n_1024)
);

AO21x2_ASAP7_75t_L g1025 ( 
.A1(n_946),
.A2(n_953),
.B(n_935),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_968),
.B(n_962),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_961),
.Y(n_1027)
);

INVxp67_ASAP7_75t_SL g1028 ( 
.A(n_974),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_982),
.A2(n_947),
.B1(n_969),
.B2(n_942),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_996),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_943),
.Y(n_1031)
);

AO21x2_ASAP7_75t_L g1032 ( 
.A1(n_1008),
.A2(n_981),
.B(n_985),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_982),
.B(n_969),
.Y(n_1033)
);

HB1xp67_ASAP7_75t_L g1034 ( 
.A(n_974),
.Y(n_1034)
);

OR2x2_ASAP7_75t_L g1035 ( 
.A(n_956),
.B(n_963),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_997),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1000),
.Y(n_1037)
);

BUFx2_ASAP7_75t_SL g1038 ( 
.A(n_980),
.Y(n_1038)
);

AO21x2_ASAP7_75t_L g1039 ( 
.A1(n_1008),
.A2(n_955),
.B(n_979),
.Y(n_1039)
);

INVxp33_ASAP7_75t_L g1040 ( 
.A(n_1006),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_984),
.B(n_976),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_940),
.Y(n_1042)
);

NOR2x1_ASAP7_75t_R g1043 ( 
.A(n_938),
.B(n_954),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_990),
.Y(n_1044)
);

BUFx2_ASAP7_75t_SL g1045 ( 
.A(n_939),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_992),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_956),
.B(n_963),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_999),
.Y(n_1048)
);

INVx5_ASAP7_75t_L g1049 ( 
.A(n_951),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_993),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_943),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1030),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_1022),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_1014),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_1021),
.B(n_941),
.Y(n_1055)
);

OR2x2_ASAP7_75t_L g1056 ( 
.A(n_1035),
.B(n_995),
.Y(n_1056)
);

INVxp67_ASAP7_75t_SL g1057 ( 
.A(n_1015),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_1027),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1036),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_1050),
.B(n_1032),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_1029),
.A2(n_1007),
.B1(n_971),
.B2(n_972),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_1046),
.B(n_965),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_1035),
.B(n_952),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1047),
.B(n_975),
.Y(n_1064)
);

INVx1_ASAP7_75t_SL g1065 ( 
.A(n_1048),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_1033),
.A2(n_945),
.B1(n_970),
.B2(n_975),
.Y(n_1066)
);

NOR2xp67_ASAP7_75t_L g1067 ( 
.A(n_1049),
.B(n_1004),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_1019),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1037),
.B(n_936),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_SL g1070 ( 
.A(n_1023),
.Y(n_1070)
);

HB1xp67_ASAP7_75t_L g1071 ( 
.A(n_1034),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_1025),
.B(n_1016),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_1025),
.B(n_936),
.Y(n_1073)
);

INVxp67_ASAP7_75t_SL g1074 ( 
.A(n_1028),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_1042),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_1025),
.B(n_936),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1054),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_1061),
.A2(n_1020),
.B1(n_1018),
.B2(n_1017),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1052),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1052),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1063),
.B(n_1044),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_1060),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1069),
.B(n_1016),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_1065),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1063),
.B(n_1064),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1069),
.B(n_1016),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_1075),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1069),
.B(n_1016),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1063),
.B(n_1039),
.Y(n_1089)
);

INVxp67_ASAP7_75t_SL g1090 ( 
.A(n_1057),
.Y(n_1090)
);

OR2x2_ASAP7_75t_L g1091 ( 
.A(n_1056),
.B(n_1039),
.Y(n_1091)
);

NOR2x1_ASAP7_75t_L g1092 ( 
.A(n_1067),
.B(n_1045),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_1064),
.B(n_1039),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1064),
.B(n_1073),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1073),
.B(n_1032),
.Y(n_1095)
);

NOR2x1_ASAP7_75t_SL g1096 ( 
.A(n_1059),
.B(n_1045),
.Y(n_1096)
);

INVx2_ASAP7_75t_SL g1097 ( 
.A(n_1068),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_1068),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1079),
.Y(n_1099)
);

INVx4_ASAP7_75t_L g1100 ( 
.A(n_1098),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1079),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1080),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1094),
.B(n_1076),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1094),
.B(n_1076),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1094),
.B(n_1062),
.Y(n_1105)
);

INVxp67_ASAP7_75t_SL g1106 ( 
.A(n_1090),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1085),
.B(n_1089),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_1087),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1077),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1083),
.B(n_1072),
.Y(n_1110)
);

INVxp67_ASAP7_75t_L g1111 ( 
.A(n_1098),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1085),
.B(n_1062),
.Y(n_1112)
);

NOR2x1_ASAP7_75t_L g1113 ( 
.A(n_1092),
.B(n_1038),
.Y(n_1113)
);

OR2x2_ASAP7_75t_L g1114 ( 
.A(n_1091),
.B(n_1056),
.Y(n_1114)
);

OR2x2_ASAP7_75t_L g1115 ( 
.A(n_1091),
.B(n_1081),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1083),
.B(n_1072),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1083),
.B(n_1072),
.Y(n_1117)
);

INVxp67_ASAP7_75t_SL g1118 ( 
.A(n_1090),
.Y(n_1118)
);

OR2x2_ASAP7_75t_L g1119 ( 
.A(n_1091),
.B(n_1056),
.Y(n_1119)
);

INVxp67_ASAP7_75t_L g1120 ( 
.A(n_1108),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1103),
.B(n_1089),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1099),
.Y(n_1122)
);

AO22x1_ASAP7_75t_L g1123 ( 
.A1(n_1113),
.A2(n_964),
.B1(n_1092),
.B2(n_1074),
.Y(n_1123)
);

AOI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1113),
.A2(n_1078),
.B1(n_1026),
.B2(n_1061),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1099),
.Y(n_1125)
);

INVxp67_ASAP7_75t_L g1126 ( 
.A(n_1115),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1101),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_1100),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_SL g1129 ( 
.A(n_1100),
.B(n_964),
.Y(n_1129)
);

NOR2xp67_ASAP7_75t_L g1130 ( 
.A(n_1100),
.B(n_1097),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1109),
.Y(n_1131)
);

OR2x2_ASAP7_75t_L g1132 ( 
.A(n_1115),
.B(n_1095),
.Y(n_1132)
);

OR2x2_ASAP7_75t_L g1133 ( 
.A(n_1110),
.B(n_1095),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1109),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1101),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1102),
.Y(n_1136)
);

NAND3xp33_ASAP7_75t_SL g1137 ( 
.A(n_1100),
.B(n_1031),
.C(n_1051),
.Y(n_1137)
);

OR2x2_ASAP7_75t_L g1138 ( 
.A(n_1110),
.B(n_1095),
.Y(n_1138)
);

INVx1_ASAP7_75t_SL g1139 ( 
.A(n_1114),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1103),
.B(n_1093),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_1139),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1131),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1124),
.A2(n_1078),
.B1(n_1119),
.B2(n_1114),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1126),
.B(n_1104),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1131),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_1129),
.A2(n_1055),
.B1(n_1104),
.B2(n_1107),
.Y(n_1146)
);

INVxp67_ASAP7_75t_L g1147 ( 
.A(n_1137),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1122),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1134),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1133),
.B(n_1116),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1133),
.B(n_1138),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1130),
.A2(n_1119),
.B1(n_1105),
.B2(n_1107),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1132),
.A2(n_1093),
.B1(n_1088),
.B2(n_1086),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1134),
.Y(n_1154)
);

AOI31xp33_ASAP7_75t_L g1155 ( 
.A1(n_1123),
.A2(n_1043),
.A3(n_1031),
.B(n_1106),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1125),
.Y(n_1156)
);

AOI211xp5_ASAP7_75t_L g1157 ( 
.A1(n_1128),
.A2(n_1111),
.B(n_1118),
.C(n_1055),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1120),
.A2(n_1111),
.B(n_1074),
.Y(n_1158)
);

NOR2x1_ASAP7_75t_L g1159 ( 
.A(n_1128),
.B(n_1038),
.Y(n_1159)
);

INVxp67_ASAP7_75t_SL g1160 ( 
.A(n_1128),
.Y(n_1160)
);

OAI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1155),
.A2(n_1138),
.B1(n_1132),
.B2(n_1121),
.Y(n_1161)
);

XOR2x2_ASAP7_75t_L g1162 ( 
.A(n_1146),
.B(n_1096),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1159),
.A2(n_1096),
.B(n_1116),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1156),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1143),
.A2(n_1093),
.B1(n_1086),
.B2(n_1088),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1156),
.Y(n_1166)
);

AOI221xp5_ASAP7_75t_L g1167 ( 
.A1(n_1152),
.A2(n_1140),
.B1(n_1117),
.B2(n_1013),
.C(n_1127),
.Y(n_1167)
);

OAI211xp5_ASAP7_75t_SL g1168 ( 
.A1(n_1147),
.A2(n_1002),
.B(n_1066),
.C(n_991),
.Y(n_1168)
);

O2A1O1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1141),
.A2(n_1058),
.B(n_1071),
.C(n_1053),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1157),
.A2(n_1117),
.B1(n_1112),
.B2(n_1105),
.Y(n_1170)
);

OAI211xp5_ASAP7_75t_SL g1171 ( 
.A1(n_1161),
.A2(n_1153),
.B(n_1158),
.C(n_1160),
.Y(n_1171)
);

OAI21xp33_ASAP7_75t_L g1172 ( 
.A1(n_1165),
.A2(n_1151),
.B(n_1144),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1163),
.B(n_1151),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_1169),
.B(n_1150),
.Y(n_1174)
);

AOI221xp5_ASAP7_75t_L g1175 ( 
.A1(n_1167),
.A2(n_1148),
.B1(n_1150),
.B2(n_1142),
.C(n_1154),
.Y(n_1175)
);

AOI221xp5_ASAP7_75t_L g1176 ( 
.A1(n_1170),
.A2(n_1154),
.B1(n_1145),
.B2(n_1142),
.C(n_1135),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1168),
.A2(n_1086),
.B1(n_1088),
.B2(n_1082),
.Y(n_1177)
);

O2A1O1Ixp5_ASAP7_75t_L g1178 ( 
.A1(n_1164),
.A2(n_1149),
.B(n_1145),
.C(n_1136),
.Y(n_1178)
);

O2A1O1Ixp33_ASAP7_75t_SL g1179 ( 
.A1(n_1162),
.A2(n_958),
.B(n_1070),
.C(n_1024),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1166),
.A2(n_1070),
.B1(n_1041),
.B2(n_1149),
.Y(n_1180)
);

OAI21xp33_ASAP7_75t_SL g1181 ( 
.A1(n_1167),
.A2(n_1097),
.B(n_1084),
.Y(n_1181)
);

INVxp67_ASAP7_75t_L g1182 ( 
.A(n_1164),
.Y(n_1182)
);

NAND4xp75_ASAP7_75t_L g1183 ( 
.A(n_1181),
.B(n_1012),
.C(n_1070),
.D(n_1002),
.Y(n_1183)
);

INVx1_ASAP7_75t_SL g1184 ( 
.A(n_1173),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1178),
.A2(n_958),
.B(n_989),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1182),
.Y(n_1186)
);

NAND4xp25_ASAP7_75t_L g1187 ( 
.A(n_1171),
.B(n_998),
.C(n_1066),
.D(n_1011),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1174),
.Y(n_1188)
);

NOR3xp33_ASAP7_75t_L g1189 ( 
.A(n_1179),
.B(n_987),
.C(n_1009),
.Y(n_1189)
);

NAND3xp33_ASAP7_75t_SL g1190 ( 
.A(n_1175),
.B(n_960),
.C(n_1070),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1186),
.Y(n_1191)
);

NOR4xp75_ASAP7_75t_L g1192 ( 
.A(n_1183),
.B(n_1172),
.C(n_1012),
.D(n_937),
.Y(n_1192)
);

AOI211xp5_ASAP7_75t_L g1193 ( 
.A1(n_1188),
.A2(n_1176),
.B(n_1180),
.C(n_1012),
.Y(n_1193)
);

NOR3xp33_ASAP7_75t_L g1194 ( 
.A(n_1187),
.B(n_986),
.C(n_994),
.Y(n_1194)
);

NAND4xp75_ASAP7_75t_L g1195 ( 
.A(n_1185),
.B(n_1012),
.C(n_1023),
.D(n_937),
.Y(n_1195)
);

NOR2x1_ASAP7_75t_L g1196 ( 
.A(n_1185),
.B(n_973),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1184),
.Y(n_1197)
);

NOR3xp33_ASAP7_75t_SL g1198 ( 
.A(n_1190),
.B(n_1023),
.C(n_1010),
.Y(n_1198)
);

NAND4xp75_ASAP7_75t_L g1199 ( 
.A(n_1196),
.B(n_1010),
.C(n_1003),
.D(n_1189),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1191),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1197),
.Y(n_1201)
);

NOR3xp33_ASAP7_75t_SL g1202 ( 
.A(n_1195),
.B(n_1070),
.C(n_977),
.Y(n_1202)
);

OR2x2_ASAP7_75t_L g1203 ( 
.A(n_1197),
.B(n_1177),
.Y(n_1203)
);

INVxp67_ASAP7_75t_L g1204 ( 
.A(n_1194),
.Y(n_1204)
);

NOR2x1_ASAP7_75t_L g1205 ( 
.A(n_1198),
.B(n_977),
.Y(n_1205)
);

AND3x2_ASAP7_75t_L g1206 ( 
.A(n_1201),
.B(n_1193),
.C(n_1192),
.Y(n_1206)
);

OR2x6_ASAP7_75t_L g1207 ( 
.A(n_1204),
.B(n_977),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_1199),
.Y(n_1208)
);

XOR2x2_ASAP7_75t_L g1209 ( 
.A(n_1205),
.B(n_960),
.Y(n_1209)
);

BUFx12f_ASAP7_75t_L g1210 ( 
.A(n_1207),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1206),
.B(n_1200),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_1211),
.B(n_1208),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1212),
.A2(n_1203),
.B1(n_1210),
.B2(n_1207),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1213),
.A2(n_1209),
.B1(n_1202),
.B2(n_978),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1214),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1215),
.B(n_978),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1216),
.A2(n_978),
.B1(n_1040),
.B2(n_1058),
.Y(n_1217)
);


endmodule