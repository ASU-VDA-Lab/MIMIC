module fake_jpeg_29716_n_316 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_316);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_316;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_11),
.B(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_0),
.B(n_2),
.Y(n_46)
);

OR2x4_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_41),
.Y(n_64)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_28),
.B1(n_39),
.B2(n_34),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_53),
.A2(n_39),
.B1(n_25),
.B2(n_36),
.Y(n_68)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_18),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_33),
.Y(n_82)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

FAx1_ASAP7_75t_SL g138 ( 
.A(n_64),
.B(n_67),
.CI(n_13),
.CON(n_138),
.SN(n_138)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_31),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_65),
.B(n_68),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_SL g66 ( 
.A(n_51),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_66),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_26),
.B(n_32),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_25),
.B1(n_20),
.B2(n_23),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_75),
.A2(n_78),
.B1(n_5),
.B2(n_8),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_77),
.B(n_80),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_54),
.A2(n_20),
.B1(n_26),
.B2(n_32),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_19),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_51),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_81),
.B(n_82),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_24),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_104),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_24),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_85),
.B(n_87),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_42),
.A2(n_40),
.B1(n_33),
.B2(n_38),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_86),
.A2(n_88),
.B1(n_94),
.B2(n_101),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_49),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_47),
.A2(n_40),
.B1(n_32),
.B2(n_26),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_41),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_92),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_62),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_44),
.A2(n_40),
.B1(n_38),
.B2(n_29),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_29),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_97),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_30),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_30),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_100),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_61),
.A2(n_32),
.B1(n_2),
.B2(n_3),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_48),
.B(n_0),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_0),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_3),
.Y(n_118)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_109),
.Y(n_157)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_110),
.Y(n_161)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_67),
.A2(n_65),
.B(n_84),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_93),
.B(n_91),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_113),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_104),
.A2(n_61),
.B1(n_57),
.B2(n_6),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_116),
.A2(n_119),
.B1(n_124),
.B2(n_131),
.Y(n_156)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_120),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_129),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_64),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

NAND2xp33_ASAP7_75t_SL g122 ( 
.A(n_74),
.B(n_83),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_138),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_65),
.B(n_5),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_128),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_63),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_126),
.A2(n_134),
.B1(n_137),
.B2(n_76),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_9),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_132),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_68),
.A2(n_100),
.B1(n_99),
.B2(n_89),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_88),
.B(n_10),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_135),
.C(n_72),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_79),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_12),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_79),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_91),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_151),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_142),
.A2(n_173),
.B(n_127),
.Y(n_181)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_147),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_138),
.B(n_15),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_148),
.B(n_152),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_106),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_150),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_123),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_70),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_125),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_138),
.B(n_16),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_154),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_70),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_155),
.B(n_159),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_102),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_73),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_162),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_73),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_114),
.B(n_16),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_166),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_112),
.A2(n_72),
.B(n_98),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_111),
.B(n_120),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_114),
.B(n_76),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_98),
.C(n_99),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_169),
.C(n_172),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_102),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_171),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_119),
.B(n_76),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_133),
.A2(n_127),
.B(n_140),
.C(n_118),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_178),
.Y(n_228)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_180),
.B(n_187),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_155),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_141),
.A2(n_127),
.B1(n_131),
.B2(n_107),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_184),
.A2(n_188),
.B1(n_192),
.B2(n_196),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_156),
.A2(n_159),
.B1(n_150),
.B2(n_172),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_186),
.A2(n_173),
.B1(n_146),
.B2(n_163),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_145),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_170),
.A2(n_107),
.B1(n_116),
.B2(n_122),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_189),
.B(n_190),
.Y(n_205)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_117),
.B1(n_109),
.B2(n_110),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_193),
.A2(n_199),
.B(n_167),
.Y(n_209)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_197),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_170),
.A2(n_132),
.B1(n_129),
.B2(n_130),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_165),
.A2(n_142),
.B(n_170),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_201),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_146),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_203),
.Y(n_217)
);

AO22x1_ASAP7_75t_L g203 ( 
.A1(n_156),
.A2(n_108),
.B1(n_173),
.B2(n_151),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_147),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_158),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_209),
.A2(n_212),
.B(n_218),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_156),
.B1(n_171),
.B2(n_169),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_210),
.A2(n_214),
.B1(n_220),
.B2(n_176),
.Y(n_247)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_155),
.B(n_154),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_203),
.A2(n_167),
.B1(n_152),
.B2(n_143),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_183),
.B(n_143),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_215),
.B(n_222),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_186),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_219),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_144),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_203),
.A2(n_145),
.B1(n_162),
.B2(n_160),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_149),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_221),
.B(n_185),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_182),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_175),
.B(n_144),
.Y(n_224)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_224),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_225),
.A2(n_226),
.B1(n_180),
.B2(n_177),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_201),
.A2(n_148),
.B1(n_153),
.B2(n_145),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_164),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_198),
.C(n_175),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_229),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_223),
.Y(n_233)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_233),
.Y(n_260)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_234),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_214),
.Y(n_253)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_236),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_181),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_247),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_220),
.A2(n_176),
.B1(n_210),
.B2(n_229),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_238),
.A2(n_217),
.B(n_209),
.Y(n_256)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_206),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_240),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_192),
.C(n_202),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_213),
.C(n_219),
.Y(n_262)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_223),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_249),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_245),
.A2(n_213),
.B1(n_222),
.B2(n_215),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_207),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_246),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_208),
.B(n_196),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_248),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_217),
.Y(n_249)
);

MAJx2_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_224),
.C(n_217),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_252),
.B(n_242),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_262),
.C(n_244),
.Y(n_273)
);

A2O1A1Ixp33_ASAP7_75t_SL g268 ( 
.A1(n_256),
.A2(n_259),
.B(n_264),
.C(n_248),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_248),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_238),
.A2(n_216),
.B(n_212),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_225),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_244),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_250),
.A2(n_226),
.B(n_188),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_241),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_269),
.Y(n_284)
);

NOR2xp67_ASAP7_75t_SL g291 ( 
.A(n_268),
.B(n_280),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_254),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_247),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_270),
.A2(n_250),
.B(n_242),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_234),
.Y(n_271)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_271),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_273),
.C(n_275),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_274),
.A2(n_257),
.B1(n_255),
.B2(n_266),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_231),
.C(n_239),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_236),
.Y(n_276)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_276),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_231),
.C(n_232),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_278),
.C(n_251),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_232),
.Y(n_278)
);

XOR2x2_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_230),
.Y(n_279)
);

OAI21x1_ASAP7_75t_L g281 ( 
.A1(n_279),
.A2(n_264),
.B(n_256),
.Y(n_281)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_287),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_195),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_255),
.C(n_258),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_258),
.C(n_263),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_290),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_289),
.B(n_287),
.Y(n_292)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_292),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_276),
.B(n_271),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_295),
.A2(n_286),
.B1(n_285),
.B2(n_190),
.Y(n_303)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_283),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_297),
.A2(n_299),
.B(n_285),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_288),
.A2(n_250),
.B1(n_268),
.B2(n_260),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_298),
.A2(n_268),
.B1(n_228),
.B2(n_243),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_300),
.B(n_293),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_303),
.Y(n_306)
);

NOR2x1_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_189),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_305),
.Y(n_308)
);

OAI31xp33_ASAP7_75t_SL g305 ( 
.A1(n_292),
.A2(n_191),
.A3(n_178),
.B(n_204),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_307),
.B(n_309),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_294),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_306),
.A2(n_301),
.B(n_305),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_310),
.B(n_312),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_308),
.B(n_191),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_158),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_158),
.C(n_108),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_313),
.Y(n_316)
);


endmodule