module real_jpeg_28752_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_312, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_312;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_0),
.A2(n_55),
.B1(n_56),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_0),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_0),
.A2(n_65),
.B1(n_67),
.B2(n_71),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_0),
.A2(n_35),
.B1(n_36),
.B2(n_71),
.Y(n_111)
);

INVx11_ASAP7_75t_SL g66 ( 
.A(n_1),
.Y(n_66)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_2),
.Y(n_95)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_5),
.Y(n_156)
);

AOI21xp33_ASAP7_75t_SL g162 ( 
.A1(n_5),
.A2(n_32),
.B(n_36),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_5),
.B(n_34),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_5),
.A2(n_55),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_5),
.B(n_55),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_5),
.B(n_60),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_5),
.A2(n_92),
.B1(n_96),
.B2(n_239),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_5),
.A2(n_35),
.B(n_254),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_6),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_6),
.A2(n_35),
.B1(n_36),
.B2(n_159),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_6),
.A2(n_55),
.B1(n_56),
.B2(n_159),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_6),
.A2(n_65),
.B1(n_67),
.B2(n_159),
.Y(n_239)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_8),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_135),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_8),
.A2(n_65),
.B1(n_67),
.B2(n_135),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_8),
.A2(n_55),
.B1(n_56),
.B2(n_135),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_L g146 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_9),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_147),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_9),
.A2(n_55),
.B1(n_56),
.B2(n_147),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_9),
.A2(n_65),
.B1(n_67),
.B2(n_147),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_10),
.A2(n_46),
.B1(n_55),
.B2(n_56),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_46),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_10),
.A2(n_46),
.B1(n_65),
.B2(n_67),
.Y(n_166)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_12),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_12),
.A2(n_55),
.B1(n_56),
.B2(n_102),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_102),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_12),
.A2(n_65),
.B1(n_67),
.B2(n_102),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_13),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_13),
.A2(n_55),
.B1(n_56),
.B2(n_59),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_13),
.A2(n_59),
.B1(n_65),
.B2(n_67),
.Y(n_128)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_15),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_16),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_16),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_L g153 ( 
.A1(n_16),
.A2(n_29),
.B1(n_55),
.B2(n_56),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_16),
.A2(n_29),
.B1(n_65),
.B2(n_67),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_17),
.A2(n_27),
.B1(n_28),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_17),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_17),
.A2(n_40),
.B1(n_55),
.B2(n_56),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_17),
.A2(n_40),
.B1(n_65),
.B2(n_67),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_116),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_115),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_103),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_22),
.B(n_103),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_75),
.C(n_81),
.Y(n_22)
);

FAx1_ASAP7_75t_SL g136 ( 
.A(n_23),
.B(n_75),
.CI(n_81),
.CON(n_136),
.SN(n_136)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_42),
.B2(n_74),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_24),
.A2(n_25),
.B1(n_105),
.B2(n_113),
.Y(n_104)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_25),
.B(n_43),
.C(n_73),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_39),
.B2(n_41),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_26),
.A2(n_30),
.B1(n_41),
.B2(n_100),
.Y(n_99)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

O2A1O1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_31)
);

NAND2xp33_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_32),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_28),
.A2(n_38),
.B(n_156),
.C(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_30),
.A2(n_41),
.B1(n_158),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_31),
.A2(n_34),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_31),
.A2(n_34),
.B1(n_101),
.B2(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_31),
.A2(n_34),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_31),
.A2(n_34),
.B1(n_134),
.B2(n_187),
.Y(n_201)
);

AO22x1_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_34)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_49),
.B(n_51),
.C(n_54),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_52),
.Y(n_51)
);

OAI32xp33_ASAP7_75t_L g262 ( 
.A1(n_35),
.A2(n_49),
.A3(n_56),
.B1(n_255),
.B2(n_263),
.Y(n_262)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_36),
.B(n_156),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_39),
.Y(n_107)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_61),
.B1(n_72),
.B2(n_73),
.Y(n_42)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_58),
.B2(n_60),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_45),
.A2(n_48),
.B1(n_54),
.B2(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_47),
.A2(n_58),
.B1(n_60),
.B2(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_47),
.A2(n_60),
.B1(n_78),
.B2(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_47),
.A2(n_60),
.B1(n_146),
.B2(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_47),
.A2(n_60),
.B1(n_132),
.B2(n_190),
.Y(n_202)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_48),
.A2(n_54),
.B1(n_145),
.B2(n_148),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_48),
.A2(n_54),
.B1(n_148),
.B2(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_48),
.A2(n_54),
.B1(n_171),
.B2(n_253),
.Y(n_252)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_56),
.B1(n_63),
.B2(n_64),
.Y(n_69)
);

OAI32xp33_ASAP7_75t_L g216 ( 
.A1(n_55),
.A2(n_63),
.A3(n_67),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_55),
.B(n_57),
.Y(n_263)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_61),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_61),
.A2(n_73),
.B1(n_110),
.B2(n_112),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_68),
.B(n_70),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_62),
.A2(n_68),
.B1(n_70),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_62),
.A2(n_68),
.B1(n_87),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_62),
.A2(n_68),
.B1(n_130),
.B2(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_62),
.A2(n_68),
.B1(n_212),
.B2(n_214),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_62),
.A2(n_68),
.B1(n_214),
.B2(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_62),
.B(n_156),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_62),
.A2(n_68),
.B1(n_152),
.B2(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_64),
.B(n_65),
.Y(n_218)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_65),
.B(n_244),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_75),
.A2(n_76),
.B(n_79),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_80),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_98),
.B(n_99),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_83),
.B1(n_120),
.B2(n_122),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_91),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_84),
.A2(n_85),
.B1(n_91),
.B2(n_98),
.Y(n_292)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_88),
.A2(n_90),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_88),
.A2(n_90),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_98),
.B1(n_99),
.B2(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_96),
.B(n_97),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_92),
.A2(n_96),
.B1(n_97),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_92),
.A2(n_96),
.B1(n_128),
.B2(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_92),
.A2(n_96),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_92),
.A2(n_96),
.B1(n_233),
.B2(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_92),
.A2(n_96),
.B1(n_228),
.B2(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_93),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_93),
.A2(n_94),
.B1(n_164),
.B2(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_93),
.A2(n_165),
.B1(n_232),
.B2(n_234),
.Y(n_231)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_96),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_96),
.B(n_156),
.Y(n_244)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_114),
.Y(n_103)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_109),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_110),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_137),
.B(n_308),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_136),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_118),
.B(n_136),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.C(n_124),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_119),
.B(n_123),
.Y(n_296)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_124),
.A2(n_125),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_131),
.C(n_133),
.Y(n_125)
);

FAx1_ASAP7_75t_SL g291 ( 
.A(n_126),
.B(n_131),
.CI(n_133),
.CON(n_291),
.SN(n_291)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_127),
.B(n_129),
.Y(n_197)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_136),
.Y(n_310)
);

AOI321xp33_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_289),
.A3(n_297),
.B1(n_302),
.B2(n_307),
.C(n_312),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_192),
.C(n_204),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_175),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_140),
.B(n_175),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_160),
.C(n_167),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_141),
.B(n_286),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_154),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_149),
.B2(n_150),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_150),
.C(n_154),
.Y(n_182)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_153),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_160),
.A2(n_167),
.B1(n_168),
.B2(n_287),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_160),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_163),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_166),
.Y(n_181)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.C(n_174),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_169),
.B(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_172),
.B(n_174),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_173),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_183),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_182),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_182),
.C(n_183),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_180),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_191),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_188),
.C(n_191),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AOI21xp33_ASAP7_75t_L g303 ( 
.A1(n_193),
.A2(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_194),
.B(n_195),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_203),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_197),
.B(n_198),
.C(n_203),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_199),
.B(n_201),
.C(n_202),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_283),
.B(n_288),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_269),
.B(n_282),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_248),
.B(n_268),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_229),
.B(n_247),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_219),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_209),
.B(n_219),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_215),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_210),
.A2(n_211),
.B1(n_215),
.B2(n_216),
.Y(n_235)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_213),
.Y(n_217)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_226),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_224),
.C(n_226),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_225),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_227),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_236),
.B(n_246),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_235),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_231),
.B(n_235),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_241),
.B(n_245),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_238),
.B(n_240),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_249),
.B(n_250),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_261),
.B1(n_266),
.B2(n_267),
.Y(n_250)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_256),
.B1(n_259),
.B2(n_260),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_252),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_256),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_260),
.C(n_267),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_258),
.Y(n_279)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_261),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_264),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_270),
.B(n_271),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_275),
.B2(n_276),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_278),
.C(n_280),
.Y(n_284)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_280),
.B2(n_281),
.Y(n_276)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_277),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_278),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_294),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_294),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.C(n_293),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_292),
.Y(n_301)
);

BUFx24_ASAP7_75t_SL g309 ( 
.A(n_291),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_298),
.A2(n_303),
.B(n_306),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_299),
.B(n_300),
.Y(n_306)
);


endmodule