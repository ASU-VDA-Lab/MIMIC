module fake_ariane_203_n_1748 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1748);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1748;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx2_ASAP7_75t_SL g155 ( 
.A(n_129),
.Y(n_155)
);

BUFx10_ASAP7_75t_L g156 ( 
.A(n_8),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_100),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_135),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_1),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_139),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_61),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_48),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_18),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_136),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_56),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_5),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_27),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_9),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_6),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_114),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_122),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_11),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_116),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_62),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_78),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_32),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_83),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_1),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_126),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_70),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_89),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_19),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_34),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_51),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_30),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_0),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_25),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_92),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_106),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_105),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_151),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_85),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_102),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_120),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_3),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_29),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_35),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_84),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_88),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_52),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_112),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_39),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_72),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_8),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_50),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_13),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_63),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_111),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_35),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_47),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_58),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_125),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_98),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_2),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_21),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_16),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_149),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_37),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_94),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_39),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_55),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_69),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_123),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_47),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_79),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_68),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_95),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_74),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_6),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_104),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_54),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_142),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_59),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_38),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_75),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_31),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_31),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_99),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_16),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_15),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_55),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_40),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_145),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_2),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_130),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_87),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_147),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_76),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_20),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g252 ( 
.A(n_108),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_58),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_80),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_22),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_115),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_44),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_59),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_143),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_49),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_26),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_118),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_60),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_103),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_14),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_101),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_86),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_96),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_41),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_41),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_57),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_51),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_26),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_81),
.Y(n_274)
);

BUFx10_ASAP7_75t_L g275 ( 
.A(n_131),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_50),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_17),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_54),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_15),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_18),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_137),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_20),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_67),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_24),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_66),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_64),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_144),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_82),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_10),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_93),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_141),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_4),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_4),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_146),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_124),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_5),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_14),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_32),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_77),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_45),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_117),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_128),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_138),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_148),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_38),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_65),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_33),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_11),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_204),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_161),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_173),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_228),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_165),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_174),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_263),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_216),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_174),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_290),
.Y(n_318)
);

INVxp33_ASAP7_75t_SL g319 ( 
.A(n_206),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_205),
.B(n_175),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_165),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_167),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_175),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_182),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_182),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_161),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_183),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_172),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_205),
.B(n_183),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_191),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_299),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_191),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_169),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_179),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_159),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_221),
.B(n_0),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_242),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_224),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_162),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_163),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_212),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_221),
.B(n_3),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_R g343 ( 
.A(n_227),
.B(n_154),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_225),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_277),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_167),
.B(n_7),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_171),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_166),
.Y(n_348)
);

INVxp33_ASAP7_75t_SL g349 ( 
.A(n_168),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_225),
.B(n_7),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_293),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_185),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_224),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_186),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_240),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_240),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_230),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_172),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_286),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_188),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_198),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_230),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_167),
.B(n_9),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_199),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_286),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_232),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_232),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_237),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_237),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_268),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_252),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_177),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_293),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_207),
.Y(n_374)
);

INVxp33_ASAP7_75t_L g375 ( 
.A(n_177),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_247),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_247),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_252),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_252),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_248),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_252),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_314),
.B(n_248),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_347),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_314),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_346),
.B(n_184),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_317),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_347),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_347),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_317),
.B(n_184),
.Y(n_389)
);

AND2x6_ASAP7_75t_L g390 ( 
.A(n_346),
.B(n_268),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_323),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_323),
.B(n_259),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_333),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_324),
.B(n_184),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_347),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_343),
.B(n_320),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_347),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_347),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_324),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_325),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_325),
.B(n_223),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_327),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_327),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_330),
.B(n_259),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_370),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_337),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_330),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g408 ( 
.A(n_321),
.B(n_337),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_332),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_332),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_344),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_344),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_357),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_357),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_329),
.B(n_264),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_353),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_362),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_363),
.B(n_241),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_362),
.B(n_264),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_366),
.B(n_285),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_366),
.B(n_367),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_367),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_368),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_368),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_369),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_369),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_376),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_376),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_377),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_377),
.B(n_285),
.Y(n_430)
);

BUFx8_ASAP7_75t_L g431 ( 
.A(n_373),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_380),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_380),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_370),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_342),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_363),
.Y(n_436)
);

OA21x2_ASAP7_75t_L g437 ( 
.A1(n_336),
.A2(n_303),
.B(n_250),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_370),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_322),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_350),
.Y(n_440)
);

BUFx8_ASAP7_75t_L g441 ( 
.A(n_373),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_335),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_328),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_358),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_372),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_351),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_400),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_400),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_400),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_396),
.B(n_349),
.Y(n_450)
);

BUFx4f_ASAP7_75t_L g451 ( 
.A(n_442),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_406),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_415),
.A2(n_319),
.B1(n_321),
.B2(n_265),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_408),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_408),
.B(n_310),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_400),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_400),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_405),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_405),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_400),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_400),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_400),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_400),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_415),
.A2(n_310),
.B1(n_326),
.B2(n_338),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_390),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_428),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_428),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_442),
.B(n_326),
.Y(n_468)
);

OAI22xp33_ASAP7_75t_L g469 ( 
.A1(n_408),
.A2(n_338),
.B1(n_375),
.B2(n_339),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_435),
.B(n_340),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_428),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_442),
.B(n_348),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_428),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_L g474 ( 
.A1(n_390),
.A2(n_313),
.B1(n_379),
.B2(n_378),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_428),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_442),
.B(n_352),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_390),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_406),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_428),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_428),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_428),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_435),
.B(n_354),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_428),
.Y(n_483)
);

BUFx10_ASAP7_75t_L g484 ( 
.A(n_442),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_435),
.B(n_360),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_384),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_399),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_384),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_442),
.B(n_361),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_384),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_439),
.B(n_364),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_406),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_439),
.B(n_374),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_399),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_405),
.Y(n_495)
);

CKINVDCx6p67_ASAP7_75t_R g496 ( 
.A(n_393),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_442),
.B(n_311),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_405),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_396),
.B(n_309),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_416),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_386),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_431),
.B(n_371),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_386),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_399),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_383),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_399),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_386),
.Y(n_507)
);

OAI22xp33_ASAP7_75t_L g508 ( 
.A1(n_440),
.A2(n_444),
.B1(n_445),
.B2(n_443),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_442),
.B(n_312),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_402),
.Y(n_510)
);

BUFx4f_ASAP7_75t_L g511 ( 
.A(n_442),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_391),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_391),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_402),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_421),
.B(n_401),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_402),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_402),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_403),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_434),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_443),
.B(n_315),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_403),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_439),
.B(n_209),
.Y(n_522)
);

INVx4_ASAP7_75t_L g523 ( 
.A(n_390),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_403),
.Y(n_524)
);

OAI22xp33_ASAP7_75t_L g525 ( 
.A1(n_440),
.A2(n_365),
.B1(n_359),
.B2(n_356),
.Y(n_525)
);

INVx5_ASAP7_75t_L g526 ( 
.A(n_390),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_421),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_439),
.B(n_316),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_440),
.A2(n_197),
.B1(n_246),
.B2(n_208),
.Y(n_529)
);

OAI22xp33_ASAP7_75t_SL g530 ( 
.A1(n_440),
.A2(n_279),
.B1(n_284),
.B2(n_251),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_434),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_383),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_443),
.B(n_318),
.Y(n_533)
);

NAND2xp33_ASAP7_75t_L g534 ( 
.A(n_390),
.B(n_391),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_434),
.Y(n_535)
);

BUFx10_ASAP7_75t_L g536 ( 
.A(n_390),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_403),
.Y(n_537)
);

NAND2xp33_ASAP7_75t_L g538 ( 
.A(n_390),
.B(n_241),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_407),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_383),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_444),
.A2(n_257),
.B1(n_220),
.B2(n_226),
.Y(n_541)
);

NAND3xp33_ASAP7_75t_L g542 ( 
.A(n_409),
.B(n_241),
.C(n_178),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_407),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_436),
.B(n_381),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_407),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_446),
.B(n_331),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_407),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_410),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_446),
.B(n_187),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_431),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_436),
.B(n_303),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_444),
.B(n_355),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_390),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_446),
.B(n_187),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_410),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_410),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_410),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_390),
.A2(n_279),
.B1(n_284),
.B2(n_276),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_427),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_409),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_390),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_434),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_390),
.A2(n_238),
.B1(n_308),
.B2(n_253),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_437),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_427),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_421),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_409),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_427),
.Y(n_568)
);

CKINVDCx6p67_ASAP7_75t_R g569 ( 
.A(n_393),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_427),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_446),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_438),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_431),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_416),
.Y(n_574)
);

NAND2xp33_ASAP7_75t_SL g575 ( 
.A(n_445),
.B(n_411),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_416),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_411),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_445),
.B(n_156),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_411),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_412),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_436),
.A2(n_235),
.B1(n_233),
.B2(n_239),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_438),
.Y(n_582)
);

INVx6_ASAP7_75t_L g583 ( 
.A(n_418),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_389),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_426),
.B(n_155),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_438),
.B(n_155),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_412),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_412),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_426),
.B(n_211),
.Y(n_589)
);

AO22x2_ASAP7_75t_L g590 ( 
.A1(n_385),
.A2(n_255),
.B1(n_189),
.B2(n_202),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_438),
.B(n_157),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_413),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_437),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_413),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_450),
.B(n_431),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_519),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_486),
.Y(n_597)
);

INVxp67_ASAP7_75t_SL g598 ( 
.A(n_495),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_465),
.B(n_413),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_486),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_465),
.B(n_414),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_465),
.B(n_414),
.Y(n_602)
);

NAND2xp33_ASAP7_75t_L g603 ( 
.A(n_480),
.B(n_470),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_452),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_488),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_465),
.B(n_477),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_571),
.B(n_508),
.Y(n_607)
);

NAND2xp33_ASAP7_75t_L g608 ( 
.A(n_480),
.B(n_414),
.Y(n_608)
);

AND2x6_ASAP7_75t_SL g609 ( 
.A(n_499),
.B(n_189),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_571),
.B(n_385),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_488),
.Y(n_611)
);

BUFx6f_ASAP7_75t_SL g612 ( 
.A(n_454),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_490),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_478),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_496),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_477),
.B(n_417),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_477),
.B(n_417),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_491),
.B(n_385),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_478),
.B(n_401),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_519),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_590),
.A2(n_437),
.B1(n_441),
.B2(n_431),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_492),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_493),
.B(n_385),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_482),
.A2(n_423),
.B1(n_422),
.B2(n_433),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_485),
.B(n_431),
.Y(n_625)
);

NAND3xp33_ASAP7_75t_L g626 ( 
.A(n_453),
.B(n_441),
.C(n_422),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_583),
.B(n_441),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_515),
.B(n_389),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_490),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_527),
.B(n_566),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_527),
.B(n_385),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_566),
.B(n_385),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_515),
.B(n_394),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_477),
.B(n_417),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_523),
.B(n_422),
.Y(n_635)
);

AND2x6_ASAP7_75t_SL g636 ( 
.A(n_544),
.B(n_202),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_SL g637 ( 
.A(n_502),
.B(n_550),
.Y(n_637)
);

NOR2xp67_ASAP7_75t_SL g638 ( 
.A(n_526),
.B(n_523),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_583),
.B(n_441),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_492),
.B(n_401),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_501),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_519),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_522),
.B(n_423),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_531),
.Y(n_644)
);

OR2x6_ASAP7_75t_L g645 ( 
.A(n_454),
.B(n_441),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_589),
.B(n_423),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_501),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_531),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_583),
.B(n_441),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_528),
.B(n_424),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_531),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_503),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_526),
.Y(n_653)
);

OAI22xp33_ASAP7_75t_L g654 ( 
.A1(n_453),
.A2(n_419),
.B1(n_382),
.B2(n_392),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_583),
.B(n_424),
.Y(n_655)
);

BUFx5_ASAP7_75t_L g656 ( 
.A(n_536),
.Y(n_656)
);

NOR3xp33_ASAP7_75t_L g657 ( 
.A(n_529),
.B(n_217),
.C(n_213),
.Y(n_657)
);

AND2x4_ASAP7_75t_SL g658 ( 
.A(n_573),
.B(n_334),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_536),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_455),
.B(n_394),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_535),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_584),
.B(n_424),
.Y(n_662)
);

NOR2xp67_ASAP7_75t_L g663 ( 
.A(n_455),
.B(n_382),
.Y(n_663)
);

A2O1A1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_563),
.A2(n_429),
.B(n_433),
.C(n_432),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_503),
.B(n_507),
.Y(n_665)
);

AND2x4_ASAP7_75t_SL g666 ( 
.A(n_573),
.B(n_341),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_578),
.B(n_425),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_468),
.B(n_425),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_507),
.B(n_425),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_575),
.A2(n_418),
.B1(n_437),
.B2(n_432),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_535),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_535),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_512),
.B(n_513),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_512),
.B(n_513),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_562),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_560),
.B(n_567),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_523),
.B(n_429),
.Y(n_677)
);

INVxp67_ASAP7_75t_SL g678 ( 
.A(n_495),
.Y(n_678)
);

INVxp67_ASAP7_75t_L g679 ( 
.A(n_500),
.Y(n_679)
);

AO221x1_ASAP7_75t_L g680 ( 
.A1(n_469),
.A2(n_241),
.B1(n_243),
.B2(n_251),
.C(n_255),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_560),
.B(n_429),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_563),
.A2(n_418),
.B1(n_437),
.B2(n_432),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_567),
.B(n_433),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_523),
.B(n_418),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_577),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_577),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_497),
.B(n_418),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_536),
.Y(n_688)
);

OR2x6_ASAP7_75t_L g689 ( 
.A(n_550),
.B(n_394),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_579),
.B(n_418),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_579),
.B(n_580),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_580),
.B(n_392),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_587),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_587),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_588),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_562),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_562),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_588),
.B(n_404),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_592),
.B(n_404),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_592),
.B(n_594),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_553),
.B(n_419),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_594),
.B(n_420),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_494),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_509),
.B(n_420),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_520),
.B(n_430),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_553),
.B(n_430),
.Y(n_706)
);

AND2x4_ASAP7_75t_SL g707 ( 
.A(n_464),
.B(n_345),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_533),
.B(n_437),
.Y(n_708)
);

NAND2xp33_ASAP7_75t_SL g709 ( 
.A(n_472),
.B(n_231),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_546),
.B(n_156),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_564),
.B(n_593),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_494),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_L g713 ( 
.A(n_480),
.B(n_241),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_536),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_572),
.Y(n_715)
);

OAI21xp5_ASAP7_75t_L g716 ( 
.A1(n_564),
.A2(n_387),
.B(n_395),
.Y(n_716)
);

BUFx2_ASAP7_75t_L g717 ( 
.A(n_576),
.Y(n_717)
);

NOR3xp33_ASAP7_75t_L g718 ( 
.A(n_541),
.B(n_213),
.C(n_217),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_553),
.B(n_219),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_451),
.A2(n_398),
.B(n_395),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_590),
.A2(n_244),
.B1(n_276),
.B2(n_296),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_SL g722 ( 
.A1(n_590),
.A2(n_307),
.B1(n_156),
.B2(n_275),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_582),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_516),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_574),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_451),
.A2(n_398),
.B(n_395),
.Y(n_726)
);

NAND3xp33_ASAP7_75t_L g727 ( 
.A(n_464),
.B(n_258),
.C(n_271),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_516),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_516),
.Y(n_729)
);

BUFx5_ASAP7_75t_L g730 ( 
.A(n_484),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_526),
.B(n_218),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_516),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_524),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_546),
.B(n_218),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_458),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_526),
.B(n_222),
.Y(n_736)
);

BUFx6f_ASAP7_75t_SL g737 ( 
.A(n_496),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_582),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_564),
.B(n_236),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_524),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_524),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_552),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_553),
.B(n_219),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_537),
.B(n_296),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_537),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_549),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_545),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_545),
.B(n_222),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_545),
.B(n_243),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_561),
.B(n_250),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_545),
.B(n_260),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_549),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_548),
.Y(n_753)
);

A2O1A1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_534),
.A2(n_272),
.B(n_260),
.C(n_261),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_SL g755 ( 
.A(n_525),
.B(n_275),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_548),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_548),
.B(n_261),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_564),
.B(n_269),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_474),
.B(n_156),
.Y(n_759)
);

O2A1O1Ixp5_ASAP7_75t_L g760 ( 
.A1(n_624),
.A2(n_511),
.B(n_451),
.C(n_476),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_725),
.B(n_569),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_663),
.B(n_554),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_598),
.A2(n_511),
.B(n_561),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_678),
.A2(n_511),
.B(n_561),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_705),
.B(n_554),
.Y(n_765)
);

AO21x1_ASAP7_75t_L g766 ( 
.A1(n_595),
.A2(n_593),
.B(n_489),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_705),
.B(n_590),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_715),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_595),
.A2(n_561),
.B1(n_538),
.B2(n_593),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_654),
.B(n_551),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_742),
.B(n_710),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_654),
.B(n_593),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_597),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_650),
.B(n_585),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_735),
.Y(n_775)
);

A2O1A1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_625),
.A2(n_510),
.B(n_543),
.C(n_548),
.Y(n_776)
);

AOI21x1_ASAP7_75t_L g777 ( 
.A1(n_719),
.A2(n_586),
.B(n_460),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_628),
.B(n_559),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_692),
.A2(n_558),
.B1(n_498),
.B2(n_559),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_725),
.Y(n_780)
);

BUFx12f_ASAP7_75t_L g781 ( 
.A(n_615),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_665),
.A2(n_498),
.B(n_484),
.Y(n_782)
);

OAI21x1_ASAP7_75t_L g783 ( 
.A1(n_716),
.A2(n_481),
.B(n_449),
.Y(n_783)
);

NOR2xp67_ASAP7_75t_SL g784 ( 
.A(n_717),
.B(n_526),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_628),
.B(n_633),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_673),
.A2(n_676),
.B(n_674),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_633),
.B(n_559),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_600),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_730),
.B(n_484),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_730),
.B(n_484),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_619),
.B(n_640),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_622),
.B(n_581),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_735),
.Y(n_793)
);

BUFx12f_ASAP7_75t_L g794 ( 
.A(n_604),
.Y(n_794)
);

BUFx4f_ASAP7_75t_L g795 ( 
.A(n_614),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_605),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_611),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_691),
.A2(n_460),
.B(n_457),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_700),
.A2(n_461),
.B(n_457),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_662),
.B(n_559),
.Y(n_800)
);

OAI22xp5_ASAP7_75t_L g801 ( 
.A1(n_698),
.A2(n_459),
.B1(n_458),
.B2(n_526),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_727),
.B(n_530),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_599),
.A2(n_462),
.B(n_461),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_662),
.B(n_530),
.Y(n_804)
);

INVx11_ASAP7_75t_L g805 ( 
.A(n_737),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_711),
.A2(n_473),
.B(n_462),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_599),
.A2(n_475),
.B(n_473),
.Y(n_807)
);

AO21x1_ASAP7_75t_L g808 ( 
.A1(n_625),
.A2(n_708),
.B(n_607),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_689),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_755),
.B(n_458),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_746),
.B(n_510),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_601),
.A2(n_479),
.B(n_475),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_601),
.A2(n_616),
.B(n_602),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_613),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_602),
.A2(n_483),
.B(n_479),
.Y(n_815)
);

AO21x1_ASAP7_75t_L g816 ( 
.A1(n_708),
.A2(n_483),
.B(n_510),
.Y(n_816)
);

O2A1O1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_618),
.A2(n_543),
.B(n_570),
.C(n_568),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_SL g818 ( 
.A1(n_759),
.A2(n_707),
.B1(n_626),
.B2(n_680),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_616),
.A2(n_463),
.B(n_456),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_660),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_752),
.B(n_543),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_707),
.B(n_569),
.Y(n_822)
);

BUFx12f_ASAP7_75t_L g823 ( 
.A(n_636),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_630),
.B(n_487),
.Y(n_824)
);

AOI21xp33_ASAP7_75t_L g825 ( 
.A1(n_739),
.A2(n_591),
.B(n_504),
.Y(n_825)
);

NOR3xp33_ASAP7_75t_L g826 ( 
.A(n_657),
.B(n_272),
.C(n_270),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_623),
.B(n_459),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_689),
.B(n_459),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_629),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_689),
.B(n_570),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_641),
.Y(n_831)
);

AOI21x1_ASAP7_75t_L g832 ( 
.A1(n_719),
.A2(n_504),
.B(n_487),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_L g833 ( 
.A1(n_711),
.A2(n_514),
.B(n_506),
.Y(n_833)
);

NOR2x2_ASAP7_75t_L g834 ( 
.A(n_645),
.B(n_506),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_627),
.A2(n_568),
.B1(n_565),
.B2(n_557),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_730),
.B(n_480),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_617),
.A2(n_463),
.B(n_456),
.Y(n_837)
);

O2A1O1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_664),
.A2(n_565),
.B(n_557),
.C(n_556),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_617),
.A2(n_471),
.B(n_467),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_634),
.A2(n_471),
.B(n_467),
.Y(n_840)
);

AO21x1_ASAP7_75t_L g841 ( 
.A1(n_758),
.A2(n_556),
.B(n_555),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_646),
.B(n_555),
.Y(n_842)
);

A2O1A1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_664),
.A2(n_547),
.B(n_514),
.C(n_539),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_627),
.A2(n_547),
.B1(n_517),
.B2(n_539),
.Y(n_844)
);

CKINVDCx10_ASAP7_75t_R g845 ( 
.A(n_737),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_730),
.B(n_656),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_704),
.A2(n_517),
.B(n_518),
.C(n_521),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_648),
.Y(n_848)
);

INVx4_ASAP7_75t_L g849 ( 
.A(n_645),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_704),
.B(n_518),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_653),
.Y(n_851)
);

AO21x1_ASAP7_75t_L g852 ( 
.A1(n_739),
.A2(n_521),
.B(n_262),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_647),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_631),
.B(n_447),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_740),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_635),
.A2(n_466),
.B(n_447),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_632),
.B(n_447),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_701),
.A2(n_466),
.B(n_448),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_745),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_677),
.A2(n_466),
.B(n_447),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_699),
.B(n_448),
.Y(n_861)
);

AO21x1_ASAP7_75t_L g862 ( 
.A1(n_758),
.A2(n_262),
.B(n_304),
.Y(n_862)
);

BUFx4f_ASAP7_75t_L g863 ( 
.A(n_645),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_639),
.A2(n_466),
.B1(n_448),
.B2(n_542),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_730),
.B(n_480),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_702),
.B(n_448),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_658),
.Y(n_867)
);

NAND2xp33_ASAP7_75t_L g868 ( 
.A(n_730),
.B(n_656),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_677),
.A2(n_540),
.B(n_532),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_658),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_652),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_685),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_701),
.A2(n_540),
.B(n_532),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_706),
.A2(n_540),
.B(n_532),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_612),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_706),
.A2(n_540),
.B(n_532),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_667),
.B(n_270),
.Y(n_877)
);

NOR2xp67_ASAP7_75t_L g878 ( 
.A(n_679),
.B(n_158),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_643),
.A2(n_540),
.B(n_532),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_684),
.B(n_278),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_603),
.A2(n_505),
.B(n_387),
.Y(n_881)
);

OR2x2_ASAP7_75t_L g882 ( 
.A(n_734),
.B(n_666),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_666),
.B(n_273),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_669),
.A2(n_505),
.B(n_387),
.Y(n_884)
);

OAI21xp33_ASAP7_75t_L g885 ( 
.A1(n_667),
.A2(n_282),
.B(n_289),
.Y(n_885)
);

INVx4_ASAP7_75t_L g886 ( 
.A(n_612),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_747),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_681),
.A2(n_505),
.B(n_387),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_683),
.A2(n_505),
.B(n_398),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_610),
.B(n_273),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_670),
.A2(n_398),
.B(n_395),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_656),
.B(n_505),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_L g893 ( 
.A1(n_686),
.A2(n_297),
.B1(n_298),
.B2(n_300),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_656),
.B(n_395),
.Y(n_894)
);

AOI21x1_ASAP7_75t_L g895 ( 
.A1(n_743),
.A2(n_304),
.B(n_280),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_693),
.Y(n_896)
);

O2A1O1Ixp5_ASAP7_75t_L g897 ( 
.A1(n_668),
.A2(n_398),
.B(n_395),
.C(n_280),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_609),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_606),
.A2(n_398),
.B(n_160),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_639),
.B(n_292),
.Y(n_900)
);

AOI21xp33_ASAP7_75t_L g901 ( 
.A1(n_687),
.A2(n_305),
.B(n_249),
.Y(n_901)
);

O2A1O1Ixp5_ASAP7_75t_L g902 ( 
.A1(n_668),
.A2(n_241),
.B(n_388),
.C(n_383),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_648),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_753),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_671),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_649),
.B(n_307),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_649),
.A2(n_245),
.B1(n_170),
.B2(n_176),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_694),
.B(n_307),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_671),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_695),
.B(n_307),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_655),
.B(n_164),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_690),
.A2(n_682),
.B(n_684),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_731),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_721),
.B(n_180),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_606),
.A2(n_256),
.B(n_181),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_723),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_687),
.B(n_10),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_718),
.B(n_275),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_721),
.B(n_190),
.Y(n_919)
);

NAND2xp33_ASAP7_75t_L g920 ( 
.A(n_656),
.B(n_192),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_720),
.A2(n_267),
.B(n_193),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_726),
.A2(n_274),
.B(n_194),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_703),
.A2(n_281),
.B(n_201),
.Y(n_923)
);

INVx4_ASAP7_75t_L g924 ( 
.A(n_731),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_738),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_736),
.B(n_195),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_712),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_724),
.A2(n_287),
.B(n_210),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_736),
.B(n_196),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_656),
.B(n_383),
.Y(n_930)
);

INVx1_ASAP7_75t_SL g931 ( 
.A(n_748),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_596),
.B(n_200),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_728),
.A2(n_283),
.B(n_203),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_744),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_729),
.B(n_12),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_732),
.A2(n_288),
.B(n_214),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_733),
.B(n_12),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_768),
.Y(n_938)
);

AND2x2_ASAP7_75t_SL g939 ( 
.A(n_863),
.B(n_621),
.Y(n_939)
);

CKINVDCx16_ASAP7_75t_R g940 ( 
.A(n_781),
.Y(n_940)
);

INVx4_ASAP7_75t_L g941 ( 
.A(n_805),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_771),
.A2(n_917),
.B1(n_792),
.B2(n_770),
.Y(n_942)
);

NAND2x1p5_ASAP7_75t_L g943 ( 
.A(n_924),
.B(n_620),
.Y(n_943)
);

BUFx2_ASAP7_75t_L g944 ( 
.A(n_780),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_SL g945 ( 
.A1(n_898),
.A2(n_722),
.B1(n_621),
.B2(n_637),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_765),
.B(n_749),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_897),
.A2(n_741),
.B(n_756),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_771),
.B(n_642),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_791),
.B(n_751),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_R g950 ( 
.A(n_845),
.B(n_709),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_912),
.B(n_644),
.Y(n_951)
);

AO21x2_ASAP7_75t_L g952 ( 
.A1(n_841),
.A2(n_750),
.B(n_743),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_775),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_868),
.A2(n_608),
.B(n_750),
.Y(n_954)
);

BUFx12f_ASAP7_75t_L g955 ( 
.A(n_794),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_785),
.B(n_651),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_772),
.B(n_661),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_917),
.A2(n_802),
.B(n_826),
.C(n_792),
.Y(n_958)
);

AO21x1_ASAP7_75t_L g959 ( 
.A1(n_786),
.A2(n_757),
.B(n_675),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_774),
.A2(n_688),
.B1(n_714),
.B2(n_659),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_842),
.A2(n_688),
.B(n_714),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_761),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_SL g963 ( 
.A1(n_935),
.A2(n_713),
.B(n_697),
.C(n_696),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_800),
.A2(n_714),
.B1(n_688),
.B2(n_659),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_802),
.A2(n_754),
.B(n_672),
.C(n_638),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_820),
.B(n_754),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_820),
.A2(n_714),
.B1(n_688),
.B2(n_659),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_826),
.A2(n_767),
.B1(n_804),
.B2(n_818),
.Y(n_968)
);

INVx4_ASAP7_75t_L g969 ( 
.A(n_828),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_775),
.Y(n_970)
);

BUFx8_ASAP7_75t_SL g971 ( 
.A(n_795),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_846),
.A2(n_659),
.B(n_653),
.Y(n_972)
);

NOR3xp33_ASAP7_75t_SL g973 ( 
.A(n_935),
.B(n_215),
.C(n_229),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_808),
.B(n_766),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_931),
.B(n_13),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_846),
.A2(n_397),
.B(n_388),
.Y(n_976)
);

AOI221xp5_ASAP7_75t_L g977 ( 
.A1(n_885),
.A2(n_291),
.B1(n_234),
.B2(n_302),
.C(n_266),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_916),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_773),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_882),
.B(n_17),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_762),
.B(n_19),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_788),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_925),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_796),
.Y(n_984)
);

BUFx8_ASAP7_75t_SL g985 ( 
.A(n_795),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_880),
.B(n_21),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_L g987 ( 
.A1(n_818),
.A2(n_275),
.B1(n_171),
.B2(n_254),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_927),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_SL g989 ( 
.A1(n_823),
.A2(n_294),
.B1(n_295),
.B2(n_301),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_848),
.B(n_254),
.Y(n_990)
);

HB1xp67_ASAP7_75t_L g991 ( 
.A(n_830),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_797),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_877),
.A2(n_22),
.B(n_23),
.C(n_25),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_913),
.B(n_23),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_SL g995 ( 
.A(n_863),
.B(n_306),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_901),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_R g997 ( 
.A(n_867),
.B(n_90),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_775),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_880),
.A2(n_28),
.B(n_30),
.C(n_33),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_814),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_822),
.B(n_34),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_829),
.B(n_36),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_831),
.B(n_36),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_867),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_903),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_900),
.A2(n_37),
.B(n_40),
.C(n_42),
.Y(n_1006)
);

INVxp67_ASAP7_75t_L g1007 ( 
.A(n_903),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_827),
.A2(n_388),
.B(n_383),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_870),
.B(n_42),
.Y(n_1009)
);

INVx3_ASAP7_75t_SL g1010 ( 
.A(n_886),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_937),
.A2(n_254),
.B(n_171),
.C(n_383),
.Y(n_1011)
);

INVxp67_ASAP7_75t_L g1012 ( 
.A(n_830),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_853),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_775),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_827),
.A2(n_397),
.B(n_388),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_855),
.Y(n_1016)
);

INVx2_ASAP7_75t_SL g1017 ( 
.A(n_870),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_871),
.B(n_43),
.Y(n_1018)
);

NAND3xp33_ASAP7_75t_SL g1019 ( 
.A(n_907),
.B(n_43),
.C(n_44),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_872),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_809),
.B(n_45),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_859),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_763),
.A2(n_388),
.B(n_383),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_896),
.B(n_46),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_810),
.B(n_46),
.Y(n_1025)
);

CKINVDCx20_ASAP7_75t_R g1026 ( 
.A(n_886),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_778),
.A2(n_171),
.B1(n_254),
.B2(n_52),
.Y(n_1027)
);

OR2x6_ASAP7_75t_L g1028 ( 
.A(n_828),
.B(n_254),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_809),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_764),
.A2(n_388),
.B(n_383),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_883),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_787),
.A2(n_254),
.B1(n_171),
.B2(n_53),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_810),
.B(n_48),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_890),
.A2(n_49),
.B(n_53),
.C(n_56),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_918),
.B(n_57),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_887),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_930),
.A2(n_397),
.B(n_388),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_883),
.Y(n_1038)
);

AOI21x1_ASAP7_75t_L g1039 ( 
.A1(n_852),
.A2(n_862),
.B(n_816),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_SL g1040 ( 
.A1(n_875),
.A2(n_171),
.B1(n_397),
.B2(n_388),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_924),
.A2(n_397),
.B1(n_388),
.B2(n_91),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_906),
.B(n_397),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_811),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_850),
.B(n_821),
.Y(n_1044)
);

OAI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_908),
.A2(n_910),
.B1(n_914),
.B2(n_919),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_861),
.A2(n_397),
.B1(n_73),
.B2(n_97),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_866),
.A2(n_397),
.B1(n_107),
.B2(n_109),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_848),
.B(n_397),
.Y(n_1048)
);

OR2x6_ASAP7_75t_L g1049 ( 
.A(n_849),
.B(n_71),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_875),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_783),
.A2(n_110),
.B(n_113),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_904),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_813),
.A2(n_119),
.B(n_121),
.C(n_127),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_930),
.A2(n_133),
.B(n_134),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_848),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_793),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_937),
.A2(n_140),
.B(n_150),
.C(n_153),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_793),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_934),
.B(n_878),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_848),
.Y(n_1060)
);

INVx4_ASAP7_75t_L g1061 ( 
.A(n_793),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_793),
.Y(n_1062)
);

OR2x6_ASAP7_75t_L g1063 ( 
.A(n_849),
.B(n_905),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_776),
.A2(n_760),
.B(n_838),
.C(n_897),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_824),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_911),
.A2(n_769),
.B1(n_776),
.B2(n_806),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_905),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_SL g1068 ( 
.A(n_784),
.B(n_933),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_905),
.B(n_909),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_834),
.Y(n_1070)
);

OR2x6_ASAP7_75t_L g1071 ( 
.A(n_905),
.B(n_909),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_909),
.B(n_929),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_779),
.A2(n_857),
.B1(n_854),
.B2(n_864),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_920),
.A2(n_892),
.B(n_790),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_932),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_926),
.B(n_893),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_909),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_1051),
.A2(n_832),
.B(n_881),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_942),
.B(n_936),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_958),
.B(n_948),
.Y(n_1080)
);

INVx5_ASAP7_75t_L g1081 ( 
.A(n_971),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_SL g1082 ( 
.A1(n_986),
.A2(n_966),
.B(n_1025),
.Y(n_1082)
);

AOI221x1_ASAP7_75t_L g1083 ( 
.A1(n_958),
.A2(n_1019),
.B1(n_1033),
.B2(n_945),
.C(n_1011),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_968),
.A2(n_835),
.B1(n_844),
.B2(n_843),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1066),
.A2(n_789),
.B(n_790),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1073),
.A2(n_789),
.B(n_892),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_948),
.B(n_915),
.Y(n_1087)
);

O2A1O1Ixp33_ASAP7_75t_SL g1088 ( 
.A1(n_1076),
.A2(n_865),
.B(n_836),
.C(n_894),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1064),
.A2(n_847),
.B(n_843),
.Y(n_1089)
);

AO32x2_ASAP7_75t_L g1090 ( 
.A1(n_1027),
.A2(n_801),
.A3(n_834),
.B1(n_847),
.B2(n_902),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1064),
.A2(n_760),
.B(n_817),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_1023),
.A2(n_777),
.B(n_884),
.Y(n_1092)
);

NAND3x1_ASAP7_75t_L g1093 ( 
.A(n_1035),
.B(n_891),
.C(n_923),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_946),
.A2(n_954),
.B(n_1074),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_979),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1042),
.A2(n_865),
.B(n_836),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1042),
.A2(n_782),
.B(n_879),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_982),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_951),
.A2(n_833),
.B(n_825),
.Y(n_1099)
);

CKINVDCx11_ASAP7_75t_R g1100 ( 
.A(n_955),
.Y(n_1100)
);

BUFx10_ASAP7_75t_L g1101 ( 
.A(n_994),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1007),
.B(n_928),
.Y(n_1102)
);

AO31x2_ASAP7_75t_L g1103 ( 
.A1(n_959),
.A2(n_876),
.A3(n_874),
.B(n_873),
.Y(n_1103)
);

AO32x2_ASAP7_75t_L g1104 ( 
.A1(n_1032),
.A2(n_902),
.A3(n_895),
.B1(n_888),
.B2(n_799),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_973),
.A2(n_899),
.B(n_922),
.C(n_921),
.Y(n_1105)
);

AOI221xp5_ASAP7_75t_SL g1106 ( 
.A1(n_999),
.A2(n_798),
.B1(n_889),
.B2(n_858),
.C(n_812),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_SL g1107 ( 
.A1(n_1057),
.A2(n_894),
.B(n_869),
.C(n_860),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_944),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_938),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_962),
.B(n_851),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1031),
.B(n_851),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_985),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_SL g1113 ( 
.A(n_939),
.B(n_856),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_973),
.A2(n_803),
.B(n_807),
.C(n_815),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_941),
.Y(n_1115)
);

AOI221xp5_ASAP7_75t_SL g1116 ( 
.A1(n_993),
.A2(n_819),
.B1(n_837),
.B2(n_839),
.C(n_840),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_984),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_969),
.B(n_994),
.Y(n_1118)
);

NAND3xp33_ASAP7_75t_L g1119 ( 
.A(n_996),
.B(n_1006),
.C(n_1034),
.Y(n_1119)
);

AO31x2_ASAP7_75t_L g1120 ( 
.A1(n_1011),
.A2(n_965),
.A3(n_1072),
.B(n_961),
.Y(n_1120)
);

CKINVDCx20_ASAP7_75t_R g1121 ( 
.A(n_940),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1065),
.B(n_1044),
.Y(n_1122)
);

AO31x2_ASAP7_75t_L g1123 ( 
.A1(n_965),
.A2(n_1072),
.A3(n_1046),
.B(n_1047),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_992),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_968),
.A2(n_987),
.B(n_1075),
.C(n_981),
.Y(n_1125)
);

OAI22x1_ASAP7_75t_L g1126 ( 
.A1(n_1070),
.A2(n_1021),
.B1(n_1029),
.B2(n_1001),
.Y(n_1126)
);

AOI21xp33_ASAP7_75t_L g1127 ( 
.A1(n_987),
.A2(n_1045),
.B(n_939),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_951),
.A2(n_1068),
.B(n_1015),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1000),
.Y(n_1129)
);

OR2x2_ASAP7_75t_L g1130 ( 
.A(n_1038),
.B(n_1005),
.Y(n_1130)
);

BUFx12f_ASAP7_75t_L g1131 ( 
.A(n_941),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1008),
.A2(n_963),
.B(n_964),
.Y(n_1132)
);

AO22x2_ASAP7_75t_L g1133 ( 
.A1(n_974),
.A2(n_1019),
.B1(n_957),
.B2(n_1059),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_957),
.A2(n_974),
.B(n_947),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_998),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1007),
.B(n_949),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1039),
.A2(n_976),
.B(n_1037),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_963),
.A2(n_960),
.B(n_972),
.Y(n_1138)
);

OAI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_980),
.A2(n_975),
.B1(n_1009),
.B2(n_995),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_967),
.A2(n_1048),
.B(n_1045),
.Y(n_1140)
);

AO31x2_ASAP7_75t_L g1141 ( 
.A1(n_1055),
.A2(n_1067),
.A3(n_1060),
.B(n_1053),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1048),
.A2(n_1054),
.B(n_1069),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_969),
.B(n_1012),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_978),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1021),
.B(n_1050),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1043),
.B(n_1012),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1069),
.A2(n_990),
.B(n_1071),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_950),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_991),
.B(n_1013),
.Y(n_1149)
);

AOI21x1_ASAP7_75t_L g1150 ( 
.A1(n_990),
.A2(n_1077),
.B(n_1071),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_956),
.B(n_1020),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_956),
.B(n_1062),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_983),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_991),
.B(n_1017),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1016),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1002),
.A2(n_1024),
.B(n_1018),
.C(n_1003),
.Y(n_1156)
);

AO21x1_ASAP7_75t_L g1157 ( 
.A1(n_1041),
.A2(n_943),
.B(n_1061),
.Y(n_1157)
);

AOI21x1_ASAP7_75t_SL g1158 ( 
.A1(n_1010),
.A2(n_950),
.B(n_997),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1022),
.B(n_1036),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_1010),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1028),
.A2(n_1049),
.B1(n_1040),
.B2(n_943),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1052),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1058),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_998),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_953),
.A2(n_970),
.B(n_1014),
.Y(n_1165)
);

BUFx12f_ASAP7_75t_L g1166 ( 
.A(n_1028),
.Y(n_1166)
);

AO31x2_ASAP7_75t_L g1167 ( 
.A1(n_952),
.A2(n_1061),
.A3(n_1071),
.B(n_1063),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_953),
.A2(n_1014),
.B(n_970),
.Y(n_1168)
);

OA21x2_ASAP7_75t_L g1169 ( 
.A1(n_952),
.A2(n_977),
.B(n_1063),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_1063),
.B(n_1004),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1028),
.A2(n_1049),
.B(n_998),
.Y(n_1171)
);

AOI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1049),
.A2(n_998),
.B(n_1056),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1056),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1026),
.A2(n_1056),
.B(n_1062),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1056),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1062),
.A2(n_989),
.B(n_997),
.Y(n_1176)
);

O2A1O1Ixp5_ASAP7_75t_L g1177 ( 
.A1(n_1062),
.A2(n_958),
.B(n_595),
.C(n_986),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1051),
.A2(n_1030),
.B(n_1023),
.Y(n_1178)
);

AOI221x1_ASAP7_75t_L g1179 ( 
.A1(n_958),
.A2(n_1019),
.B1(n_986),
.B2(n_595),
.C(n_1025),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_958),
.A2(n_511),
.B(n_451),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_958),
.A2(n_511),
.B(n_451),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_979),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_958),
.A2(n_511),
.B(n_451),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_944),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1051),
.A2(n_1030),
.B(n_1023),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_944),
.Y(n_1186)
);

NOR4xp25_ASAP7_75t_L g1187 ( 
.A(n_958),
.B(n_999),
.C(n_1019),
.D(n_996),
.Y(n_1187)
);

AOI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1039),
.A2(n_974),
.B(n_852),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_958),
.A2(n_511),
.B(n_451),
.Y(n_1189)
);

AOI221xp5_ASAP7_75t_L g1190 ( 
.A1(n_958),
.A2(n_654),
.B1(n_453),
.B2(n_942),
.C(n_469),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_942),
.A2(n_958),
.B1(n_595),
.B2(n_576),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_958),
.A2(n_942),
.B(n_770),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1051),
.A2(n_1030),
.B(n_1023),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_942),
.B(n_454),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_944),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_958),
.A2(n_511),
.B(n_451),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_969),
.B(n_828),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_958),
.A2(n_942),
.B(n_625),
.C(n_595),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_979),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_944),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_SL g1201 ( 
.A1(n_958),
.A2(n_942),
.B(n_770),
.C(n_986),
.Y(n_1201)
);

NAND3x1_ASAP7_75t_L g1202 ( 
.A(n_942),
.B(n_453),
.C(n_1035),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_958),
.A2(n_511),
.B(n_451),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_958),
.A2(n_511),
.B(n_451),
.Y(n_1204)
);

INVx1_ASAP7_75t_SL g1205 ( 
.A(n_944),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1051),
.A2(n_1030),
.B(n_1023),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1051),
.A2(n_1030),
.B(n_1023),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_942),
.A2(n_958),
.B1(n_770),
.B2(n_917),
.Y(n_1208)
);

INVx3_ASAP7_75t_SL g1209 ( 
.A(n_940),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_958),
.A2(n_511),
.B(n_451),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_979),
.Y(n_1211)
);

OR2x6_ASAP7_75t_L g1212 ( 
.A(n_1028),
.B(n_645),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_958),
.A2(n_511),
.B(n_451),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_958),
.A2(n_450),
.B(n_396),
.C(n_986),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_988),
.Y(n_1215)
);

AO32x2_ASAP7_75t_L g1216 ( 
.A1(n_945),
.A2(n_1066),
.A3(n_1073),
.B1(n_1032),
.B2(n_1027),
.Y(n_1216)
);

CKINVDCx6p67_ASAP7_75t_R g1217 ( 
.A(n_1081),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1122),
.B(n_1136),
.Y(n_1218)
);

BUFx8_ASAP7_75t_SL g1219 ( 
.A(n_1121),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_1197),
.Y(n_1220)
);

BUFx8_ASAP7_75t_L g1221 ( 
.A(n_1112),
.Y(n_1221)
);

BUFx4f_ASAP7_75t_L g1222 ( 
.A(n_1131),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_SL g1223 ( 
.A1(n_1198),
.A2(n_1208),
.B(n_1125),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1190),
.A2(n_1127),
.B1(n_1208),
.B2(n_1192),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1127),
.A2(n_1192),
.B1(n_1080),
.B2(n_1191),
.Y(n_1225)
);

CKINVDCx11_ASAP7_75t_R g1226 ( 
.A(n_1100),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1202),
.A2(n_1079),
.B1(n_1194),
.B2(n_1145),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1186),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1095),
.Y(n_1229)
);

BUFx8_ASAP7_75t_L g1230 ( 
.A(n_1115),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1098),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1117),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_1170),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_SL g1234 ( 
.A1(n_1214),
.A2(n_1179),
.B(n_1083),
.Y(n_1234)
);

CKINVDCx11_ASAP7_75t_R g1235 ( 
.A(n_1209),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1124),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1122),
.B(n_1151),
.Y(n_1237)
);

CKINVDCx6p67_ASAP7_75t_R g1238 ( 
.A(n_1101),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1151),
.B(n_1118),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1101),
.B(n_1108),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1129),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1133),
.A2(n_1084),
.B1(n_1139),
.B2(n_1119),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_1148),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_1184),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_1195),
.Y(n_1245)
);

INVx1_ASAP7_75t_SL g1246 ( 
.A(n_1108),
.Y(n_1246)
);

INVx6_ASAP7_75t_L g1247 ( 
.A(n_1197),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1133),
.A2(n_1084),
.B1(n_1119),
.B2(n_1126),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_SL g1249 ( 
.A1(n_1161),
.A2(n_1113),
.B1(n_1082),
.B2(n_1212),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_1200),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1174),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1120),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1161),
.A2(n_1212),
.B1(n_1146),
.B2(n_1170),
.Y(n_1253)
);

INVx4_ASAP7_75t_L g1254 ( 
.A(n_1143),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1188),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_SL g1256 ( 
.A1(n_1113),
.A2(n_1212),
.B1(n_1166),
.B2(n_1169),
.Y(n_1256)
);

INVx6_ASAP7_75t_L g1257 ( 
.A(n_1143),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_1160),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_SL g1259 ( 
.A(n_1177),
.B(n_1187),
.Y(n_1259)
);

INVx6_ASAP7_75t_L g1260 ( 
.A(n_1130),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1182),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1199),
.A2(n_1211),
.B1(n_1155),
.B2(n_1162),
.Y(n_1262)
);

INVx1_ASAP7_75t_SL g1263 ( 
.A(n_1200),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1149),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_SL g1265 ( 
.A1(n_1187),
.A2(n_1205),
.B1(n_1158),
.B2(n_1174),
.Y(n_1265)
);

CKINVDCx11_ASAP7_75t_R g1266 ( 
.A(n_1205),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1159),
.Y(n_1267)
);

INVxp67_ASAP7_75t_L g1268 ( 
.A(n_1154),
.Y(n_1268)
);

INVx3_ASAP7_75t_L g1269 ( 
.A(n_1172),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1159),
.Y(n_1270)
);

NAND2x1p5_ASAP7_75t_L g1271 ( 
.A(n_1110),
.B(n_1111),
.Y(n_1271)
);

AOI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1201),
.A2(n_1176),
.B1(n_1163),
.B2(n_1152),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1215),
.A2(n_1153),
.B1(n_1144),
.B2(n_1109),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1141),
.Y(n_1274)
);

INVx1_ASAP7_75t_SL g1275 ( 
.A(n_1135),
.Y(n_1275)
);

INVx6_ASAP7_75t_L g1276 ( 
.A(n_1171),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1141),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1156),
.B(n_1102),
.Y(n_1278)
);

AOI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1093),
.A2(n_1087),
.B1(n_1157),
.B2(n_1140),
.Y(n_1279)
);

BUFx10_ASAP7_75t_L g1280 ( 
.A(n_1173),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_1135),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1175),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1165),
.Y(n_1283)
);

BUFx8_ASAP7_75t_L g1284 ( 
.A(n_1216),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1168),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1089),
.A2(n_1091),
.B1(n_1134),
.B2(n_1169),
.Y(n_1286)
);

INVx1_ASAP7_75t_SL g1287 ( 
.A(n_1164),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1180),
.A2(n_1196),
.B1(n_1189),
.B2(n_1183),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_1164),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1181),
.A2(n_1203),
.B1(n_1213),
.B2(n_1210),
.Y(n_1290)
);

NAND2x1p5_ASAP7_75t_L g1291 ( 
.A(n_1150),
.B(n_1147),
.Y(n_1291)
);

BUFx12f_ASAP7_75t_L g1292 ( 
.A(n_1167),
.Y(n_1292)
);

BUFx8_ASAP7_75t_L g1293 ( 
.A(n_1216),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1134),
.A2(n_1204),
.B1(n_1099),
.B2(n_1086),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1090),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_SL g1296 ( 
.A1(n_1090),
.A2(n_1085),
.B1(n_1128),
.B2(n_1123),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1094),
.A2(n_1096),
.B1(n_1132),
.B2(n_1090),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1142),
.A2(n_1138),
.B1(n_1097),
.B2(n_1123),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1103),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_1120),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_SL g1301 ( 
.A1(n_1123),
.A2(n_1120),
.B1(n_1137),
.B2(n_1105),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1088),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1103),
.Y(n_1303)
);

OAI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1106),
.A2(n_1114),
.B1(n_1104),
.B2(n_1116),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_SL g1305 ( 
.A1(n_1178),
.A2(n_1207),
.B1(n_1206),
.B2(n_1193),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1092),
.Y(n_1306)
);

INVx4_ASAP7_75t_L g1307 ( 
.A(n_1106),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_SL g1308 ( 
.A1(n_1107),
.A2(n_1116),
.B(n_1104),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1104),
.B(n_1185),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1078),
.A2(n_1190),
.B1(n_1127),
.B2(n_1208),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1095),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1190),
.A2(n_1127),
.B1(n_1208),
.B2(n_759),
.Y(n_1312)
);

OAI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1190),
.A2(n_942),
.B1(n_1191),
.B2(n_1208),
.Y(n_1313)
);

AOI22xp5_ASAP7_75t_SL g1314 ( 
.A1(n_1121),
.A2(n_1126),
.B1(n_393),
.B2(n_169),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1131),
.Y(n_1315)
);

INVx1_ASAP7_75t_SL g1316 ( 
.A(n_1108),
.Y(n_1316)
);

BUFx8_ASAP7_75t_SL g1317 ( 
.A(n_1121),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1190),
.A2(n_1127),
.B1(n_1208),
.B2(n_759),
.Y(n_1318)
);

INVx6_ASAP7_75t_L g1319 ( 
.A(n_1131),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1190),
.A2(n_942),
.B1(n_595),
.B2(n_958),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1190),
.A2(n_1127),
.B1(n_1208),
.B2(n_759),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1190),
.A2(n_1127),
.B1(n_1208),
.B2(n_759),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1122),
.B(n_942),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1190),
.A2(n_1127),
.B1(n_1208),
.B2(n_759),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1095),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_SL g1326 ( 
.A1(n_1208),
.A2(n_945),
.B1(n_707),
.B2(n_755),
.Y(n_1326)
);

INVx4_ASAP7_75t_L g1327 ( 
.A(n_1131),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_1186),
.Y(n_1328)
);

CKINVDCx11_ASAP7_75t_R g1329 ( 
.A(n_1100),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1095),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1095),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1190),
.A2(n_1127),
.B1(n_1208),
.B2(n_759),
.Y(n_1332)
);

INVx6_ASAP7_75t_L g1333 ( 
.A(n_1131),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1131),
.Y(n_1334)
);

INVx1_ASAP7_75t_SL g1335 ( 
.A(n_1108),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1145),
.B(n_1101),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1208),
.A2(n_945),
.B1(n_707),
.B2(n_755),
.Y(n_1337)
);

INVx8_ASAP7_75t_L g1338 ( 
.A(n_1081),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1283),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1276),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1285),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1303),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1295),
.B(n_1286),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1276),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1239),
.B(n_1218),
.Y(n_1345)
);

INVx2_ASAP7_75t_SL g1346 ( 
.A(n_1280),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1266),
.B(n_1250),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1298),
.A2(n_1290),
.B(n_1288),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1295),
.B(n_1286),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1295),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1244),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1320),
.A2(n_1313),
.B1(n_1337),
.B2(n_1326),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1229),
.B(n_1231),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1252),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_1245),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1252),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1232),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1236),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1241),
.Y(n_1359)
);

OAI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1313),
.A2(n_1227),
.B1(n_1323),
.B2(n_1234),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1298),
.A2(n_1306),
.B(n_1299),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1261),
.Y(n_1362)
);

NOR2xp67_ASAP7_75t_L g1363 ( 
.A(n_1279),
.B(n_1278),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1311),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_SL g1365 ( 
.A1(n_1284),
.A2(n_1293),
.B1(n_1314),
.B2(n_1265),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1237),
.B(n_1264),
.Y(n_1366)
);

INVx2_ASAP7_75t_SL g1367 ( 
.A(n_1280),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1300),
.B(n_1233),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1325),
.Y(n_1369)
);

AO21x2_ASAP7_75t_L g1370 ( 
.A1(n_1304),
.A2(n_1274),
.B(n_1277),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1233),
.B(n_1269),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1330),
.Y(n_1372)
);

OR2x6_ASAP7_75t_L g1373 ( 
.A(n_1223),
.B(n_1291),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1331),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1219),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1267),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1270),
.Y(n_1377)
);

INVx4_ASAP7_75t_L g1378 ( 
.A(n_1254),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1306),
.A2(n_1297),
.B(n_1294),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1297),
.A2(n_1294),
.B(n_1302),
.Y(n_1380)
);

AO21x2_ASAP7_75t_L g1381 ( 
.A1(n_1304),
.A2(n_1277),
.B(n_1255),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1268),
.Y(n_1382)
);

INVx3_ASAP7_75t_L g1383 ( 
.A(n_1307),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1291),
.A2(n_1310),
.B(n_1308),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1307),
.B(n_1248),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1246),
.B(n_1263),
.Y(n_1386)
);

INVx4_ASAP7_75t_L g1387 ( 
.A(n_1254),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1248),
.B(n_1309),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1225),
.B(n_1224),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1225),
.B(n_1224),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1282),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1269),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1276),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1281),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1262),
.Y(n_1395)
);

AO21x1_ASAP7_75t_L g1396 ( 
.A1(n_1259),
.A2(n_1242),
.B(n_1272),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1262),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1259),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1242),
.B(n_1310),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1301),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1271),
.B(n_1296),
.Y(n_1401)
);

AOI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1240),
.A2(n_1336),
.B(n_1251),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_SL g1403 ( 
.A1(n_1312),
.A2(n_1318),
.B(n_1332),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1292),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1271),
.B(n_1316),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1292),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1312),
.A2(n_1321),
.B(n_1332),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1338),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1284),
.Y(n_1409)
);

AND2x4_ASAP7_75t_SL g1410 ( 
.A(n_1253),
.B(n_1220),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1249),
.B(n_1328),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1293),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1228),
.B(n_1335),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1260),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1256),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1305),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1260),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1260),
.B(n_1318),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1351),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1382),
.B(n_1253),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1389),
.A2(n_1321),
.B1(n_1324),
.B2(n_1322),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1352),
.A2(n_1322),
.B(n_1324),
.Y(n_1422)
);

O2A1O1Ixp33_ASAP7_75t_L g1423 ( 
.A1(n_1360),
.A2(n_1258),
.B(n_1287),
.C(n_1275),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1368),
.B(n_1289),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1394),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1398),
.B(n_1238),
.Y(n_1426)
);

INVxp67_ASAP7_75t_SL g1427 ( 
.A(n_1363),
.Y(n_1427)
);

NAND2xp33_ASAP7_75t_R g1428 ( 
.A(n_1375),
.B(n_1329),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1413),
.B(n_1217),
.Y(n_1429)
);

A2O1A1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1352),
.A2(n_1222),
.B(n_1334),
.C(n_1315),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1355),
.B(n_1317),
.Y(n_1431)
);

OA21x2_ASAP7_75t_L g1432 ( 
.A1(n_1348),
.A2(n_1273),
.B(n_1257),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1405),
.B(n_1338),
.Y(n_1433)
);

AND2x4_ASAP7_75t_L g1434 ( 
.A(n_1368),
.B(n_1334),
.Y(n_1434)
);

AO32x2_ASAP7_75t_L g1435 ( 
.A1(n_1346),
.A2(n_1327),
.A3(n_1235),
.B1(n_1230),
.B2(n_1221),
.Y(n_1435)
);

O2A1O1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1390),
.A2(n_1315),
.B(n_1243),
.C(n_1230),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1398),
.B(n_1220),
.Y(n_1437)
);

AO32x2_ASAP7_75t_L g1438 ( 
.A1(n_1346),
.A2(n_1327),
.A3(n_1221),
.B1(n_1329),
.B2(n_1319),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1376),
.B(n_1247),
.Y(n_1439)
);

AOI221xp5_ASAP7_75t_L g1440 ( 
.A1(n_1399),
.A2(n_1226),
.B1(n_1319),
.B2(n_1333),
.C(n_1247),
.Y(n_1440)
);

AO22x2_ASAP7_75t_L g1441 ( 
.A1(n_1404),
.A2(n_1319),
.B1(n_1333),
.B2(n_1406),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1376),
.B(n_1377),
.Y(n_1442)
);

AOI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1399),
.A2(n_1396),
.B1(n_1365),
.B2(n_1407),
.Y(n_1443)
);

AO21x2_ASAP7_75t_L g1444 ( 
.A1(n_1416),
.A2(n_1363),
.B(n_1400),
.Y(n_1444)
);

O2A1O1Ixp33_ASAP7_75t_L g1445 ( 
.A1(n_1396),
.A2(n_1403),
.B(n_1385),
.C(n_1416),
.Y(n_1445)
);

AO32x2_ASAP7_75t_L g1446 ( 
.A1(n_1367),
.A2(n_1408),
.A3(n_1378),
.B1(n_1387),
.B2(n_1388),
.Y(n_1446)
);

AO32x2_ASAP7_75t_L g1447 ( 
.A1(n_1367),
.A2(n_1408),
.A3(n_1378),
.B1(n_1387),
.B2(n_1388),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1377),
.B(n_1345),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1366),
.B(n_1353),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1347),
.B(n_1386),
.Y(n_1450)
);

AOI221xp5_ASAP7_75t_L g1451 ( 
.A1(n_1403),
.A2(n_1385),
.B1(n_1400),
.B2(n_1395),
.C(n_1397),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1350),
.Y(n_1452)
);

NAND4xp25_ASAP7_75t_L g1453 ( 
.A(n_1383),
.B(n_1411),
.C(n_1339),
.D(n_1341),
.Y(n_1453)
);

OA21x2_ASAP7_75t_L g1454 ( 
.A1(n_1348),
.A2(n_1384),
.B(n_1379),
.Y(n_1454)
);

O2A1O1Ixp33_ASAP7_75t_SL g1455 ( 
.A1(n_1405),
.A2(n_1394),
.B(n_1357),
.C(n_1372),
.Y(n_1455)
);

AO32x2_ASAP7_75t_L g1456 ( 
.A1(n_1378),
.A2(n_1387),
.A3(n_1402),
.B1(n_1343),
.B2(n_1349),
.Y(n_1456)
);

INVx4_ASAP7_75t_L g1457 ( 
.A(n_1394),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1357),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1371),
.B(n_1394),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1358),
.B(n_1359),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1371),
.B(n_1414),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1358),
.B(n_1359),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1401),
.B(n_1349),
.Y(n_1463)
);

O2A1O1Ixp33_ASAP7_75t_L g1464 ( 
.A1(n_1373),
.A2(n_1383),
.B(n_1418),
.C(n_1393),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1409),
.B(n_1412),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1409),
.B(n_1412),
.Y(n_1466)
);

A2O1A1Ixp33_ASAP7_75t_L g1467 ( 
.A1(n_1415),
.A2(n_1397),
.B(n_1395),
.C(n_1410),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1362),
.B(n_1364),
.Y(n_1468)
);

AOI211xp5_ASAP7_75t_L g1469 ( 
.A1(n_1415),
.A2(n_1380),
.B(n_1379),
.C(n_1362),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1402),
.B(n_1417),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_SL g1471 ( 
.A(n_1378),
.B(n_1387),
.Y(n_1471)
);

AOI221xp5_ASAP7_75t_L g1472 ( 
.A1(n_1369),
.A2(n_1374),
.B1(n_1391),
.B2(n_1356),
.C(n_1354),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1448),
.B(n_1369),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1458),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1452),
.Y(n_1475)
);

OAI221xp5_ASAP7_75t_SL g1476 ( 
.A1(n_1443),
.A2(n_1391),
.B1(n_1354),
.B2(n_1356),
.C(n_1340),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1459),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1454),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1446),
.Y(n_1479)
);

INVxp67_ASAP7_75t_SL g1480 ( 
.A(n_1427),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1462),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1454),
.B(n_1341),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1446),
.B(n_1392),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1422),
.A2(n_1421),
.B1(n_1451),
.B2(n_1443),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1449),
.B(n_1381),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1456),
.B(n_1381),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1456),
.B(n_1381),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1462),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1449),
.B(n_1342),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1419),
.B(n_1370),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1456),
.B(n_1446),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1447),
.B(n_1370),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1447),
.B(n_1361),
.Y(n_1493)
);

INVxp67_ASAP7_75t_L g1494 ( 
.A(n_1470),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1442),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1442),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1447),
.B(n_1370),
.Y(n_1497)
);

NOR2x1p5_ASAP7_75t_L g1498 ( 
.A(n_1453),
.B(n_1344),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1460),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1468),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1425),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1481),
.B(n_1472),
.Y(n_1502)
);

OA21x2_ASAP7_75t_L g1503 ( 
.A1(n_1478),
.A2(n_1467),
.B(n_1453),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1501),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1489),
.B(n_1437),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1482),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1489),
.B(n_1437),
.Y(n_1507)
);

CKINVDCx16_ASAP7_75t_R g1508 ( 
.A(n_1477),
.Y(n_1508)
);

AND2x2_ASAP7_75t_SL g1509 ( 
.A(n_1491),
.B(n_1479),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1481),
.B(n_1488),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1491),
.B(n_1463),
.Y(n_1511)
);

AO21x2_ASAP7_75t_L g1512 ( 
.A1(n_1478),
.A2(n_1445),
.B(n_1444),
.Y(n_1512)
);

BUFx3_ASAP7_75t_L g1513 ( 
.A(n_1501),
.Y(n_1513)
);

OAI221xp5_ASAP7_75t_L g1514 ( 
.A1(n_1484),
.A2(n_1423),
.B1(n_1469),
.B2(n_1430),
.C(n_1420),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1474),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1491),
.B(n_1469),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1478),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1478),
.Y(n_1518)
);

AOI221xp5_ASAP7_75t_L g1519 ( 
.A1(n_1484),
.A2(n_1440),
.B1(n_1436),
.B2(n_1455),
.C(n_1450),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1479),
.B(n_1466),
.Y(n_1520)
);

NOR2xp67_ASAP7_75t_L g1521 ( 
.A(n_1492),
.B(n_1457),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1479),
.B(n_1465),
.Y(n_1522)
);

OAI322xp33_ASAP7_75t_L g1523 ( 
.A1(n_1490),
.A2(n_1426),
.A3(n_1439),
.B1(n_1428),
.B2(n_1464),
.C1(n_1433),
.C2(n_1431),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1473),
.B(n_1429),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1500),
.B(n_1439),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1474),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1483),
.B(n_1461),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1483),
.B(n_1457),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1482),
.Y(n_1529)
);

AOI21xp33_ASAP7_75t_L g1530 ( 
.A1(n_1490),
.A2(n_1426),
.B(n_1492),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1474),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1481),
.B(n_1342),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1485),
.B(n_1424),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1480),
.B(n_1434),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1483),
.B(n_1424),
.Y(n_1535)
);

NOR3xp33_ASAP7_75t_SL g1536 ( 
.A(n_1476),
.B(n_1435),
.C(n_1471),
.Y(n_1536)
);

NAND2x1p5_ASAP7_75t_L g1537 ( 
.A(n_1498),
.B(n_1432),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1482),
.Y(n_1538)
);

INVxp67_ASAP7_75t_SL g1539 ( 
.A(n_1490),
.Y(n_1539)
);

BUFx3_ASAP7_75t_L g1540 ( 
.A(n_1501),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1509),
.B(n_1480),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1510),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1509),
.B(n_1493),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1509),
.B(n_1493),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1516),
.B(n_1511),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1516),
.B(n_1493),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1516),
.B(n_1493),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1502),
.B(n_1488),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1502),
.B(n_1510),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1532),
.B(n_1495),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1515),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1511),
.B(n_1492),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_L g1553 ( 
.A(n_1524),
.B(n_1434),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1532),
.B(n_1495),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1511),
.B(n_1497),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1515),
.B(n_1495),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1526),
.B(n_1496),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1526),
.B(n_1496),
.Y(n_1558)
);

INVxp67_ASAP7_75t_L g1559 ( 
.A(n_1512),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1528),
.B(n_1497),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1528),
.B(n_1497),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1521),
.B(n_1498),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1531),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1529),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1528),
.B(n_1494),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1531),
.B(n_1496),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1506),
.B(n_1485),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1506),
.B(n_1475),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1539),
.B(n_1482),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1505),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1505),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1527),
.B(n_1498),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1529),
.B(n_1538),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1527),
.B(n_1535),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1539),
.B(n_1499),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1529),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1507),
.Y(n_1577)
);

NOR2x1_ASAP7_75t_L g1578 ( 
.A(n_1541),
.B(n_1523),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1551),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1551),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1545),
.B(n_1508),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1563),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1549),
.B(n_1520),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1563),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1549),
.B(n_1523),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1573),
.Y(n_1586)
);

AOI21xp33_ASAP7_75t_SL g1587 ( 
.A1(n_1541),
.A2(n_1508),
.B(n_1534),
.Y(n_1587)
);

OAI21xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1543),
.A2(n_1522),
.B(n_1520),
.Y(n_1588)
);

AND2x4_ASAP7_75t_SL g1589 ( 
.A(n_1562),
.B(n_1536),
.Y(n_1589)
);

AOI31xp33_ASAP7_75t_L g1590 ( 
.A1(n_1541),
.A2(n_1519),
.A3(n_1537),
.B(n_1520),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1545),
.B(n_1535),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1545),
.B(n_1536),
.Y(n_1592)
);

INVx2_ASAP7_75t_SL g1593 ( 
.A(n_1562),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1548),
.B(n_1507),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1573),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1573),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1548),
.B(n_1522),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1543),
.A2(n_1514),
.B(n_1519),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1543),
.B(n_1535),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1544),
.B(n_1574),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1570),
.B(n_1522),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1564),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1570),
.B(n_1525),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1556),
.Y(n_1604)
);

NAND4xp25_ASAP7_75t_L g1605 ( 
.A(n_1544),
.B(n_1540),
.C(n_1504),
.D(n_1513),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1571),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1571),
.B(n_1475),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1577),
.Y(n_1608)
);

INVxp33_ASAP7_75t_L g1609 ( 
.A(n_1544),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1577),
.Y(n_1610)
);

INVx1_ASAP7_75t_SL g1611 ( 
.A(n_1572),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1556),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1546),
.B(n_1525),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1550),
.B(n_1533),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1550),
.B(n_1533),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1554),
.B(n_1533),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1564),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1557),
.Y(n_1618)
);

NOR2xp67_ASAP7_75t_SL g1619 ( 
.A(n_1572),
.B(n_1514),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1585),
.B(n_1546),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1582),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1600),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1582),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1581),
.B(n_1574),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1598),
.B(n_1546),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1581),
.B(n_1600),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1594),
.B(n_1554),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1619),
.B(n_1547),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1619),
.B(n_1547),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1579),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1580),
.Y(n_1631)
);

CKINVDCx16_ASAP7_75t_R g1632 ( 
.A(n_1592),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1590),
.B(n_1553),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1594),
.B(n_1547),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1584),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1606),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_L g1637 ( 
.A(n_1592),
.B(n_1578),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1591),
.B(n_1574),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1603),
.B(n_1575),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1591),
.B(n_1552),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1599),
.B(n_1552),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1592),
.B(n_1572),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1608),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1603),
.B(n_1575),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1583),
.B(n_1568),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1610),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1607),
.B(n_1568),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1586),
.Y(n_1648)
);

NAND2xp33_ASAP7_75t_L g1649 ( 
.A(n_1593),
.B(n_1568),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1614),
.B(n_1567),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1602),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1589),
.B(n_1562),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1597),
.B(n_1542),
.Y(n_1653)
);

OR2x6_ASAP7_75t_L g1654 ( 
.A(n_1593),
.B(n_1441),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1637),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1625),
.B(n_1620),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1637),
.B(n_1611),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1622),
.B(n_1586),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1621),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1623),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1622),
.B(n_1595),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1634),
.B(n_1601),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1626),
.B(n_1595),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1630),
.Y(n_1664)
);

NAND3xp33_ASAP7_75t_SL g1665 ( 
.A(n_1628),
.B(n_1587),
.C(n_1609),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1631),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1635),
.Y(n_1667)
);

AOI21xp33_ASAP7_75t_L g1668 ( 
.A1(n_1648),
.A2(n_1629),
.B(n_1636),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1626),
.B(n_1596),
.Y(n_1669)
);

INVx1_ASAP7_75t_SL g1670 ( 
.A(n_1632),
.Y(n_1670)
);

AOI221xp5_ASAP7_75t_L g1671 ( 
.A1(n_1633),
.A2(n_1609),
.B1(n_1559),
.B2(n_1589),
.C(n_1530),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1633),
.B(n_1596),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1643),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_SL g1674 ( 
.A1(n_1642),
.A2(n_1649),
.B1(n_1652),
.B2(n_1503),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1646),
.Y(n_1675)
);

AOI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1642),
.A2(n_1503),
.B1(n_1512),
.B2(n_1487),
.Y(n_1676)
);

OAI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1641),
.A2(n_1599),
.B1(n_1613),
.B2(n_1562),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1652),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1624),
.B(n_1612),
.Y(n_1679)
);

OAI221xp5_ASAP7_75t_L g1680 ( 
.A1(n_1674),
.A2(n_1649),
.B1(n_1654),
.B2(n_1559),
.C(n_1605),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1655),
.B(n_1624),
.Y(n_1681)
);

AOI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1670),
.A2(n_1512),
.B1(n_1654),
.B2(n_1503),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1655),
.B(n_1638),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1659),
.Y(n_1684)
);

INVx1_ASAP7_75t_SL g1685 ( 
.A(n_1678),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_SL g1686 ( 
.A(n_1657),
.B(n_1672),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1656),
.B(n_1638),
.Y(n_1687)
);

AOI21xp33_ASAP7_75t_L g1688 ( 
.A1(n_1658),
.A2(n_1651),
.B(n_1654),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1671),
.A2(n_1641),
.B1(n_1640),
.B2(n_1650),
.Y(n_1689)
);

O2A1O1Ixp33_ASAP7_75t_L g1690 ( 
.A1(n_1668),
.A2(n_1588),
.B(n_1639),
.C(n_1644),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1659),
.Y(n_1691)
);

AOI21x1_ASAP7_75t_L g1692 ( 
.A1(n_1660),
.A2(n_1651),
.B(n_1654),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1663),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1669),
.B(n_1641),
.Y(n_1694)
);

AOI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1676),
.A2(n_1512),
.B1(n_1503),
.B2(n_1486),
.Y(n_1695)
);

AOI321xp33_ASAP7_75t_SL g1696 ( 
.A1(n_1665),
.A2(n_1640),
.A3(n_1645),
.B1(n_1627),
.B2(n_1647),
.C(n_1653),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1679),
.B(n_1640),
.Y(n_1697)
);

OAI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1661),
.A2(n_1537),
.B1(n_1647),
.B2(n_1617),
.C(n_1602),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1684),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1686),
.B(n_1664),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1694),
.B(n_1662),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1684),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1683),
.Y(n_1703)
);

INVxp67_ASAP7_75t_L g1704 ( 
.A(n_1681),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1694),
.B(n_1662),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1685),
.B(n_1666),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1687),
.B(n_1667),
.Y(n_1707)
);

AND2x4_ASAP7_75t_SL g1708 ( 
.A(n_1693),
.B(n_1673),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1692),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1691),
.Y(n_1710)
);

A2O1A1Ixp33_ASAP7_75t_L g1711 ( 
.A1(n_1700),
.A2(n_1690),
.B(n_1680),
.C(n_1682),
.Y(n_1711)
);

NAND4xp25_ASAP7_75t_L g1712 ( 
.A(n_1700),
.B(n_1696),
.C(n_1697),
.D(n_1689),
.Y(n_1712)
);

NOR2x1_ASAP7_75t_SL g1713 ( 
.A(n_1701),
.B(n_1675),
.Y(n_1713)
);

NOR3xp33_ASAP7_75t_L g1714 ( 
.A(n_1706),
.B(n_1688),
.C(n_1698),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1701),
.B(n_1542),
.Y(n_1715)
);

NAND3xp33_ASAP7_75t_SL g1716 ( 
.A(n_1709),
.B(n_1695),
.C(n_1677),
.Y(n_1716)
);

NOR3xp33_ASAP7_75t_L g1717 ( 
.A(n_1704),
.B(n_1617),
.C(n_1618),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1705),
.Y(n_1718)
);

AOI221xp5_ASAP7_75t_L g1719 ( 
.A1(n_1709),
.A2(n_1530),
.B1(n_1569),
.B2(n_1618),
.C(n_1604),
.Y(n_1719)
);

OAI211xp5_ASAP7_75t_SL g1720 ( 
.A1(n_1711),
.A2(n_1703),
.B(n_1699),
.C(n_1702),
.Y(n_1720)
);

AOI222xp33_ASAP7_75t_L g1721 ( 
.A1(n_1716),
.A2(n_1710),
.B1(n_1708),
.B2(n_1705),
.C1(n_1707),
.C2(n_1486),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1718),
.B(n_1708),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1712),
.A2(n_1569),
.B(n_1604),
.Y(n_1723)
);

AOI221x1_ASAP7_75t_L g1724 ( 
.A1(n_1714),
.A2(n_1562),
.B1(n_1518),
.B2(n_1558),
.C(n_1566),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1722),
.Y(n_1725)
);

O2A1O1Ixp5_ASAP7_75t_L g1726 ( 
.A1(n_1723),
.A2(n_1715),
.B(n_1720),
.C(n_1713),
.Y(n_1726)
);

AOI222xp33_ASAP7_75t_L g1727 ( 
.A1(n_1721),
.A2(n_1719),
.B1(n_1717),
.B2(n_1486),
.C1(n_1487),
.C2(n_1552),
.Y(n_1727)
);

AOI221xp5_ASAP7_75t_L g1728 ( 
.A1(n_1724),
.A2(n_1517),
.B1(n_1518),
.B2(n_1555),
.C(n_1487),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1722),
.Y(n_1729)
);

AOI211xp5_ASAP7_75t_L g1730 ( 
.A1(n_1720),
.A2(n_1438),
.B(n_1567),
.C(n_1435),
.Y(n_1730)
);

NOR4xp25_ASAP7_75t_L g1731 ( 
.A(n_1725),
.B(n_1567),
.C(n_1615),
.D(n_1614),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1729),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1730),
.B(n_1560),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1726),
.Y(n_1734)
);

XOR2x2_ASAP7_75t_L g1735 ( 
.A(n_1728),
.B(n_1727),
.Y(n_1735)
);

AOI221xp5_ASAP7_75t_L g1736 ( 
.A1(n_1734),
.A2(n_1731),
.B1(n_1733),
.B2(n_1732),
.C(n_1735),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_SL g1737 ( 
.A(n_1731),
.B(n_1616),
.Y(n_1737)
);

OAI322xp33_ASAP7_75t_L g1738 ( 
.A1(n_1734),
.A2(n_1616),
.A3(n_1615),
.B1(n_1576),
.B2(n_1564),
.C1(n_1517),
.C2(n_1538),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1737),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1739),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1740),
.A2(n_1736),
.B1(n_1738),
.B2(n_1576),
.Y(n_1741)
);

CKINVDCx20_ASAP7_75t_R g1742 ( 
.A(n_1741),
.Y(n_1742)
);

AOI21xp5_ASAP7_75t_L g1743 ( 
.A1(n_1742),
.A2(n_1555),
.B(n_1560),
.Y(n_1743)
);

AOI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1743),
.A2(n_1555),
.B1(n_1560),
.B2(n_1561),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1744),
.B(n_1576),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1745),
.A2(n_1561),
.B1(n_1517),
.B2(n_1565),
.Y(n_1746)
);

AOI221xp5_ASAP7_75t_L g1747 ( 
.A1(n_1746),
.A2(n_1517),
.B1(n_1566),
.B2(n_1565),
.C(n_1538),
.Y(n_1747)
);

AOI211xp5_ASAP7_75t_L g1748 ( 
.A1(n_1747),
.A2(n_1438),
.B(n_1517),
.C(n_1521),
.Y(n_1748)
);


endmodule