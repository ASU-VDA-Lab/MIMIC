module fake_netlist_1_7777_n_19 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_19);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_19;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_7;
INVx5_ASAP7_75t_L g7 ( .A(n_3), .Y(n_7) );
AND2x4_ASAP7_75t_L g8 ( .A(n_5), .B(n_1), .Y(n_8) );
INVx3_ASAP7_75t_L g9 ( .A(n_4), .Y(n_9) );
INVx4_ASAP7_75t_SL g10 ( .A(n_0), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_6), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_2), .Y(n_12) );
INVx3_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
AND2x4_ASAP7_75t_L g14 ( .A(n_10), .B(n_9), .Y(n_14) );
OAI22xp5_ASAP7_75t_L g15 ( .A1(n_13), .A2(n_11), .B1(n_12), .B2(n_7), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_15), .B(n_13), .Y(n_16) );
AOI222xp33_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_7), .B1(n_14), .B2(n_13), .C1(n_10), .C2(n_15), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
endmodule