module fake_jpeg_14278_n_83 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_83);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_83;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_24),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_40),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_30),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_44),
.B(n_35),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_35),
.C(n_30),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_4),
.C(n_5),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_49),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_47),
.A2(n_29),
.B(n_3),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_32),
.B1(n_34),
.B2(n_37),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_35),
.B(n_33),
.C(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_2),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_57),
.Y(n_66)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_61),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_60),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_53),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_22),
.B(n_23),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_50),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_64),
.B(n_25),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_54),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_67),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g67 ( 
.A(n_63),
.B(n_18),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_SL g69 ( 
.A(n_60),
.B(n_20),
.C(n_21),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_71),
.C(n_72),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_74),
.B(n_66),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_67),
.C(n_76),
.Y(n_78)
);

MAJx2_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_75),
.C(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_79),
.B(n_70),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_65),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_62),
.Y(n_83)
);


endmodule