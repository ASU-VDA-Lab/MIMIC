module fake_netlist_6_4668_n_2783 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_507, n_580, n_209, n_367, n_465, n_590, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_557, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_327, n_369, n_597, n_280, n_287, n_353, n_555, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_522, n_466, n_506, n_56, n_360, n_119, n_235, n_536, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_581, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_95, n_311, n_10, n_403, n_253, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_582, n_4, n_199, n_138, n_266, n_296, n_571, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2783);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_590;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_557;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_597;
input n_280;
input n_287;
input n_353;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_536;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_571;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2783;

wire n_992;
wire n_2542;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_2729;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_1591;
wire n_772;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_1467;
wire n_976;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_699;
wire n_1986;
wire n_2397;
wire n_824;
wire n_686;
wire n_757;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2735;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_630;
wire n_2059;
wire n_2198;
wire n_2669;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_792;
wire n_2522;
wire n_1328;
wire n_1957;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_2455;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_2459;
wire n_1111;
wire n_1713;
wire n_715;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_612;
wire n_2641;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2749;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_850;
wire n_690;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_604;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_2733;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2644;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_2619;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_627;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2728;
wire n_2349;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_2767;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_2707;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_2537;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_2517;
wire n_2713;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2590;
wire n_2643;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_765;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_797;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2675;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_614;
wire n_2307;
wire n_2069;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2771;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2718;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_2682;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_683;
wire n_811;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2780;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_1243;
wire n_848;
wire n_2732;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_2781;
wire n_1129;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_1593;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_2420;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2240;
wire n_2656;
wire n_2278;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_2755;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_2740;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2716;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2541;
wire n_654;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_2406;
wire n_2390;
wire n_806;
wire n_959;
wire n_879;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_1045;
wire n_706;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_2695;
wire n_743;
wire n_766;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_2671;
wire n_2761;
wire n_2715;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_646;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_2587;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_2752;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2186;
wire n_2163;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_2528;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_814;
wire n_2746;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_2076;
wire n_2736;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_1114;
wire n_1848;
wire n_1147;
wire n_763;
wire n_1785;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_744;
wire n_971;
wire n_2702;
wire n_946;
wire n_761;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_2741;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2255;
wire n_2112;
wire n_1464;
wire n_1737;
wire n_653;
wire n_2430;
wire n_1414;
wire n_908;
wire n_752;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_839;
wire n_2437;
wire n_2743;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_1058;
wire n_854;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_719;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_2600;
wire n_984;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_1996;
wire n_2367;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_849;
wire n_2662;
wire n_753;
wire n_1753;
wire n_2471;
wire n_2540;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_2774;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_2659;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx10_ASAP7_75t_L g599 ( 
.A(n_112),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_98),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_416),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_466),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_442),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_596),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_440),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_148),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_59),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_330),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_182),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_347),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_444),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_586),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_201),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_332),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_579),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_513),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_224),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_315),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_497),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_522),
.Y(n_620)
);

CKINVDCx16_ASAP7_75t_R g621 ( 
.A(n_506),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_232),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_455),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_322),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_448),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_144),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_306),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_303),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_452),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_571),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_172),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_63),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_384),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_367),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_564),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_35),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_502),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_18),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_219),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_211),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_340),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_581),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_429),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_28),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_306),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_167),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_521),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_233),
.Y(n_648)
);

CKINVDCx16_ASAP7_75t_R g649 ( 
.A(n_98),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_325),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_101),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_292),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_247),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_303),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_319),
.Y(n_655)
);

CKINVDCx20_ASAP7_75t_R g656 ( 
.A(n_297),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_598),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_438),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_123),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_20),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_19),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_205),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_418),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_361),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_64),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_456),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_234),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_207),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_278),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_221),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_143),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_480),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_267),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_53),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_18),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_569),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_271),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_308),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_432),
.Y(n_679)
);

CKINVDCx14_ASAP7_75t_R g680 ( 
.A(n_426),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_52),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_301),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_291),
.Y(n_683)
);

INVxp67_ASAP7_75t_SL g684 ( 
.A(n_357),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_194),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_449),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_563),
.Y(n_687)
);

CKINVDCx16_ASAP7_75t_R g688 ( 
.A(n_330),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_582),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_356),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_296),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_472),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_566),
.Y(n_693)
);

BUFx8_ASAP7_75t_SL g694 ( 
.A(n_19),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_110),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_96),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_560),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_197),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_206),
.Y(n_699)
);

CKINVDCx16_ASAP7_75t_R g700 ( 
.A(n_474),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_424),
.Y(n_701)
);

CKINVDCx16_ASAP7_75t_R g702 ( 
.A(n_531),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_507),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_329),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_407),
.Y(n_705)
);

BUFx10_ASAP7_75t_L g706 ( 
.A(n_58),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_148),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_349),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_496),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_458),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_590),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_583),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_572),
.Y(n_713)
);

BUFx10_ASAP7_75t_L g714 ( 
.A(n_147),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_504),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_382),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_27),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_548),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_59),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_518),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_475),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_459),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_258),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_595),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_30),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_83),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_319),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_576),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_379),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_464),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_261),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_43),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_199),
.Y(n_733)
);

CKINVDCx20_ASAP7_75t_R g734 ( 
.A(n_26),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_580),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_168),
.Y(n_736)
);

CKINVDCx16_ASAP7_75t_R g737 ( 
.A(n_399),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_243),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_575),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_443),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_338),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_589),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_21),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_539),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_549),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_565),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_63),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_423),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_383),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_445),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_97),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_337),
.Y(n_752)
);

BUFx10_ASAP7_75t_L g753 ( 
.A(n_302),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_570),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_329),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_30),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_246),
.Y(n_757)
);

INVx1_ASAP7_75t_SL g758 ( 
.A(n_516),
.Y(n_758)
);

BUFx5_ASAP7_75t_L g759 ( 
.A(n_70),
.Y(n_759)
);

CKINVDCx14_ASAP7_75t_R g760 ( 
.A(n_131),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_28),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_240),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_500),
.Y(n_763)
);

CKINVDCx16_ASAP7_75t_R g764 ( 
.A(n_413),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_391),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_89),
.Y(n_766)
);

BUFx10_ASAP7_75t_L g767 ( 
.A(n_453),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_457),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_192),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_574),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_6),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_376),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_508),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_282),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_216),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_197),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_246),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_446),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_447),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_75),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_137),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_262),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_415),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_115),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_540),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_505),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_322),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_545),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_551),
.Y(n_789)
);

CKINVDCx20_ASAP7_75t_R g790 ( 
.A(n_243),
.Y(n_790)
);

INVx1_ASAP7_75t_SL g791 ( 
.A(n_501),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_454),
.Y(n_792)
);

CKINVDCx14_ASAP7_75t_R g793 ( 
.A(n_451),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_117),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_311),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_519),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_492),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_384),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_379),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_289),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_372),
.Y(n_801)
);

INVx1_ASAP7_75t_SL g802 ( 
.A(n_535),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_328),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_170),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_573),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_450),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_76),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_543),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_460),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_484),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_219),
.Y(n_811)
);

BUFx10_ASAP7_75t_L g812 ( 
.A(n_468),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_308),
.Y(n_813)
);

BUFx10_ASAP7_75t_L g814 ( 
.A(n_541),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_217),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_442),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_402),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_103),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_533),
.Y(n_819)
);

CKINVDCx20_ASAP7_75t_R g820 ( 
.A(n_476),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_441),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_337),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_331),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_128),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_491),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_432),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_177),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_520),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_366),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_203),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_295),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_759),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_759),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_759),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_694),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_759),
.Y(n_836)
);

CKINVDCx16_ASAP7_75t_R g837 ( 
.A(n_649),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_759),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_694),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_759),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_680),
.Y(n_841)
);

BUFx3_ASAP7_75t_L g842 ( 
.A(n_602),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_602),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_759),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_705),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_624),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_705),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_733),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_624),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_680),
.Y(n_850)
);

CKINVDCx20_ASAP7_75t_R g851 ( 
.A(n_765),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_733),
.Y(n_852)
);

INVx1_ASAP7_75t_SL g853 ( 
.A(n_606),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_624),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_624),
.Y(n_855)
);

CKINVDCx16_ASAP7_75t_R g856 ( 
.A(n_688),
.Y(n_856)
);

INVxp33_ASAP7_75t_SL g857 ( 
.A(n_665),
.Y(n_857)
);

CKINVDCx20_ASAP7_75t_R g858 ( 
.A(n_765),
.Y(n_858)
);

INVxp67_ASAP7_75t_SL g859 ( 
.A(n_735),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_751),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_761),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_760),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_761),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_794),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_794),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_829),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_829),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_626),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_626),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_626),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_793),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_626),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_682),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_793),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_618),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_682),
.Y(n_876)
);

CKINVDCx14_ASAP7_75t_R g877 ( 
.A(n_708),
.Y(n_877)
);

CKINVDCx16_ASAP7_75t_R g878 ( 
.A(n_737),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_682),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_682),
.Y(n_880)
);

INVxp67_ASAP7_75t_L g881 ( 
.A(n_599),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_764),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_600),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_685),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_685),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_601),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_685),
.Y(n_887)
);

CKINVDCx16_ASAP7_75t_R g888 ( 
.A(n_621),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_685),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_719),
.Y(n_890)
);

CKINVDCx16_ASAP7_75t_R g891 ( 
.A(n_700),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_719),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_719),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_603),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_719),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_607),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_735),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_613),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_790),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_808),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_599),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_756),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_622),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_756),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_756),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_756),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_769),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_769),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_769),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_769),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_605),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_628),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_790),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_631),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_609),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_611),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_619),
.Y(n_917)
);

INVxp33_ASAP7_75t_L g918 ( 
.A(n_611),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_614),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_808),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_623),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_629),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_632),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_634),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_644),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_812),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_648),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_650),
.Y(n_928)
);

CKINVDCx16_ASAP7_75t_R g929 ( 
.A(n_702),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_652),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_653),
.Y(n_931)
);

CKINVDCx16_ASAP7_75t_R g932 ( 
.A(n_837),
.Y(n_932)
);

INVxp67_ASAP7_75t_L g933 ( 
.A(n_886),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_883),
.Y(n_934)
);

INVxp67_ASAP7_75t_SL g935 ( 
.A(n_842),
.Y(n_935)
);

CKINVDCx20_ASAP7_75t_R g936 ( 
.A(n_851),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_868),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_870),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_872),
.Y(n_939)
);

NOR2xp67_ASAP7_75t_L g940 ( 
.A(n_883),
.B(n_647),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_894),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_873),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_876),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_880),
.Y(n_944)
);

CKINVDCx20_ASAP7_75t_R g945 ( 
.A(n_851),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_896),
.Y(n_946)
);

CKINVDCx20_ASAP7_75t_R g947 ( 
.A(n_858),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_884),
.Y(n_948)
);

INVx1_ASAP7_75t_SL g949 ( 
.A(n_858),
.Y(n_949)
);

CKINVDCx16_ASAP7_75t_R g950 ( 
.A(n_856),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_887),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_889),
.Y(n_952)
);

NOR2xp67_ASAP7_75t_L g953 ( 
.A(n_894),
.B(n_616),
.Y(n_953)
);

CKINVDCx20_ASAP7_75t_R g954 ( 
.A(n_899),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_890),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_895),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_902),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_898),
.Y(n_958)
);

CKINVDCx20_ASAP7_75t_R g959 ( 
.A(n_899),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_882),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_898),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_904),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_905),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_903),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_903),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_906),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_842),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_907),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_908),
.Y(n_969)
);

CKINVDCx20_ASAP7_75t_R g970 ( 
.A(n_913),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_912),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_913),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_909),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_912),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_910),
.Y(n_975)
);

CKINVDCx20_ASAP7_75t_R g976 ( 
.A(n_878),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_914),
.Y(n_977)
);

CKINVDCx20_ASAP7_75t_R g978 ( 
.A(n_835),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_914),
.Y(n_979)
);

CKINVDCx20_ASAP7_75t_R g980 ( 
.A(n_835),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_882),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_846),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_839),
.Y(n_983)
);

INVxp67_ASAP7_75t_SL g984 ( 
.A(n_843),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_839),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_888),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_841),
.B(n_758),
.Y(n_987)
);

INVxp67_ASAP7_75t_SL g988 ( 
.A(n_843),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_891),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_841),
.B(n_791),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_929),
.Y(n_991)
);

INVxp67_ASAP7_75t_SL g992 ( 
.A(n_897),
.Y(n_992)
);

INVxp67_ASAP7_75t_L g993 ( 
.A(n_896),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_846),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_849),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_850),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_967),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_934),
.Y(n_998)
);

INVx2_ASAP7_75t_SL g999 ( 
.A(n_967),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_937),
.Y(n_1000)
);

CKINVDCx8_ASAP7_75t_R g1001 ( 
.A(n_932),
.Y(n_1001)
);

NAND2xp33_ASAP7_75t_SL g1002 ( 
.A(n_996),
.B(n_820),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_938),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_939),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_935),
.B(n_897),
.Y(n_1005)
);

BUFx8_ASAP7_75t_L g1006 ( 
.A(n_950),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_942),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_943),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_944),
.Y(n_1009)
);

CKINVDCx20_ASAP7_75t_R g1010 ( 
.A(n_936),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_982),
.B(n_832),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_953),
.Y(n_1012)
);

BUFx8_ASAP7_75t_L g1013 ( 
.A(n_948),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_976),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_946),
.Y(n_1015)
);

CKINVDCx20_ASAP7_75t_R g1016 ( 
.A(n_976),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_994),
.B(n_833),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_941),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_951),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_952),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_936),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_955),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_993),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_984),
.B(n_862),
.Y(n_1024)
);

OA21x2_ASAP7_75t_L g1025 ( 
.A1(n_995),
.A2(n_838),
.B(n_834),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_956),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_957),
.Y(n_1027)
);

AND2x2_ASAP7_75t_SL g1028 ( 
.A(n_987),
.B(n_604),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_962),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_963),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_990),
.A2(n_857),
.B1(n_831),
.B2(n_816),
.Y(n_1031)
);

XOR2xp5_ASAP7_75t_L g1032 ( 
.A(n_986),
.B(n_720),
.Y(n_1032)
);

AND2x6_ASAP7_75t_L g1033 ( 
.A(n_966),
.B(n_604),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_958),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_968),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_969),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_973),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_975),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_988),
.B(n_871),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_961),
.Y(n_1040)
);

CKINVDCx20_ASAP7_75t_R g1041 ( 
.A(n_945),
.Y(n_1041)
);

NOR2x1_ASAP7_75t_L g1042 ( 
.A(n_940),
.B(n_721),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_992),
.B(n_871),
.Y(n_1043)
);

AND2x2_ASAP7_75t_SL g1044 ( 
.A(n_960),
.B(n_615),
.Y(n_1044)
);

NAND2xp33_ASAP7_75t_L g1045 ( 
.A(n_996),
.B(n_874),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_933),
.B(n_900),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_949),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_964),
.B(n_874),
.Y(n_1048)
);

AND2x6_ASAP7_75t_L g1049 ( 
.A(n_965),
.B(n_615),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_971),
.A2(n_836),
.B(n_840),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_974),
.B(n_900),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_977),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_979),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_989),
.B(n_920),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_981),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_991),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_978),
.B(n_877),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_978),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_980),
.Y(n_1059)
);

CKINVDCx20_ASAP7_75t_R g1060 ( 
.A(n_945),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_980),
.A2(n_831),
.B1(n_816),
.B2(n_853),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_983),
.B(n_859),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_983),
.Y(n_1063)
);

NOR2x1_ASAP7_75t_L g1064 ( 
.A(n_985),
.B(n_754),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_985),
.Y(n_1065)
);

INVx4_ASAP7_75t_L g1066 ( 
.A(n_947),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_972),
.B(n_642),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_972),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_947),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_SL g1070 ( 
.A1(n_970),
.A2(n_641),
.B1(n_643),
.B2(n_638),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_954),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_954),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_959),
.Y(n_1073)
);

AOI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_959),
.A2(n_763),
.B1(n_820),
.B2(n_875),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_970),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_SL g1076 ( 
.A1(n_976),
.A2(n_656),
.B1(n_670),
.B2(n_654),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_937),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_937),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_976),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_937),
.Y(n_1080)
);

HB1xp67_ASAP7_75t_L g1081 ( 
.A(n_967),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_937),
.Y(n_1082)
);

AND2x4_ASAP7_75t_SL g1083 ( 
.A(n_976),
.B(n_812),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1025),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_1010),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_1006),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_1025),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1003),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1011),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_1012),
.B(n_1028),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_1044),
.B(n_619),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_997),
.Y(n_1092)
);

INVxp67_ASAP7_75t_SL g1093 ( 
.A(n_1081),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1004),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_1006),
.Y(n_1095)
);

AND2x6_ASAP7_75t_L g1096 ( 
.A(n_1042),
.B(n_1024),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1009),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1020),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1011),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_1017),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1026),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1017),
.Y(n_1102)
);

NOR3xp33_ASAP7_75t_L g1103 ( 
.A(n_1031),
.B(n_901),
.C(n_881),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1029),
.Y(n_1104)
);

INVx2_ASAP7_75t_SL g1105 ( 
.A(n_1005),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1050),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1000),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1038),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_1012),
.B(n_875),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_1044),
.B(n_619),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_1007),
.Y(n_1111)
);

INVxp33_ASAP7_75t_L g1112 ( 
.A(n_1047),
.Y(n_1112)
);

INVx4_ASAP7_75t_L g1113 ( 
.A(n_997),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1077),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_1039),
.B(n_1015),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_1047),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1022),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_997),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_1007),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1027),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1078),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1080),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1030),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_1005),
.B(n_619),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_1039),
.B(n_926),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1082),
.Y(n_1126)
);

AND3x1_ASAP7_75t_L g1127 ( 
.A(n_1074),
.B(n_847),
.C(n_845),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_1008),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1037),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1008),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_1062),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1008),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1019),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1049),
.B(n_642),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_1015),
.B(n_926),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1019),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1049),
.B(n_693),
.Y(n_1137)
);

INVx8_ASAP7_75t_L g1138 ( 
.A(n_1049),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1019),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_1051),
.B(n_730),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1043),
.B(n_920),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1035),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1035),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1081),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1035),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_1051),
.B(n_1036),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_1036),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_998),
.Y(n_1148)
);

CKINVDCx6p67_ASAP7_75t_R g1149 ( 
.A(n_1016),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1036),
.Y(n_1150)
);

CKINVDCx6p67_ASAP7_75t_R g1151 ( 
.A(n_1079),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1033),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_1033),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1049),
.B(n_693),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1033),
.Y(n_1155)
);

INVxp67_ASAP7_75t_SL g1156 ( 
.A(n_999),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1033),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_1021),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1023),
.B(n_918),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1046),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1033),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1048),
.B(n_802),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1046),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1054),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1067),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_1054),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1053),
.B(n_730),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1048),
.B(n_610),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1067),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1055),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1052),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_1018),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1056),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1040),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1040),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1053),
.B(n_848),
.Y(n_1176)
);

NOR2x1p5_ASAP7_75t_L g1177 ( 
.A(n_1053),
.B(n_684),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1013),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1013),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1045),
.Y(n_1180)
);

AND3x2_ASAP7_75t_L g1181 ( 
.A(n_1014),
.B(n_608),
.C(n_625),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1002),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1002),
.Y(n_1183)
);

AND2x6_ASAP7_75t_L g1184 ( 
.A(n_1064),
.B(n_713),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1083),
.Y(n_1185)
);

INVxp67_ASAP7_75t_R g1186 ( 
.A(n_1076),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_1041),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1072),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1001),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1034),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1068),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1069),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_1060),
.Y(n_1193)
);

INVx1_ASAP7_75t_SL g1194 ( 
.A(n_1010),
.Y(n_1194)
);

AND3x2_ASAP7_75t_L g1195 ( 
.A(n_1057),
.B(n_669),
.C(n_625),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_1031),
.B(n_730),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1071),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1075),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1057),
.B(n_796),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1073),
.Y(n_1200)
);

OAI22xp33_ASAP7_75t_SL g1201 ( 
.A1(n_1061),
.A2(n_635),
.B1(n_689),
.B2(n_676),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1073),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_1073),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1066),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1058),
.Y(n_1205)
);

INVxp33_ASAP7_75t_SL g1206 ( 
.A(n_1032),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1059),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_1066),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_1063),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1065),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1061),
.B(n_796),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1070),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1063),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_1063),
.Y(n_1214)
);

INVx2_ASAP7_75t_SL g1215 ( 
.A(n_1005),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1003),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1105),
.B(n_911),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1111),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1203),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1107),
.Y(n_1220)
);

INVx4_ASAP7_75t_L g1221 ( 
.A(n_1118),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1111),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1111),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_1116),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_1131),
.B(n_852),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1089),
.B(n_715),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1119),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1119),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1119),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1168),
.B(n_696),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1203),
.Y(n_1231)
);

INVx1_ASAP7_75t_SL g1232 ( 
.A(n_1112),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_1203),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1107),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1105),
.B(n_915),
.Y(n_1235)
);

NAND3x1_ASAP7_75t_L g1236 ( 
.A(n_1212),
.B(n_731),
.C(n_701),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1128),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1162),
.B(n_734),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1084),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1202),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_1203),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1088),
.Y(n_1242)
);

BUFx10_ASAP7_75t_L g1243 ( 
.A(n_1148),
.Y(n_1243)
);

AND2x4_ASAP7_75t_L g1244 ( 
.A(n_1215),
.B(n_919),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1117),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1128),
.Y(n_1246)
);

INVx4_ASAP7_75t_L g1247 ( 
.A(n_1118),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1094),
.Y(n_1248)
);

INVx4_ASAP7_75t_L g1249 ( 
.A(n_1118),
.Y(n_1249)
);

BUFx4f_ASAP7_75t_L g1250 ( 
.A(n_1208),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1202),
.Y(n_1251)
);

INVxp67_ASAP7_75t_SL g1252 ( 
.A(n_1128),
.Y(n_1252)
);

AND2x6_ASAP7_75t_L g1253 ( 
.A(n_1152),
.B(n_718),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1117),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1115),
.B(n_752),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1097),
.Y(n_1256)
);

INVx4_ASAP7_75t_L g1257 ( 
.A(n_1128),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1084),
.Y(n_1258)
);

INVx4_ASAP7_75t_L g1259 ( 
.A(n_1113),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1089),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1209),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1171),
.B(n_612),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1099),
.B(n_728),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1112),
.B(n_617),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_1092),
.Y(n_1265)
);

AND2x6_ASAP7_75t_SL g1266 ( 
.A(n_1190),
.B(n_658),
.Y(n_1266)
);

INVx1_ASAP7_75t_SL g1267 ( 
.A(n_1194),
.Y(n_1267)
);

AND2x6_ASAP7_75t_L g1268 ( 
.A(n_1152),
.B(n_1155),
.Y(n_1268)
);

INVx5_ASAP7_75t_L g1269 ( 
.A(n_1208),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_1148),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1159),
.B(n_1141),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1090),
.B(n_815),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1213),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1099),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1213),
.Y(n_1275)
);

OR2x2_ASAP7_75t_L g1276 ( 
.A(n_1109),
.B(n_860),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1098),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_1158),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1120),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1125),
.B(n_633),
.Y(n_1280)
);

OR2x6_ASAP7_75t_L g1281 ( 
.A(n_1208),
.B(n_861),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1120),
.Y(n_1282)
);

OAI22x1_ASAP7_75t_SL g1283 ( 
.A1(n_1206),
.A2(n_636),
.B1(n_645),
.B2(n_639),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1101),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1141),
.B(n_863),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1123),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1104),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1108),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1093),
.B(n_646),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1114),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1121),
.Y(n_1291)
);

INVx5_ASAP7_75t_L g1292 ( 
.A(n_1208),
.Y(n_1292)
);

INVx4_ASAP7_75t_L g1293 ( 
.A(n_1113),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1100),
.B(n_1102),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1122),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1130),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1102),
.B(n_745),
.Y(n_1297)
);

NAND2x1p5_ASAP7_75t_L g1298 ( 
.A(n_1113),
.B(n_921),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1123),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1215),
.B(n_922),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1164),
.B(n_923),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1129),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1176),
.B(n_864),
.Y(n_1303)
);

AND2x2_ASAP7_75t_SL g1304 ( 
.A(n_1187),
.B(n_1193),
.Y(n_1304)
);

BUFx10_ASAP7_75t_L g1305 ( 
.A(n_1172),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1129),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1087),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1164),
.B(n_1166),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1174),
.B(n_620),
.Y(n_1309)
);

AND2x4_ASAP7_75t_L g1310 ( 
.A(n_1164),
.B(n_924),
.Y(n_1310)
);

INVx4_ASAP7_75t_L g1311 ( 
.A(n_1092),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1165),
.A2(n_786),
.B1(n_788),
.B2(n_770),
.Y(n_1312)
);

OAI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1169),
.A2(n_805),
.B1(n_810),
.B2(n_797),
.Y(n_1313)
);

INVx5_ASAP7_75t_L g1314 ( 
.A(n_1096),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1172),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1087),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1166),
.B(n_925),
.Y(n_1317)
);

NOR2x1p5_ASAP7_75t_L g1318 ( 
.A(n_1166),
.B(n_1178),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1149),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1160),
.B(n_927),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_SL g1321 ( 
.A(n_1174),
.B(n_630),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1087),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1126),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1176),
.B(n_865),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1175),
.Y(n_1325)
);

INVx8_ASAP7_75t_L g1326 ( 
.A(n_1184),
.Y(n_1326)
);

AO21x2_ASAP7_75t_L g1327 ( 
.A1(n_1091),
.A2(n_828),
.B(n_844),
.Y(n_1327)
);

INVx5_ASAP7_75t_L g1328 ( 
.A(n_1096),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1135),
.B(n_866),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1169),
.B(n_637),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_1149),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_SL g1332 ( 
.A(n_1175),
.B(n_657),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1130),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1132),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1091),
.A2(n_730),
.B1(n_836),
.B2(n_814),
.Y(n_1335)
);

INVx5_ASAP7_75t_L g1336 ( 
.A(n_1096),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1216),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1096),
.B(n_1132),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1133),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1133),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_1151),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1200),
.Y(n_1342)
);

INVx5_ASAP7_75t_L g1343 ( 
.A(n_1096),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1163),
.B(n_928),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1144),
.B(n_867),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1096),
.B(n_672),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1192),
.B(n_599),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1182),
.B(n_651),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1173),
.B(n_930),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1110),
.A2(n_692),
.B1(n_697),
.B2(n_687),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1136),
.B(n_1139),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1192),
.B(n_931),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1110),
.A2(n_814),
.B1(n_812),
.B2(n_640),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1136),
.Y(n_1354)
);

INVx5_ASAP7_75t_L g1355 ( 
.A(n_1184),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1139),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1204),
.B(n_703),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1197),
.B(n_706),
.Y(n_1358)
);

AO21x2_ASAP7_75t_L g1359 ( 
.A1(n_1134),
.A2(n_855),
.B(n_854),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1142),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_SL g1361 ( 
.A(n_1204),
.B(n_709),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1142),
.B(n_711),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1143),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1143),
.Y(n_1364)
);

BUFx8_ASAP7_75t_SL g1365 ( 
.A(n_1085),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1177),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1197),
.B(n_916),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1150),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1146),
.B(n_660),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1150),
.Y(n_1370)
);

BUFx6f_ASAP7_75t_L g1371 ( 
.A(n_1147),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1146),
.B(n_661),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_SL g1373 ( 
.A(n_1204),
.B(n_712),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1198),
.B(n_706),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1183),
.B(n_655),
.Y(n_1375)
);

BUFx10_ASAP7_75t_L g1376 ( 
.A(n_1195),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1198),
.B(n_1210),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1085),
.Y(n_1378)
);

AND2x6_ASAP7_75t_L g1379 ( 
.A(n_1155),
.B(n_669),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1188),
.Y(n_1380)
);

INVx3_ASAP7_75t_L g1381 ( 
.A(n_1147),
.Y(n_1381)
);

INVx4_ASAP7_75t_L g1382 ( 
.A(n_1147),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1210),
.B(n_706),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1145),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1106),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1106),
.Y(n_1386)
);

BUFx2_ASAP7_75t_L g1387 ( 
.A(n_1214),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_1157),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1157),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1205),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1180),
.B(n_724),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1207),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1199),
.B(n_714),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1161),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1170),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1156),
.B(n_1185),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1161),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1124),
.Y(n_1398)
);

INVx5_ASAP7_75t_L g1399 ( 
.A(n_1184),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1153),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1124),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1191),
.Y(n_1402)
);

INVx5_ASAP7_75t_L g1403 ( 
.A(n_1184),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1137),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1103),
.B(n_714),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1154),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1140),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1185),
.B(n_714),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1220),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1377),
.Y(n_1410)
);

NAND3xp33_ASAP7_75t_L g1411 ( 
.A(n_1238),
.B(n_1196),
.C(n_1211),
.Y(n_1411)
);

INVxp33_ASAP7_75t_L g1412 ( 
.A(n_1224),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1260),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1271),
.B(n_1186),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1234),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1294),
.B(n_1184),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1260),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1245),
.Y(n_1418)
);

O2A1O1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1230),
.A2(n_1196),
.B(n_1201),
.C(n_1140),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1274),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_SL g1421 ( 
.A(n_1269),
.B(n_1127),
.Y(n_1421)
);

OAI221xp5_ASAP7_75t_L g1422 ( 
.A1(n_1255),
.A2(n_1189),
.B1(n_1179),
.B2(n_1178),
.C(n_1167),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_SL g1423 ( 
.A(n_1269),
.B(n_1292),
.Y(n_1423)
);

NAND3xp33_ASAP7_75t_L g1424 ( 
.A(n_1280),
.B(n_1167),
.C(n_1181),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1274),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1302),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1382),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1272),
.B(n_1184),
.Y(n_1428)
);

NAND3xp33_ASAP7_75t_L g1429 ( 
.A(n_1348),
.B(n_1375),
.C(n_1393),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1302),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1232),
.B(n_1151),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1219),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1292),
.B(n_1179),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1292),
.B(n_1250),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1306),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1254),
.Y(n_1436)
);

INVxp67_ASAP7_75t_L g1437 ( 
.A(n_1387),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1242),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1248),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1303),
.A2(n_1206),
.B1(n_1138),
.B2(n_742),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1329),
.B(n_1138),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1324),
.B(n_739),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1323),
.A2(n_814),
.B1(n_746),
.B2(n_773),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1285),
.B(n_744),
.Y(n_1444)
);

NOR2xp67_ASAP7_75t_L g1445 ( 
.A(n_1270),
.B(n_1086),
.Y(n_1445)
);

AOI221xp5_ASAP7_75t_L g1446 ( 
.A1(n_1405),
.A2(n_1264),
.B1(n_1289),
.B2(n_1353),
.C(n_1277),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1256),
.B(n_785),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1284),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1279),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1287),
.B(n_789),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1282),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1382),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1288),
.B(n_809),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1267),
.B(n_1086),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1290),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1239),
.B(n_849),
.Y(n_1456)
);

NOR2x1p5_ASAP7_75t_L g1457 ( 
.A(n_1315),
.B(n_1095),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_SL g1458 ( 
.A(n_1396),
.B(n_1095),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1396),
.B(n_819),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_SL g1460 ( 
.A(n_1308),
.B(n_825),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1291),
.B(n_627),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1278),
.B(n_659),
.Y(n_1462)
);

O2A1O1Ixp33_ASAP7_75t_L g1463 ( 
.A1(n_1402),
.A2(n_771),
.B(n_774),
.C(n_732),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1225),
.B(n_916),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1295),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1276),
.B(n_662),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_SL g1467 ( 
.A(n_1308),
.B(n_663),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1380),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1286),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1347),
.B(n_753),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1390),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_SL g1472 ( 
.A(n_1265),
.B(n_664),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_SL g1473 ( 
.A(n_1265),
.B(n_667),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1392),
.Y(n_1474)
);

INVxp67_ASAP7_75t_L g1475 ( 
.A(n_1408),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1239),
.B(n_869),
.Y(n_1476)
);

INVx2_ASAP7_75t_SL g1477 ( 
.A(n_1261),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1349),
.Y(n_1478)
);

NOR2xp67_ASAP7_75t_L g1479 ( 
.A(n_1366),
.B(n_461),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1258),
.B(n_869),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1337),
.B(n_782),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1369),
.B(n_668),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_SL g1483 ( 
.A(n_1259),
.B(n_753),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1299),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1265),
.B(n_671),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1369),
.B(n_674),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_SL g1487 ( 
.A(n_1219),
.B(n_675),
.Y(n_1487)
);

A2O1A1Ixp33_ASAP7_75t_L g1488 ( 
.A1(n_1401),
.A2(n_679),
.B(n_681),
.C(n_666),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1372),
.B(n_677),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1367),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_SL g1491 ( 
.A(n_1219),
.B(n_678),
.Y(n_1491)
);

NAND2xp33_ASAP7_75t_L g1492 ( 
.A(n_1325),
.B(n_686),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1218),
.Y(n_1493)
);

BUFx5_ASAP7_75t_L g1494 ( 
.A(n_1268),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1231),
.B(n_691),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1372),
.B(n_707),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1395),
.B(n_710),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1240),
.B(n_1251),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1358),
.B(n_1374),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1345),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1383),
.B(n_753),
.Y(n_1501)
);

NAND3xp33_ASAP7_75t_L g1502 ( 
.A(n_1226),
.B(n_690),
.C(n_683),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1389),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1389),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1325),
.B(n_722),
.Y(n_1505)
);

INVxp67_ASAP7_75t_L g1506 ( 
.A(n_1378),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1325),
.B(n_723),
.Y(n_1507)
);

INVx8_ASAP7_75t_L g1508 ( 
.A(n_1281),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_SL g1509 ( 
.A(n_1231),
.B(n_725),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1397),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_SL g1511 ( 
.A(n_1231),
.B(n_727),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1273),
.B(n_729),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1275),
.B(n_740),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1301),
.B(n_741),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1342),
.B(n_743),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1307),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1301),
.B(n_748),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1352),
.B(n_749),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1307),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1391),
.B(n_750),
.Y(n_1520)
);

BUFx6f_ASAP7_75t_L g1521 ( 
.A(n_1233),
.Y(n_1521)
);

BUFx6f_ASAP7_75t_L g1522 ( 
.A(n_1241),
.Y(n_1522)
);

INVx4_ASAP7_75t_L g1523 ( 
.A(n_1281),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1304),
.B(n_757),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1243),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1316),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1222),
.Y(n_1527)
);

OAI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1330),
.A2(n_783),
.B1(n_784),
.B2(n_673),
.Y(n_1528)
);

AOI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1310),
.A2(n_768),
.B1(n_772),
.B2(n_766),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1223),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1310),
.B(n_776),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1316),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_1365),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1398),
.A2(n_783),
.B1(n_784),
.B2(n_673),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1317),
.B(n_777),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1317),
.B(n_778),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_SL g1537 ( 
.A(n_1311),
.B(n_779),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1262),
.A2(n_795),
.B1(n_799),
.B2(n_780),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1311),
.B(n_800),
.Y(n_1539)
);

OAI221xp5_ASAP7_75t_L g1540 ( 
.A1(n_1335),
.A2(n_807),
.B1(n_813),
.B2(n_804),
.C(n_803),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_SL g1541 ( 
.A(n_1217),
.B(n_1235),
.Y(n_1541)
);

INVx2_ASAP7_75t_SL g1542 ( 
.A(n_1318),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_SL g1543 ( 
.A(n_1217),
.B(n_817),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1322),
.Y(n_1544)
);

NOR2xp67_ASAP7_75t_L g1545 ( 
.A(n_1319),
.B(n_462),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1223),
.Y(n_1546)
);

AOI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1235),
.A2(n_822),
.B1(n_823),
.B2(n_818),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_SL g1548 ( 
.A(n_1244),
.B(n_824),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1322),
.Y(n_1549)
);

NOR2x1p5_ASAP7_75t_L g1550 ( 
.A(n_1331),
.B(n_827),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_1244),
.B(n_1300),
.Y(n_1551)
);

AOI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1404),
.A2(n_917),
.B(n_885),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1258),
.Y(n_1553)
);

XOR2x2_ASAP7_75t_L g1554 ( 
.A(n_1236),
.B(n_1320),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1263),
.B(n_830),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1297),
.B(n_695),
.Y(n_1556)
);

NAND2xp33_ASAP7_75t_L g1557 ( 
.A(n_1314),
.B(n_787),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1407),
.B(n_698),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1227),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1384),
.B(n_699),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1228),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_SL g1562 ( 
.A(n_1259),
.B(n_767),
.Y(n_1562)
);

AOI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1309),
.A2(n_855),
.B1(n_893),
.B2(n_854),
.Y(n_1563)
);

INVx4_ASAP7_75t_L g1564 ( 
.A(n_1293),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1333),
.B(n_704),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1228),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1229),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1320),
.B(n_767),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1333),
.B(n_1334),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1312),
.A2(n_826),
.B1(n_787),
.B2(n_717),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1334),
.B(n_716),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1394),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1339),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1293),
.B(n_767),
.Y(n_1574)
);

INVxp33_ASAP7_75t_L g1575 ( 
.A(n_1344),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1406),
.B(n_879),
.Y(n_1576)
);

BUFx5_ASAP7_75t_L g1577 ( 
.A(n_1268),
.Y(n_1577)
);

OAI221xp5_ASAP7_75t_L g1578 ( 
.A1(n_1350),
.A2(n_738),
.B1(n_747),
.B2(n_736),
.C(n_726),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1344),
.B(n_755),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1339),
.B(n_879),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_SL g1581 ( 
.A(n_1305),
.B(n_826),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1360),
.B(n_885),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1360),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1314),
.B(n_762),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1364),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1364),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1313),
.A2(n_781),
.B1(n_792),
.B2(n_775),
.Y(n_1587)
);

BUFx3_ASAP7_75t_L g1588 ( 
.A(n_1305),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1368),
.B(n_892),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1394),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1340),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1388),
.B(n_893),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1354),
.B(n_798),
.Y(n_1593)
);

AND2x2_ASAP7_75t_SL g1594 ( 
.A(n_1346),
.B(n_801),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1356),
.B(n_806),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1385),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1363),
.B(n_811),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_SL g1598 ( 
.A(n_1328),
.B(n_821),
.Y(n_1598)
);

INVx5_ASAP7_75t_L g1599 ( 
.A(n_1326),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1429),
.B(n_1341),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1438),
.Y(n_1601)
);

A2O1A1Ixp33_ASAP7_75t_L g1602 ( 
.A1(n_1419),
.A2(n_1338),
.B(n_1332),
.C(n_1321),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1439),
.Y(n_1603)
);

AND2x6_ASAP7_75t_L g1604 ( 
.A(n_1427),
.B(n_1388),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1499),
.B(n_1351),
.Y(n_1605)
);

INVx6_ASAP7_75t_L g1606 ( 
.A(n_1508),
.Y(n_1606)
);

BUFx3_ASAP7_75t_L g1607 ( 
.A(n_1525),
.Y(n_1607)
);

INVxp67_ASAP7_75t_L g1608 ( 
.A(n_1498),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1410),
.B(n_1520),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1412),
.B(n_1283),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1448),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1553),
.Y(n_1612)
);

INVx2_ASAP7_75t_SL g1613 ( 
.A(n_1477),
.Y(n_1613)
);

AOI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1414),
.A2(n_1357),
.B1(n_1373),
.B2(n_1361),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1541),
.B(n_1551),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1503),
.Y(n_1616)
);

BUFx4f_ASAP7_75t_L g1617 ( 
.A(n_1508),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1446),
.B(n_1370),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1411),
.A2(n_1594),
.B1(n_1578),
.B2(n_1466),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_SL g1620 ( 
.A(n_1500),
.B(n_1328),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1504),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1475),
.B(n_1336),
.Y(n_1622)
);

NAND2xp33_ASAP7_75t_L g1623 ( 
.A(n_1411),
.B(n_1336),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1455),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1465),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1470),
.B(n_1376),
.Y(n_1626)
);

BUFx3_ASAP7_75t_L g1627 ( 
.A(n_1588),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1413),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1596),
.Y(n_1629)
);

AOI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1524),
.A2(n_1362),
.B1(n_1376),
.B2(n_1298),
.Y(n_1630)
);

INVx2_ASAP7_75t_SL g1631 ( 
.A(n_1508),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1490),
.B(n_1296),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_R g1633 ( 
.A(n_1533),
.B(n_1336),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1506),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1518),
.B(n_1296),
.Y(n_1635)
);

NOR2x1p5_ASAP7_75t_L g1636 ( 
.A(n_1523),
.B(n_1424),
.Y(n_1636)
);

AND2x6_ASAP7_75t_L g1637 ( 
.A(n_1427),
.B(n_1388),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1555),
.B(n_1252),
.Y(n_1638)
);

A2O1A1Ixp33_ASAP7_75t_L g1639 ( 
.A1(n_1424),
.A2(n_1343),
.B(n_1326),
.C(n_1381),
.Y(n_1639)
);

INVx2_ASAP7_75t_SL g1640 ( 
.A(n_1521),
.Y(n_1640)
);

BUFx6f_ASAP7_75t_L g1641 ( 
.A(n_1432),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1523),
.B(n_1343),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1437),
.B(n_1266),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1516),
.Y(n_1644)
);

NAND3xp33_ASAP7_75t_SL g1645 ( 
.A(n_1422),
.B(n_1257),
.C(n_1221),
.Y(n_1645)
);

NOR2x2_ASAP7_75t_L g1646 ( 
.A(n_1409),
.B(n_1379),
.Y(n_1646)
);

CKINVDCx20_ASAP7_75t_R g1647 ( 
.A(n_1431),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1575),
.B(n_1371),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1442),
.B(n_1381),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1542),
.B(n_1371),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1417),
.Y(n_1651)
);

BUFx4f_ASAP7_75t_L g1652 ( 
.A(n_1521),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1420),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1478),
.B(n_1237),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1425),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1444),
.B(n_1464),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1468),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1501),
.B(n_1237),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1471),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1474),
.B(n_1246),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1454),
.A2(n_1253),
.B1(n_1379),
.B2(n_1268),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_1521),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1556),
.B(n_1247),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1568),
.B(n_1327),
.Y(n_1664)
);

BUFx3_ASAP7_75t_L g1665 ( 
.A(n_1522),
.Y(n_1665)
);

BUFx2_ASAP7_75t_L g1666 ( 
.A(n_1522),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1457),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1519),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1426),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1522),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1430),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1462),
.B(n_1247),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1435),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1531),
.B(n_1535),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_SL g1675 ( 
.A(n_1483),
.B(n_1515),
.Y(n_1675)
);

INVxp67_ASAP7_75t_SL g1676 ( 
.A(n_1452),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_1550),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1505),
.Y(n_1678)
);

AOI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1458),
.A2(n_1253),
.B1(n_1379),
.B2(n_1268),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1526),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_SL g1681 ( 
.A(n_1440),
.B(n_1249),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1482),
.B(n_1253),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1486),
.B(n_1385),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1539),
.B(n_1386),
.Y(n_1684)
);

BUFx4f_ASAP7_75t_L g1685 ( 
.A(n_1432),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_SL g1686 ( 
.A(n_1445),
.B(n_1355),
.Y(n_1686)
);

INVx2_ASAP7_75t_SL g1687 ( 
.A(n_1579),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1428),
.B(n_1554),
.Y(n_1688)
);

NAND2xp33_ASAP7_75t_SL g1689 ( 
.A(n_1564),
.B(n_1400),
.Y(n_1689)
);

INVx1_ASAP7_75t_SL g1690 ( 
.A(n_1507),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1489),
.B(n_1386),
.Y(n_1691)
);

BUFx12f_ASAP7_75t_L g1692 ( 
.A(n_1579),
.Y(n_1692)
);

INVx1_ASAP7_75t_SL g1693 ( 
.A(n_1512),
.Y(n_1693)
);

AOI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1459),
.A2(n_1400),
.B1(n_1403),
.B2(n_1399),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_SL g1695 ( 
.A1(n_1547),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1514),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1573),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_SL g1698 ( 
.A(n_1441),
.B(n_917),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1496),
.B(n_1359),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1583),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1560),
.B(n_1359),
.Y(n_1701)
);

BUFx2_ASAP7_75t_L g1702 ( 
.A(n_1584),
.Y(n_1702)
);

INVx3_ASAP7_75t_L g1703 ( 
.A(n_1564),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1517),
.B(n_0),
.Y(n_1704)
);

AOI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1467),
.A2(n_917),
.B1(n_3),
.B2(n_1),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_1581),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1447),
.B(n_2),
.Y(n_1707)
);

INVxp67_ASAP7_75t_L g1708 ( 
.A(n_1536),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1532),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1585),
.Y(n_1710)
);

INVx3_ASAP7_75t_L g1711 ( 
.A(n_1452),
.Y(n_1711)
);

INVx3_ASAP7_75t_L g1712 ( 
.A(n_1599),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1450),
.B(n_3),
.Y(n_1713)
);

INVx2_ASAP7_75t_SL g1714 ( 
.A(n_1433),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1453),
.B(n_4),
.Y(n_1715)
);

INVx4_ASAP7_75t_L g1716 ( 
.A(n_1432),
.Y(n_1716)
);

CKINVDCx20_ASAP7_75t_R g1717 ( 
.A(n_1472),
.Y(n_1717)
);

OAI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1529),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_1718)
);

INVx3_ASAP7_75t_L g1719 ( 
.A(n_1599),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1558),
.B(n_5),
.Y(n_1720)
);

INVx3_ASAP7_75t_L g1721 ( 
.A(n_1599),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1565),
.B(n_7),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1571),
.B(n_7),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1543),
.B(n_8),
.Y(n_1724)
);

OR2x6_ASAP7_75t_L g1725 ( 
.A(n_1434),
.B(n_463),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1497),
.B(n_8),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1548),
.B(n_9),
.Y(n_1727)
);

INVx2_ASAP7_75t_SL g1728 ( 
.A(n_1584),
.Y(n_1728)
);

BUFx6f_ASAP7_75t_L g1729 ( 
.A(n_1423),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1494),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_SL g1731 ( 
.A(n_1513),
.B(n_9),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1562),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1461),
.B(n_10),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1415),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1481),
.B(n_11),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1494),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1456),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1545),
.B(n_12),
.Y(n_1738)
);

OR2x6_ASAP7_75t_L g1739 ( 
.A(n_1421),
.B(n_465),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1473),
.B(n_13),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1586),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_SL g1742 ( 
.A(n_1479),
.B(n_13),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1580),
.Y(n_1743)
);

AOI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1574),
.A2(n_1485),
.B1(n_1491),
.B2(n_1487),
.Y(n_1744)
);

OR2x6_ASAP7_75t_SL g1745 ( 
.A(n_1502),
.B(n_1593),
.Y(n_1745)
);

INVx2_ASAP7_75t_SL g1746 ( 
.A(n_1495),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1595),
.B(n_14),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1443),
.B(n_14),
.Y(n_1748)
);

BUFx8_ASAP7_75t_L g1749 ( 
.A(n_1418),
.Y(n_1749)
);

CKINVDCx8_ASAP7_75t_R g1750 ( 
.A(n_1492),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1580),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1582),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1544),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_SL g1754 ( 
.A(n_1538),
.B(n_15),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1597),
.B(n_16),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_SL g1756 ( 
.A(n_1494),
.B(n_16),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1582),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_SL g1758 ( 
.A(n_1494),
.B(n_17),
.Y(n_1758)
);

AOI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1509),
.A2(n_21),
.B1(n_17),
.B2(n_20),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1436),
.B(n_22),
.Y(n_1760)
);

BUFx6f_ASAP7_75t_SL g1761 ( 
.A(n_1591),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1449),
.B(n_22),
.Y(n_1762)
);

INVx8_ASAP7_75t_L g1763 ( 
.A(n_1511),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1589),
.Y(n_1764)
);

BUFx2_ASAP7_75t_L g1765 ( 
.A(n_1451),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1460),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1469),
.B(n_23),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1549),
.Y(n_1768)
);

BUFx6f_ASAP7_75t_L g1769 ( 
.A(n_1484),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1589),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1502),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_1771)
);

OAI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1569),
.A2(n_31),
.B1(n_27),
.B2(n_29),
.Y(n_1772)
);

NOR2x2_ASAP7_75t_L g1773 ( 
.A(n_1510),
.B(n_29),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1537),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1488),
.B(n_32),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1559),
.Y(n_1776)
);

BUFx3_ASAP7_75t_L g1777 ( 
.A(n_1592),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1534),
.B(n_33),
.Y(n_1778)
);

INVx5_ASAP7_75t_L g1779 ( 
.A(n_1572),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1561),
.Y(n_1780)
);

INVx2_ASAP7_75t_SL g1781 ( 
.A(n_1566),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1540),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_1782)
);

A2O1A1Ixp33_ASAP7_75t_L g1783 ( 
.A1(n_1619),
.A2(n_1463),
.B(n_1416),
.C(n_1557),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1678),
.B(n_1598),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1674),
.B(n_1587),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1612),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1601),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1690),
.B(n_1528),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_SL g1789 ( 
.A(n_1617),
.B(n_1577),
.Y(n_1789)
);

INVx2_ASAP7_75t_SL g1790 ( 
.A(n_1652),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1609),
.B(n_1576),
.Y(n_1791)
);

BUFx2_ASAP7_75t_L g1792 ( 
.A(n_1662),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1623),
.A2(n_1576),
.B(n_1476),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_L g1794 ( 
.A(n_1693),
.B(n_1608),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1688),
.B(n_1592),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1656),
.B(n_1567),
.Y(n_1796)
);

AOI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1684),
.A2(n_1476),
.B(n_1456),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_SL g1798 ( 
.A(n_1672),
.B(n_1577),
.Y(n_1798)
);

OAI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1602),
.A2(n_1552),
.B(n_1480),
.Y(n_1799)
);

CKINVDCx6p67_ASAP7_75t_R g1800 ( 
.A(n_1665),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1626),
.B(n_1590),
.Y(n_1801)
);

AOI21xp33_ASAP7_75t_L g1802 ( 
.A1(n_1699),
.A2(n_1480),
.B(n_1493),
.Y(n_1802)
);

AOI22x1_ASAP7_75t_L g1803 ( 
.A1(n_1636),
.A2(n_1527),
.B1(n_1546),
.B2(n_1530),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1616),
.Y(n_1804)
);

NAND2xp33_ASAP7_75t_SL g1805 ( 
.A(n_1633),
.B(n_1577),
.Y(n_1805)
);

OAI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1675),
.A2(n_1563),
.B(n_1570),
.Y(n_1806)
);

BUFx4f_ASAP7_75t_L g1807 ( 
.A(n_1606),
.Y(n_1807)
);

AOI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1600),
.A2(n_1577),
.B1(n_37),
.B2(n_34),
.Y(n_1808)
);

AND2x4_ASAP7_75t_L g1809 ( 
.A(n_1615),
.B(n_467),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1603),
.Y(n_1810)
);

O2A1O1Ixp33_ASAP7_75t_L g1811 ( 
.A1(n_1754),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1611),
.Y(n_1812)
);

NAND3xp33_ASAP7_75t_L g1813 ( 
.A(n_1782),
.B(n_38),
.C(n_39),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1605),
.B(n_39),
.Y(n_1814)
);

AOI22x1_ASAP7_75t_L g1815 ( 
.A1(n_1746),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_1815)
);

AOI33xp33_ASAP7_75t_L g1816 ( 
.A1(n_1771),
.A2(n_42),
.A3(n_44),
.B1(n_40),
.B2(n_41),
.B3(n_43),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1683),
.B(n_44),
.Y(n_1817)
);

AO32x1_ASAP7_75t_L g1818 ( 
.A1(n_1772),
.A2(n_47),
.A3(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_SL g1819 ( 
.A(n_1617),
.B(n_45),
.Y(n_1819)
);

INVxp67_ASAP7_75t_L g1820 ( 
.A(n_1634),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1624),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1734),
.B(n_46),
.Y(n_1822)
);

INVxp67_ASAP7_75t_SL g1823 ( 
.A(n_1777),
.Y(n_1823)
);

AOI21xp5_ASAP7_75t_L g1824 ( 
.A1(n_1689),
.A2(n_594),
.B(n_593),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1621),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1691),
.B(n_47),
.Y(n_1826)
);

OAI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1635),
.A2(n_48),
.B(n_49),
.Y(n_1827)
);

O2A1O1Ixp33_ASAP7_75t_L g1828 ( 
.A1(n_1718),
.A2(n_51),
.B(n_49),
.C(n_50),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1696),
.B(n_50),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_R g1830 ( 
.A(n_1667),
.B(n_469),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1649),
.A2(n_578),
.B(n_577),
.Y(n_1831)
);

NOR2x1_ASAP7_75t_L g1832 ( 
.A(n_1712),
.B(n_470),
.Y(n_1832)
);

O2A1O1Ixp33_ASAP7_75t_L g1833 ( 
.A1(n_1731),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1765),
.B(n_54),
.Y(n_1834)
);

INVx3_ASAP7_75t_L g1835 ( 
.A(n_1712),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1708),
.B(n_54),
.Y(n_1836)
);

AOI21x1_ASAP7_75t_L g1837 ( 
.A1(n_1701),
.A2(n_473),
.B(n_471),
.Y(n_1837)
);

O2A1O1Ixp33_ASAP7_75t_L g1838 ( 
.A1(n_1724),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_1838)
);

O2A1O1Ixp33_ASAP7_75t_SL g1839 ( 
.A1(n_1639),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_1839)
);

A2O1A1Ixp33_ASAP7_75t_L g1840 ( 
.A1(n_1707),
.A2(n_61),
.B(n_58),
.C(n_60),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1638),
.A2(n_597),
.B(n_478),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1625),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1615),
.B(n_60),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1726),
.B(n_61),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1657),
.Y(n_1845)
);

OAI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1630),
.A2(n_65),
.B1(n_62),
.B2(n_64),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1659),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_SL g1848 ( 
.A(n_1614),
.B(n_62),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_1706),
.B(n_477),
.Y(n_1849)
);

AOI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1698),
.A2(n_1681),
.B(n_1645),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1629),
.Y(n_1851)
);

CKINVDCx10_ASAP7_75t_R g1852 ( 
.A(n_1761),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1628),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1647),
.B(n_479),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1748),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1702),
.B(n_66),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1713),
.B(n_67),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1644),
.Y(n_1858)
);

OAI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1744),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1668),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1715),
.B(n_68),
.Y(n_1861)
);

NOR2xp33_ASAP7_75t_L g1862 ( 
.A(n_1750),
.B(n_481),
.Y(n_1862)
);

OAI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1663),
.A2(n_69),
.B(n_71),
.Y(n_1863)
);

OAI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1618),
.A2(n_483),
.B(n_482),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1775),
.B(n_71),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1687),
.B(n_72),
.Y(n_1866)
);

INVxp67_ASAP7_75t_L g1867 ( 
.A(n_1670),
.Y(n_1867)
);

OR2x6_ASAP7_75t_L g1868 ( 
.A(n_1725),
.B(n_485),
.Y(n_1868)
);

OAI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1714),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1651),
.Y(n_1870)
);

O2A1O1Ixp5_ASAP7_75t_L g1871 ( 
.A1(n_1756),
.A2(n_75),
.B(n_73),
.C(n_74),
.Y(n_1871)
);

OAI21x1_ASAP7_75t_L g1872 ( 
.A1(n_1730),
.A2(n_1736),
.B(n_1737),
.Y(n_1872)
);

OR2x6_ASAP7_75t_SL g1873 ( 
.A(n_1677),
.B(n_76),
.Y(n_1873)
);

O2A1O1Ixp5_ASAP7_75t_L g1874 ( 
.A1(n_1758),
.A2(n_79),
.B(n_77),
.C(n_78),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1664),
.B(n_77),
.Y(n_1875)
);

AOI21x1_ASAP7_75t_L g1876 ( 
.A1(n_1682),
.A2(n_487),
.B(n_486),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1727),
.B(n_78),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1728),
.B(n_1704),
.Y(n_1878)
);

BUFx8_ASAP7_75t_L g1879 ( 
.A(n_1761),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1648),
.B(n_79),
.Y(n_1880)
);

AO21x1_ASAP7_75t_L g1881 ( 
.A1(n_1722),
.A2(n_80),
.B(n_81),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_L g1882 ( 
.A(n_1643),
.B(n_488),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1723),
.B(n_80),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1658),
.B(n_81),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_L g1885 ( 
.A(n_1717),
.B(n_489),
.Y(n_1885)
);

OAI21xp5_ASAP7_75t_L g1886 ( 
.A1(n_1737),
.A2(n_493),
.B(n_490),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1680),
.Y(n_1887)
);

INVxp67_ASAP7_75t_L g1888 ( 
.A(n_1666),
.Y(n_1888)
);

AOI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1676),
.A2(n_495),
.B(n_494),
.Y(n_1889)
);

OAI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1743),
.A2(n_499),
.B(n_498),
.Y(n_1890)
);

NAND2xp33_ASAP7_75t_L g1891 ( 
.A(n_1729),
.B(n_82),
.Y(n_1891)
);

OAI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1739),
.A2(n_1622),
.B1(n_1695),
.B2(n_1745),
.Y(n_1892)
);

INVx1_ASAP7_75t_SL g1893 ( 
.A(n_1646),
.Y(n_1893)
);

NOR2x1_ASAP7_75t_L g1894 ( 
.A(n_1719),
.B(n_503),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1739),
.B(n_1740),
.Y(n_1895)
);

INVx1_ASAP7_75t_SL g1896 ( 
.A(n_1632),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1778),
.B(n_82),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1709),
.B(n_1753),
.Y(n_1898)
);

AO22x1_ASAP7_75t_L g1899 ( 
.A1(n_1749),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1653),
.Y(n_1900)
);

AOI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1751),
.A2(n_592),
.B(n_510),
.Y(n_1901)
);

BUFx4f_ASAP7_75t_L g1902 ( 
.A(n_1606),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1768),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1720),
.B(n_84),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1747),
.B(n_85),
.Y(n_1905)
);

INVxp67_ASAP7_75t_L g1906 ( 
.A(n_1613),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1752),
.A2(n_591),
.B(n_511),
.Y(n_1907)
);

AO21x1_ASAP7_75t_L g1908 ( 
.A1(n_1738),
.A2(n_86),
.B(n_87),
.Y(n_1908)
);

AOI21x1_ASAP7_75t_L g1909 ( 
.A1(n_1757),
.A2(n_512),
.B(n_509),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1755),
.B(n_86),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1776),
.B(n_87),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_SL g1912 ( 
.A(n_1729),
.B(n_88),
.Y(n_1912)
);

OAI22xp5_ASAP7_75t_L g1913 ( 
.A1(n_1661),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_SL g1914 ( 
.A(n_1729),
.B(n_90),
.Y(n_1914)
);

INVx3_ASAP7_75t_L g1915 ( 
.A(n_1719),
.Y(n_1915)
);

A2O1A1Ixp33_ASAP7_75t_L g1916 ( 
.A1(n_1733),
.A2(n_93),
.B(n_91),
.C(n_92),
.Y(n_1916)
);

AOI21xp5_ASAP7_75t_L g1917 ( 
.A1(n_1764),
.A2(n_515),
.B(n_514),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1770),
.B(n_91),
.Y(n_1918)
);

NAND2x1p5_ASAP7_75t_L g1919 ( 
.A(n_1721),
.B(n_517),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1655),
.Y(n_1920)
);

BUFx3_ASAP7_75t_L g1921 ( 
.A(n_1652),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1669),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1671),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1735),
.B(n_92),
.Y(n_1924)
);

NOR2xp33_ASAP7_75t_L g1925 ( 
.A(n_1610),
.B(n_523),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1763),
.B(n_93),
.Y(n_1926)
);

OAI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1705),
.A2(n_94),
.B(n_95),
.Y(n_1927)
);

HB1xp67_ASAP7_75t_L g1928 ( 
.A(n_1640),
.Y(n_1928)
);

AOI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1694),
.A2(n_588),
.B(n_525),
.Y(n_1929)
);

AOI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1711),
.A2(n_587),
.B(n_526),
.Y(n_1930)
);

BUFx3_ASAP7_75t_L g1931 ( 
.A(n_1607),
.Y(n_1931)
);

OAI21xp33_ASAP7_75t_L g1932 ( 
.A1(n_1766),
.A2(n_1774),
.B(n_1759),
.Y(n_1932)
);

AOI21xp5_ASAP7_75t_L g1933 ( 
.A1(n_1711),
.A2(n_585),
.B(n_527),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_SL g1934 ( 
.A(n_1769),
.B(n_94),
.Y(n_1934)
);

AOI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1620),
.A2(n_1660),
.B(n_1686),
.Y(n_1935)
);

AOI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1679),
.A2(n_1654),
.B(n_1725),
.Y(n_1936)
);

AOI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1703),
.A2(n_528),
.B(n_524),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1742),
.B(n_529),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1780),
.Y(n_1939)
);

AOI21xp5_ASAP7_75t_L g1940 ( 
.A1(n_1703),
.A2(n_584),
.B(n_530),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1763),
.B(n_1673),
.Y(n_1941)
);

INVx5_ASAP7_75t_L g1942 ( 
.A(n_1604),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1697),
.B(n_95),
.Y(n_1943)
);

OAI22x1_ASAP7_75t_L g1944 ( 
.A1(n_1815),
.A2(n_1732),
.B1(n_1710),
.B2(n_1700),
.Y(n_1944)
);

OAI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1813),
.A2(n_1762),
.B(n_1760),
.Y(n_1945)
);

OAI21x1_ASAP7_75t_SL g1946 ( 
.A1(n_1881),
.A2(n_1767),
.B(n_1741),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1853),
.Y(n_1947)
);

AND3x2_ASAP7_75t_L g1948 ( 
.A(n_1819),
.B(n_1642),
.C(n_1650),
.Y(n_1948)
);

A2O1A1Ixp33_ASAP7_75t_L g1949 ( 
.A1(n_1932),
.A2(n_1642),
.B(n_1631),
.C(n_1685),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1896),
.B(n_1781),
.Y(n_1950)
);

OAI21xp5_ASAP7_75t_L g1951 ( 
.A1(n_1813),
.A2(n_1685),
.B(n_1637),
.Y(n_1951)
);

AOI21xp5_ASAP7_75t_L g1952 ( 
.A1(n_1797),
.A2(n_1779),
.B(n_1769),
.Y(n_1952)
);

BUFx3_ASAP7_75t_L g1953 ( 
.A(n_1931),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_L g1954 ( 
.A(n_1794),
.B(n_1692),
.Y(n_1954)
);

NOR2xp67_ASAP7_75t_L g1955 ( 
.A(n_1906),
.B(n_1627),
.Y(n_1955)
);

A2O1A1Ixp33_ASAP7_75t_L g1956 ( 
.A1(n_1927),
.A2(n_1650),
.B(n_1779),
.C(n_1769),
.Y(n_1956)
);

NAND2x1p5_ASAP7_75t_L g1957 ( 
.A(n_1942),
.B(n_1779),
.Y(n_1957)
);

NAND2xp33_ASAP7_75t_L g1958 ( 
.A(n_1895),
.B(n_1892),
.Y(n_1958)
);

AOI21xp5_ASAP7_75t_L g1959 ( 
.A1(n_1793),
.A2(n_1864),
.B(n_1850),
.Y(n_1959)
);

BUFx6f_ASAP7_75t_L g1960 ( 
.A(n_1921),
.Y(n_1960)
);

BUFx3_ASAP7_75t_L g1961 ( 
.A(n_1792),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1870),
.Y(n_1962)
);

OAI21x1_ASAP7_75t_L g1963 ( 
.A1(n_1799),
.A2(n_1637),
.B(n_1604),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1896),
.B(n_1749),
.Y(n_1964)
);

OAI21x1_ASAP7_75t_L g1965 ( 
.A1(n_1799),
.A2(n_1637),
.B(n_1604),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1796),
.B(n_1791),
.Y(n_1966)
);

OA21x2_ASAP7_75t_L g1967 ( 
.A1(n_1802),
.A2(n_1637),
.B(n_1604),
.Y(n_1967)
);

OR2x2_ASAP7_75t_L g1968 ( 
.A(n_1875),
.B(n_1641),
.Y(n_1968)
);

OAI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1783),
.A2(n_1848),
.B(n_1864),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1872),
.Y(n_1970)
);

O2A1O1Ixp5_ASAP7_75t_L g1971 ( 
.A1(n_1827),
.A2(n_1863),
.B(n_1846),
.C(n_1859),
.Y(n_1971)
);

A2O1A1Ixp33_ASAP7_75t_L g1972 ( 
.A1(n_1828),
.A2(n_1641),
.B(n_1773),
.C(n_99),
.Y(n_1972)
);

OAI21x1_ASAP7_75t_L g1973 ( 
.A1(n_1837),
.A2(n_1876),
.B(n_1909),
.Y(n_1973)
);

AND2x6_ASAP7_75t_L g1974 ( 
.A(n_1809),
.B(n_1641),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1900),
.Y(n_1975)
);

INVx3_ASAP7_75t_L g1976 ( 
.A(n_1942),
.Y(n_1976)
);

OR2x2_ASAP7_75t_L g1977 ( 
.A(n_1823),
.B(n_1716),
.Y(n_1977)
);

NAND2x1p5_ASAP7_75t_L g1978 ( 
.A(n_1942),
.B(n_1716),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1865),
.B(n_532),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1795),
.B(n_96),
.Y(n_1980)
);

BUFx2_ASAP7_75t_L g1981 ( 
.A(n_1820),
.Y(n_1981)
);

AOI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1789),
.A2(n_536),
.B(n_534),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1920),
.Y(n_1983)
);

A2O1A1Ixp33_ASAP7_75t_L g1984 ( 
.A1(n_1838),
.A2(n_100),
.B(n_97),
.C(n_99),
.Y(n_1984)
);

A2O1A1Ixp33_ASAP7_75t_L g1985 ( 
.A1(n_1811),
.A2(n_102),
.B(n_100),
.C(n_101),
.Y(n_1985)
);

OAI21xp5_ASAP7_75t_L g1986 ( 
.A1(n_1806),
.A2(n_102),
.B(n_103),
.Y(n_1986)
);

A2O1A1Ixp33_ASAP7_75t_L g1987 ( 
.A1(n_1938),
.A2(n_106),
.B(n_104),
.C(n_105),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1817),
.B(n_104),
.Y(n_1988)
);

AOI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1789),
.A2(n_538),
.B(n_537),
.Y(n_1989)
);

OAI21xp5_ASAP7_75t_L g1990 ( 
.A1(n_1841),
.A2(n_105),
.B(n_106),
.Y(n_1990)
);

AOI21x1_ASAP7_75t_L g1991 ( 
.A1(n_1936),
.A2(n_544),
.B(n_542),
.Y(n_1991)
);

NOR2xp33_ASAP7_75t_L g1992 ( 
.A(n_1893),
.B(n_546),
.Y(n_1992)
);

AND2x4_ASAP7_75t_L g1993 ( 
.A(n_1809),
.B(n_547),
.Y(n_1993)
);

BUFx6f_ASAP7_75t_L g1994 ( 
.A(n_1807),
.Y(n_1994)
);

BUFx4_ASAP7_75t_SL g1995 ( 
.A(n_1868),
.Y(n_1995)
);

INVx4_ASAP7_75t_L g1996 ( 
.A(n_1807),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1826),
.B(n_107),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1814),
.B(n_107),
.Y(n_1998)
);

OAI22x1_ASAP7_75t_L g1999 ( 
.A1(n_1803),
.A2(n_1808),
.B1(n_1893),
.B2(n_1912),
.Y(n_1999)
);

AOI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1868),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_2000)
);

NAND3xp33_ASAP7_75t_L g2001 ( 
.A(n_1840),
.B(n_108),
.C(n_109),
.Y(n_2001)
);

AOI21x1_ASAP7_75t_SL g2002 ( 
.A1(n_1926),
.A2(n_111),
.B(n_112),
.Y(n_2002)
);

OAI21xp5_ASAP7_75t_L g2003 ( 
.A1(n_1788),
.A2(n_111),
.B(n_113),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1898),
.B(n_113),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1816),
.B(n_114),
.Y(n_2005)
);

A2O1A1Ixp33_ASAP7_75t_L g2006 ( 
.A1(n_1833),
.A2(n_116),
.B(n_114),
.C(n_115),
.Y(n_2006)
);

INVx2_ASAP7_75t_SL g2007 ( 
.A(n_1902),
.Y(n_2007)
);

OAI21xp5_ASAP7_75t_L g2008 ( 
.A1(n_1935),
.A2(n_1890),
.B(n_1831),
.Y(n_2008)
);

NAND3xp33_ASAP7_75t_L g2009 ( 
.A(n_1916),
.B(n_116),
.C(n_117),
.Y(n_2009)
);

OAI21xp5_ASAP7_75t_L g2010 ( 
.A1(n_1890),
.A2(n_118),
.B(n_119),
.Y(n_2010)
);

AOI21xp5_ASAP7_75t_L g2011 ( 
.A1(n_1886),
.A2(n_552),
.B(n_550),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_L g2012 ( 
.A(n_1785),
.B(n_553),
.Y(n_2012)
);

AOI21xp5_ASAP7_75t_L g2013 ( 
.A1(n_1886),
.A2(n_555),
.B(n_554),
.Y(n_2013)
);

INVx2_ASAP7_75t_SL g2014 ( 
.A(n_1902),
.Y(n_2014)
);

INVx4_ASAP7_75t_L g2015 ( 
.A(n_1800),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1922),
.Y(n_2016)
);

AOI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_1798),
.A2(n_1805),
.B(n_1824),
.Y(n_2017)
);

BUFx2_ASAP7_75t_L g2018 ( 
.A(n_1888),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1897),
.B(n_118),
.Y(n_2019)
);

NOR2x1_ASAP7_75t_SL g2020 ( 
.A(n_1868),
.B(n_556),
.Y(n_2020)
);

AOI21xp5_ASAP7_75t_L g2021 ( 
.A1(n_1929),
.A2(n_558),
.B(n_557),
.Y(n_2021)
);

AO31x2_ASAP7_75t_L g2022 ( 
.A1(n_1913),
.A2(n_561),
.A3(n_562),
.B(n_559),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1923),
.Y(n_2023)
);

INVx6_ASAP7_75t_SL g2024 ( 
.A(n_1852),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_SL g2025 ( 
.A(n_1941),
.B(n_567),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1878),
.B(n_119),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1918),
.B(n_120),
.Y(n_2027)
);

NAND3xp33_ASAP7_75t_SL g2028 ( 
.A(n_1819),
.B(n_120),
.C(n_121),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1786),
.Y(n_2029)
);

OAI22x1_ASAP7_75t_L g2030 ( 
.A1(n_1914),
.A2(n_1877),
.B1(n_1787),
.B2(n_1812),
.Y(n_2030)
);

BUFx3_ASAP7_75t_L g2031 ( 
.A(n_1879),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1880),
.B(n_568),
.Y(n_2032)
);

BUFx4f_ASAP7_75t_SL g2033 ( 
.A(n_1879),
.Y(n_2033)
);

INVx5_ASAP7_75t_L g2034 ( 
.A(n_1835),
.Y(n_2034)
);

OA22x2_ASAP7_75t_L g2035 ( 
.A1(n_1843),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1804),
.B(n_122),
.Y(n_2036)
);

AND3x4_ASAP7_75t_L g2037 ( 
.A(n_1873),
.B(n_124),
.C(n_125),
.Y(n_2037)
);

AOI21xp33_ASAP7_75t_L g2038 ( 
.A1(n_1844),
.A2(n_124),
.B(n_125),
.Y(n_2038)
);

INVx3_ASAP7_75t_L g2039 ( 
.A(n_1835),
.Y(n_2039)
);

INVx1_ASAP7_75t_SL g2040 ( 
.A(n_1801),
.Y(n_2040)
);

OAI21x1_ASAP7_75t_SL g2041 ( 
.A1(n_1908),
.A2(n_126),
.B(n_127),
.Y(n_2041)
);

BUFx3_ASAP7_75t_L g2042 ( 
.A(n_1790),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1825),
.B(n_126),
.Y(n_2043)
);

A2O1A1Ixp33_ASAP7_75t_L g2044 ( 
.A1(n_1857),
.A2(n_129),
.B(n_127),
.C(n_128),
.Y(n_2044)
);

A2O1A1Ixp33_ASAP7_75t_L g2045 ( 
.A1(n_1861),
.A2(n_131),
.B(n_129),
.C(n_130),
.Y(n_2045)
);

O2A1O1Ixp5_ASAP7_75t_L g2046 ( 
.A1(n_1871),
.A2(n_133),
.B(n_130),
.C(n_132),
.Y(n_2046)
);

AOI22xp33_ASAP7_75t_L g2047 ( 
.A1(n_1891),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1851),
.B(n_134),
.Y(n_2048)
);

OR2x6_ASAP7_75t_L g2049 ( 
.A(n_1959),
.B(n_1919),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1966),
.B(n_2040),
.Y(n_2050)
);

BUFx3_ASAP7_75t_L g2051 ( 
.A(n_1961),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1947),
.Y(n_2052)
);

BUFx2_ASAP7_75t_L g2053 ( 
.A(n_1964),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1962),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1975),
.B(n_1810),
.Y(n_2055)
);

BUFx2_ASAP7_75t_L g2056 ( 
.A(n_1970),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1983),
.Y(n_2057)
);

AO21x1_ASAP7_75t_L g2058 ( 
.A1(n_2010),
.A2(n_1869),
.B(n_1883),
.Y(n_2058)
);

NAND2x1p5_ASAP7_75t_L g2059 ( 
.A(n_1963),
.B(n_1832),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2016),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_2023),
.B(n_1821),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1950),
.B(n_1842),
.Y(n_2062)
);

BUFx3_ASAP7_75t_L g2063 ( 
.A(n_1953),
.Y(n_2063)
);

BUFx2_ASAP7_75t_SL g2064 ( 
.A(n_1955),
.Y(n_2064)
);

BUFx3_ASAP7_75t_L g2065 ( 
.A(n_1957),
.Y(n_2065)
);

INVx5_ASAP7_75t_L g2066 ( 
.A(n_1976),
.Y(n_2066)
);

BUFx6f_ASAP7_75t_L g2067 ( 
.A(n_1994),
.Y(n_2067)
);

NAND2x1p5_ASAP7_75t_L g2068 ( 
.A(n_1965),
.B(n_1894),
.Y(n_2068)
);

NAND2x1p5_ASAP7_75t_L g2069 ( 
.A(n_1967),
.B(n_1915),
.Y(n_2069)
);

BUFx6f_ASAP7_75t_L g2070 ( 
.A(n_1994),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2029),
.Y(n_2071)
);

BUFx6f_ASAP7_75t_L g2072 ( 
.A(n_1994),
.Y(n_2072)
);

BUFx2_ASAP7_75t_L g2073 ( 
.A(n_1981),
.Y(n_2073)
);

AO21x1_ASAP7_75t_L g2074 ( 
.A1(n_1969),
.A2(n_1905),
.B(n_1904),
.Y(n_2074)
);

BUFx3_ASAP7_75t_L g2075 ( 
.A(n_2034),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2030),
.Y(n_2076)
);

BUFx3_ASAP7_75t_L g2077 ( 
.A(n_2034),
.Y(n_2077)
);

INVxp67_ASAP7_75t_SL g2078 ( 
.A(n_1952),
.Y(n_2078)
);

BUFx3_ASAP7_75t_L g2079 ( 
.A(n_2034),
.Y(n_2079)
);

BUFx2_ASAP7_75t_L g2080 ( 
.A(n_2018),
.Y(n_2080)
);

BUFx12f_ASAP7_75t_L g2081 ( 
.A(n_1996),
.Y(n_2081)
);

INVx6_ASAP7_75t_L g2082 ( 
.A(n_1996),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1980),
.B(n_1845),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2036),
.Y(n_2084)
);

INVx4_ASAP7_75t_L g2085 ( 
.A(n_1976),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1967),
.Y(n_2086)
);

INVxp67_ASAP7_75t_SL g2087 ( 
.A(n_2039),
.Y(n_2087)
);

BUFx2_ASAP7_75t_L g2088 ( 
.A(n_1968),
.Y(n_2088)
);

NOR2xp33_ASAP7_75t_L g2089 ( 
.A(n_2012),
.B(n_1910),
.Y(n_2089)
);

INVxp67_ASAP7_75t_SL g2090 ( 
.A(n_2039),
.Y(n_2090)
);

INVx2_ASAP7_75t_SL g2091 ( 
.A(n_1977),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1973),
.Y(n_2092)
);

CKINVDCx5p33_ASAP7_75t_R g2093 ( 
.A(n_2024),
.Y(n_2093)
);

INVx3_ASAP7_75t_L g2094 ( 
.A(n_1991),
.Y(n_2094)
);

INVx4_ASAP7_75t_L g2095 ( 
.A(n_1948),
.Y(n_2095)
);

BUFx3_ASAP7_75t_L g2096 ( 
.A(n_1960),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_2008),
.B(n_1847),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2043),
.Y(n_2098)
);

BUFx3_ASAP7_75t_L g2099 ( 
.A(n_1960),
.Y(n_2099)
);

BUFx2_ASAP7_75t_R g2100 ( 
.A(n_2031),
.Y(n_2100)
);

INVx4_ASAP7_75t_L g2101 ( 
.A(n_1974),
.Y(n_2101)
);

AOI22xp33_ASAP7_75t_L g2102 ( 
.A1(n_2003),
.A2(n_1855),
.B1(n_1924),
.B2(n_1925),
.Y(n_2102)
);

AND2x4_ASAP7_75t_L g2103 ( 
.A(n_2020),
.B(n_1915),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2004),
.B(n_1884),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_1958),
.B(n_1911),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1998),
.B(n_1784),
.Y(n_2106)
);

INVx6_ASAP7_75t_SL g2107 ( 
.A(n_1993),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2048),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1946),
.Y(n_2109)
);

AOI22xp33_ASAP7_75t_L g2110 ( 
.A1(n_1986),
.A2(n_1882),
.B1(n_1836),
.B2(n_1829),
.Y(n_2110)
);

BUFx3_ASAP7_75t_L g2111 ( 
.A(n_1960),
.Y(n_2111)
);

BUFx3_ASAP7_75t_L g2112 ( 
.A(n_2042),
.Y(n_2112)
);

NAND2x1p5_ASAP7_75t_L g2113 ( 
.A(n_2017),
.B(n_1934),
.Y(n_2113)
);

BUFx3_ASAP7_75t_L g2114 ( 
.A(n_1974),
.Y(n_2114)
);

INVx1_ASAP7_75t_SL g2115 ( 
.A(n_1954),
.Y(n_2115)
);

AOI22xp33_ASAP7_75t_L g2116 ( 
.A1(n_2001),
.A2(n_1885),
.B1(n_1854),
.B2(n_1849),
.Y(n_2116)
);

BUFx6f_ASAP7_75t_L g2117 ( 
.A(n_1974),
.Y(n_2117)
);

OAI21xp33_ASAP7_75t_L g2118 ( 
.A1(n_1987),
.A2(n_1943),
.B(n_1862),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2052),
.Y(n_2119)
);

HB1xp67_ASAP7_75t_L g2120 ( 
.A(n_2091),
.Y(n_2120)
);

OAI21xp5_ASAP7_75t_L g2121 ( 
.A1(n_2110),
.A2(n_1990),
.B(n_1971),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2097),
.B(n_2022),
.Y(n_2122)
);

CKINVDCx5p33_ASAP7_75t_R g2123 ( 
.A(n_2093),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2097),
.B(n_1988),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_2052),
.Y(n_2125)
);

OAI21xp5_ASAP7_75t_L g2126 ( 
.A1(n_2110),
.A2(n_2013),
.B(n_2011),
.Y(n_2126)
);

INVx3_ASAP7_75t_L g2127 ( 
.A(n_2103),
.Y(n_2127)
);

CKINVDCx16_ASAP7_75t_R g2128 ( 
.A(n_2063),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_2091),
.B(n_1997),
.Y(n_2129)
);

OAI22xp33_ASAP7_75t_L g2130 ( 
.A1(n_2095),
.A2(n_2000),
.B1(n_2009),
.B2(n_2028),
.Y(n_2130)
);

INVx8_ASAP7_75t_L g2131 ( 
.A(n_2081),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2054),
.Y(n_2132)
);

BUFx6f_ASAP7_75t_L g2133 ( 
.A(n_2117),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2057),
.Y(n_2134)
);

INVx3_ASAP7_75t_L g2135 ( 
.A(n_2103),
.Y(n_2135)
);

AO21x2_ASAP7_75t_L g2136 ( 
.A1(n_2092),
.A2(n_1984),
.B(n_2041),
.Y(n_2136)
);

BUFx3_ASAP7_75t_L g2137 ( 
.A(n_2081),
.Y(n_2137)
);

AO31x2_ASAP7_75t_L g2138 ( 
.A1(n_2086),
.A2(n_1944),
.A3(n_2020),
.B(n_1985),
.Y(n_2138)
);

BUFx12f_ASAP7_75t_L g2139 ( 
.A(n_2093),
.Y(n_2139)
);

AO22x1_ASAP7_75t_L g2140 ( 
.A1(n_2095),
.A2(n_2037),
.B1(n_2015),
.B2(n_1951),
.Y(n_2140)
);

BUFx2_ASAP7_75t_L g2141 ( 
.A(n_2076),
.Y(n_2141)
);

AOI22xp33_ASAP7_75t_L g2142 ( 
.A1(n_2058),
.A2(n_2047),
.B1(n_1999),
.B2(n_2038),
.Y(n_2142)
);

AOI222xp33_ASAP7_75t_L g2143 ( 
.A1(n_2102),
.A2(n_1972),
.B1(n_2005),
.B2(n_1945),
.C1(n_2045),
.C2(n_2044),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_2060),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2086),
.B(n_2056),
.Y(n_2145)
);

BUFx12f_ASAP7_75t_L g2146 ( 
.A(n_2067),
.Y(n_2146)
);

AOI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_2058),
.A2(n_1974),
.B1(n_1993),
.B2(n_1992),
.Y(n_2147)
);

AND2x6_ASAP7_75t_L g2148 ( 
.A(n_2117),
.B(n_1995),
.Y(n_2148)
);

OAI21x1_ASAP7_75t_L g2149 ( 
.A1(n_2094),
.A2(n_2021),
.B(n_2002),
.Y(n_2149)
);

AOI22xp33_ASAP7_75t_L g2150 ( 
.A1(n_2118),
.A2(n_2035),
.B1(n_2025),
.B2(n_2032),
.Y(n_2150)
);

OA21x2_ASAP7_75t_L g2151 ( 
.A1(n_2092),
.A2(n_2109),
.B(n_2056),
.Y(n_2151)
);

OAI21x1_ASAP7_75t_L g2152 ( 
.A1(n_2094),
.A2(n_2068),
.B(n_2059),
.Y(n_2152)
);

OAI21x1_ASAP7_75t_L g2153 ( 
.A1(n_2094),
.A2(n_1989),
.B(n_1982),
.Y(n_2153)
);

NOR2xp33_ASAP7_75t_L g2154 ( 
.A(n_2115),
.B(n_2015),
.Y(n_2154)
);

AOI21xp33_ASAP7_75t_L g2155 ( 
.A1(n_2078),
.A2(n_2027),
.B(n_2026),
.Y(n_2155)
);

OAI21x1_ASAP7_75t_L g2156 ( 
.A1(n_2059),
.A2(n_1889),
.B(n_1930),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2125),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2125),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2134),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2134),
.Y(n_2160)
);

AOI22xp33_ASAP7_75t_L g2161 ( 
.A1(n_2121),
.A2(n_2074),
.B1(n_2102),
.B2(n_2049),
.Y(n_2161)
);

INVx2_ASAP7_75t_SL g2162 ( 
.A(n_2127),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2144),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_2145),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2144),
.Y(n_2165)
);

BUFx6f_ASAP7_75t_L g2166 ( 
.A(n_2148),
.Y(n_2166)
);

CKINVDCx11_ASAP7_75t_R g2167 ( 
.A(n_2139),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2119),
.Y(n_2168)
);

HB1xp67_ASAP7_75t_L g2169 ( 
.A(n_2120),
.Y(n_2169)
);

BUFx2_ASAP7_75t_L g2170 ( 
.A(n_2127),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_2145),
.Y(n_2171)
);

AOI22xp33_ASAP7_75t_SL g2172 ( 
.A1(n_2126),
.A2(n_2089),
.B1(n_2095),
.B2(n_2113),
.Y(n_2172)
);

AOI22xp33_ASAP7_75t_SL g2173 ( 
.A1(n_2122),
.A2(n_2089),
.B1(n_2113),
.B2(n_2049),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_2151),
.Y(n_2174)
);

INVx1_ASAP7_75t_SL g2175 ( 
.A(n_2128),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_2151),
.Y(n_2176)
);

BUFx3_ASAP7_75t_L g2177 ( 
.A(n_2139),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2132),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_2174),
.Y(n_2179)
);

OR2x2_ASAP7_75t_L g2180 ( 
.A(n_2164),
.B(n_2141),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_2174),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2159),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_2176),
.Y(n_2183)
);

HB1xp67_ASAP7_75t_L g2184 ( 
.A(n_2169),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2178),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2178),
.Y(n_2186)
);

OAI21xp33_ASAP7_75t_SL g2187 ( 
.A1(n_2161),
.A2(n_2152),
.B(n_2122),
.Y(n_2187)
);

HB1xp67_ASAP7_75t_L g2188 ( 
.A(n_2168),
.Y(n_2188)
);

OAI21x1_ASAP7_75t_L g2189 ( 
.A1(n_2176),
.A2(n_2152),
.B(n_2151),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_2184),
.B(n_2175),
.Y(n_2190)
);

OR2x6_ASAP7_75t_L g2191 ( 
.A(n_2189),
.B(n_2166),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_2180),
.B(n_2127),
.Y(n_2192)
);

OR2x6_ASAP7_75t_L g2193 ( 
.A(n_2189),
.B(n_2166),
.Y(n_2193)
);

NAND2xp33_ASAP7_75t_R g2194 ( 
.A(n_2185),
.B(n_2123),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2186),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_2180),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2188),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_2196),
.B(n_2170),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2192),
.B(n_2170),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2191),
.B(n_2187),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_2191),
.B(n_2177),
.Y(n_2201)
);

BUFx2_ASAP7_75t_L g2202 ( 
.A(n_2190),
.Y(n_2202)
);

HB1xp67_ASAP7_75t_L g2203 ( 
.A(n_2197),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2195),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2191),
.Y(n_2205)
);

OR2x2_ASAP7_75t_L g2206 ( 
.A(n_2193),
.B(n_2141),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2193),
.Y(n_2207)
);

AND2x4_ASAP7_75t_L g2208 ( 
.A(n_2202),
.B(n_2193),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2203),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2205),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2201),
.B(n_2177),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2204),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2205),
.Y(n_2213)
);

AND2x4_ASAP7_75t_L g2214 ( 
.A(n_2201),
.B(n_2166),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2207),
.Y(n_2215)
);

INVxp67_ASAP7_75t_L g2216 ( 
.A(n_2198),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_2198),
.B(n_2167),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2206),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2210),
.Y(n_2219)
);

OR2x2_ASAP7_75t_L g2220 ( 
.A(n_2216),
.B(n_2200),
.Y(n_2220)
);

OAI21x1_ASAP7_75t_L g2221 ( 
.A1(n_2210),
.A2(n_2200),
.B(n_2199),
.Y(n_2221)
);

AOI21xp33_ASAP7_75t_L g2222 ( 
.A1(n_2218),
.A2(n_2194),
.B(n_2172),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_2208),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2213),
.Y(n_2224)
);

AOI21x1_ASAP7_75t_L g2225 ( 
.A1(n_2213),
.A2(n_2199),
.B(n_2140),
.Y(n_2225)
);

AOI21xp5_ASAP7_75t_L g2226 ( 
.A1(n_2209),
.A2(n_2130),
.B(n_1899),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_2217),
.B(n_2123),
.Y(n_2227)
);

INVx4_ASAP7_75t_L g2228 ( 
.A(n_2223),
.Y(n_2228)
);

AOI211xp5_ASAP7_75t_L g2229 ( 
.A1(n_2222),
.A2(n_2215),
.B(n_2211),
.C(n_2216),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_2223),
.B(n_2212),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_2227),
.B(n_2214),
.Y(n_2231)
);

AO21x2_ASAP7_75t_L g2232 ( 
.A1(n_2230),
.A2(n_2224),
.B(n_2219),
.Y(n_2232)
);

OR2x2_ASAP7_75t_L g2233 ( 
.A(n_2228),
.B(n_2220),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_2231),
.B(n_2214),
.Y(n_2234)
);

INVx2_ASAP7_75t_SL g2235 ( 
.A(n_2229),
.Y(n_2235)
);

NAND2x1p5_ASAP7_75t_L g2236 ( 
.A(n_2233),
.B(n_2214),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_2234),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2235),
.B(n_2226),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2232),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2232),
.Y(n_2240)
);

OR2x2_ASAP7_75t_L g2241 ( 
.A(n_2233),
.B(n_2221),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2239),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2239),
.Y(n_2243)
);

AND2x4_ASAP7_75t_L g2244 ( 
.A(n_2237),
.B(n_2208),
.Y(n_2244)
);

OAI22xp5_ASAP7_75t_L g2245 ( 
.A1(n_2236),
.A2(n_2226),
.B1(n_2208),
.B2(n_2225),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2241),
.B(n_2221),
.Y(n_2246)
);

NAND3xp33_ASAP7_75t_SL g2247 ( 
.A(n_2240),
.B(n_1830),
.C(n_2024),
.Y(n_2247)
);

INVx2_ASAP7_75t_SL g2248 ( 
.A(n_2238),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_2237),
.B(n_2154),
.Y(n_2249)
);

NOR3xp33_ASAP7_75t_L g2250 ( 
.A(n_2238),
.B(n_2019),
.C(n_2106),
.Y(n_2250)
);

OAI22xp5_ASAP7_75t_L g2251 ( 
.A1(n_2236),
.A2(n_2166),
.B1(n_2100),
.B2(n_2194),
.Y(n_2251)
);

CKINVDCx14_ASAP7_75t_R g2252 ( 
.A(n_2247),
.Y(n_2252)
);

CKINVDCx16_ASAP7_75t_R g2253 ( 
.A(n_2244),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_2249),
.B(n_2137),
.Y(n_2254)
);

OR2x2_ASAP7_75t_L g2255 ( 
.A(n_2246),
.B(n_2073),
.Y(n_2255)
);

INVx2_ASAP7_75t_SL g2256 ( 
.A(n_2245),
.Y(n_2256)
);

INVx1_ASAP7_75t_SL g2257 ( 
.A(n_2248),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_2250),
.B(n_2137),
.Y(n_2258)
);

AOI22xp33_ASAP7_75t_L g2259 ( 
.A1(n_2251),
.A2(n_2166),
.B1(n_2074),
.B2(n_2148),
.Y(n_2259)
);

AND2x4_ASAP7_75t_L g2260 ( 
.A(n_2242),
.B(n_2063),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2243),
.B(n_2080),
.Y(n_2261)
);

HB1xp67_ASAP7_75t_L g2262 ( 
.A(n_2244),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_2244),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2244),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2253),
.B(n_2179),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2262),
.B(n_2053),
.Y(n_2266)
);

NOR3xp33_ASAP7_75t_L g2267 ( 
.A(n_2252),
.B(n_2033),
.C(n_1856),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2262),
.Y(n_2268)
);

A2O1A1Ixp33_ASAP7_75t_SL g2269 ( 
.A1(n_2263),
.A2(n_137),
.B(n_135),
.C(n_136),
.Y(n_2269)
);

OAI221xp5_ASAP7_75t_L g2270 ( 
.A1(n_2256),
.A2(n_2064),
.B1(n_2142),
.B2(n_2116),
.C(n_2006),
.Y(n_2270)
);

AOI222xp33_ASAP7_75t_L g2271 ( 
.A1(n_2264),
.A2(n_2116),
.B1(n_2150),
.B2(n_2108),
.C1(n_2098),
.C2(n_2084),
.Y(n_2271)
);

INVxp67_ASAP7_75t_SL g2272 ( 
.A(n_2260),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_2254),
.B(n_2258),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2261),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_2257),
.B(n_2051),
.Y(n_2275)
);

OAI221xp5_ASAP7_75t_L g2276 ( 
.A1(n_2259),
.A2(n_2257),
.B1(n_2255),
.B2(n_2260),
.C(n_2155),
.Y(n_2276)
);

AOI21xp33_ASAP7_75t_SL g2277 ( 
.A1(n_2253),
.A2(n_2014),
.B(n_2007),
.Y(n_2277)
);

AOI211xp5_ASAP7_75t_L g2278 ( 
.A1(n_2262),
.A2(n_1834),
.B(n_2104),
.C(n_1822),
.Y(n_2278)
);

INVx1_ASAP7_75t_SL g2279 ( 
.A(n_2262),
.Y(n_2279)
);

OAI32xp33_ASAP7_75t_L g2280 ( 
.A1(n_2279),
.A2(n_2181),
.A3(n_2183),
.B1(n_2179),
.B2(n_2112),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_2279),
.B(n_2268),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2266),
.Y(n_2282)
);

OAI221xp5_ASAP7_75t_L g2283 ( 
.A1(n_2267),
.A2(n_2147),
.B1(n_2173),
.B2(n_2051),
.C(n_2112),
.Y(n_2283)
);

BUFx2_ASAP7_75t_L g2284 ( 
.A(n_2272),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2275),
.Y(n_2285)
);

OAI221xp5_ASAP7_75t_L g2286 ( 
.A1(n_2276),
.A2(n_2143),
.B1(n_2082),
.B2(n_2129),
.C(n_1867),
.Y(n_2286)
);

AOI21xp33_ASAP7_75t_L g2287 ( 
.A1(n_2274),
.A2(n_2131),
.B(n_1979),
.Y(n_2287)
);

OAI22xp5_ASAP7_75t_L g2288 ( 
.A1(n_2265),
.A2(n_2183),
.B1(n_2181),
.B2(n_2131),
.Y(n_2288)
);

HB1xp67_ASAP7_75t_L g2289 ( 
.A(n_2273),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2278),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2277),
.Y(n_2291)
);

OAI22xp33_ASAP7_75t_SL g2292 ( 
.A1(n_2270),
.A2(n_2082),
.B1(n_2182),
.B2(n_2099),
.Y(n_2292)
);

AOI22xp5_ASAP7_75t_L g2293 ( 
.A1(n_2271),
.A2(n_2131),
.B1(n_2148),
.B2(n_2082),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_SL g2294 ( 
.A(n_2284),
.B(n_2269),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2289),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2282),
.B(n_2281),
.Y(n_2296)
);

NAND2xp33_ASAP7_75t_L g2297 ( 
.A(n_2285),
.B(n_2291),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2290),
.B(n_2182),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_SL g2299 ( 
.A(n_2292),
.B(n_2067),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2287),
.B(n_2124),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2286),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2280),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2293),
.Y(n_2303)
);

NOR2x1p5_ASAP7_75t_L g2304 ( 
.A(n_2283),
.B(n_2096),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_L g2305 ( 
.A(n_2288),
.B(n_2131),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2284),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2284),
.Y(n_2307)
);

INVx1_ASAP7_75t_SL g2308 ( 
.A(n_2284),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_2284),
.B(n_2083),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2284),
.B(n_1928),
.Y(n_2310)
);

INVx1_ASAP7_75t_SL g2311 ( 
.A(n_2284),
.Y(n_2311)
);

INVxp67_ASAP7_75t_L g2312 ( 
.A(n_2284),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2284),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_2289),
.B(n_2162),
.Y(n_2314)
);

INVx1_ASAP7_75t_SL g2315 ( 
.A(n_2284),
.Y(n_2315)
);

NOR3x1_ASAP7_75t_L g2316 ( 
.A(n_2294),
.B(n_135),
.C(n_136),
.Y(n_2316)
);

NAND3xp33_ASAP7_75t_L g2317 ( 
.A(n_2297),
.B(n_1866),
.C(n_2067),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2314),
.Y(n_2318)
);

AOI211xp5_ASAP7_75t_L g2319 ( 
.A1(n_2315),
.A2(n_1839),
.B(n_2070),
.C(n_2067),
.Y(n_2319)
);

AOI211xp5_ASAP7_75t_L g2320 ( 
.A1(n_2315),
.A2(n_2072),
.B(n_2070),
.C(n_140),
.Y(n_2320)
);

NAND4xp25_ASAP7_75t_L g2321 ( 
.A(n_2296),
.B(n_2096),
.C(n_2111),
.D(n_2099),
.Y(n_2321)
);

NAND4xp25_ASAP7_75t_L g2322 ( 
.A(n_2305),
.B(n_2111),
.C(n_1874),
.D(n_1940),
.Y(n_2322)
);

NOR3x1_ASAP7_75t_L g2323 ( 
.A(n_2295),
.B(n_138),
.C(n_139),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2313),
.Y(n_2324)
);

AOI221x1_ASAP7_75t_L g2325 ( 
.A1(n_2306),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.C(n_141),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2307),
.Y(n_2326)
);

AOI211xp5_ASAP7_75t_L g2327 ( 
.A1(n_2308),
.A2(n_2072),
.B(n_2070),
.C(n_143),
.Y(n_2327)
);

NAND4xp25_ASAP7_75t_SL g2328 ( 
.A(n_2311),
.B(n_1949),
.C(n_1956),
.D(n_1937),
.Y(n_2328)
);

AOI211xp5_ASAP7_75t_L g2329 ( 
.A1(n_2312),
.A2(n_2072),
.B(n_2070),
.C(n_144),
.Y(n_2329)
);

NOR4xp25_ASAP7_75t_SL g2330 ( 
.A(n_2302),
.B(n_145),
.C(n_141),
.D(n_142),
.Y(n_2330)
);

AOI21xp5_ASAP7_75t_L g2331 ( 
.A1(n_2310),
.A2(n_1907),
.B(n_1901),
.Y(n_2331)
);

OAI22xp5_ASAP7_75t_L g2332 ( 
.A1(n_2303),
.A2(n_2072),
.B1(n_2162),
.B2(n_2133),
.Y(n_2332)
);

INVxp67_ASAP7_75t_L g2333 ( 
.A(n_2298),
.Y(n_2333)
);

NOR3xp33_ASAP7_75t_L g2334 ( 
.A(n_2301),
.B(n_2046),
.C(n_1933),
.Y(n_2334)
);

NAND4xp25_ASAP7_75t_L g2335 ( 
.A(n_2309),
.B(n_1917),
.C(n_146),
.D(n_142),
.Y(n_2335)
);

OAI21xp5_ASAP7_75t_L g2336 ( 
.A1(n_2299),
.A2(n_1919),
.B(n_2148),
.Y(n_2336)
);

OAI21xp5_ASAP7_75t_SL g2337 ( 
.A1(n_2300),
.A2(n_2304),
.B(n_1978),
.Y(n_2337)
);

OAI211xp5_ASAP7_75t_L g2338 ( 
.A1(n_2312),
.A2(n_147),
.B(n_145),
.C(n_146),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2314),
.Y(n_2339)
);

NOR2xp33_ASAP7_75t_L g2340 ( 
.A(n_2315),
.B(n_149),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2314),
.Y(n_2341)
);

NAND3xp33_ASAP7_75t_L g2342 ( 
.A(n_2297),
.B(n_149),
.C(n_150),
.Y(n_2342)
);

NOR2xp33_ASAP7_75t_L g2343 ( 
.A(n_2315),
.B(n_150),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2314),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2315),
.B(n_151),
.Y(n_2345)
);

NAND3xp33_ASAP7_75t_L g2346 ( 
.A(n_2297),
.B(n_151),
.C(n_152),
.Y(n_2346)
);

AOI21xp5_ASAP7_75t_L g2347 ( 
.A1(n_2294),
.A2(n_1818),
.B(n_2050),
.Y(n_2347)
);

OAI211xp5_ASAP7_75t_SL g2348 ( 
.A1(n_2312),
.A2(n_154),
.B(n_152),
.C(n_153),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_2315),
.B(n_153),
.Y(n_2349)
);

NOR3xp33_ASAP7_75t_L g2350 ( 
.A(n_2296),
.B(n_154),
.C(n_155),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_SL g2351 ( 
.A(n_2315),
.B(n_2133),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2315),
.B(n_155),
.Y(n_2352)
);

INVx1_ASAP7_75t_SL g2353 ( 
.A(n_2345),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2349),
.Y(n_2354)
);

BUFx6f_ASAP7_75t_L g2355 ( 
.A(n_2326),
.Y(n_2355)
);

AOI21xp5_ASAP7_75t_L g2356 ( 
.A1(n_2352),
.A2(n_1818),
.B(n_156),
.Y(n_2356)
);

NOR3xp33_ASAP7_75t_SL g2357 ( 
.A(n_2340),
.B(n_156),
.C(n_157),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_2339),
.B(n_2164),
.Y(n_2358)
);

OAI21xp5_ASAP7_75t_L g2359 ( 
.A1(n_2343),
.A2(n_2148),
.B(n_2149),
.Y(n_2359)
);

AND2x2_ASAP7_75t_L g2360 ( 
.A(n_2318),
.B(n_2171),
.Y(n_2360)
);

OAI211xp5_ASAP7_75t_L g2361 ( 
.A1(n_2330),
.A2(n_159),
.B(n_157),
.C(n_158),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2323),
.Y(n_2362)
);

NOR2xp33_ASAP7_75t_L g2363 ( 
.A(n_2348),
.B(n_158),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_2316),
.Y(n_2364)
);

AOI21xp5_ASAP7_75t_L g2365 ( 
.A1(n_2324),
.A2(n_1818),
.B(n_159),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2342),
.Y(n_2366)
);

NAND4xp25_ASAP7_75t_L g2367 ( 
.A(n_2327),
.B(n_162),
.C(n_160),
.D(n_161),
.Y(n_2367)
);

NAND4xp25_ASAP7_75t_L g2368 ( 
.A(n_2320),
.B(n_162),
.C(n_160),
.D(n_161),
.Y(n_2368)
);

OAI211xp5_ASAP7_75t_L g2369 ( 
.A1(n_2329),
.A2(n_165),
.B(n_163),
.C(n_164),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2341),
.B(n_163),
.Y(n_2370)
);

CKINVDCx20_ASAP7_75t_L g2371 ( 
.A(n_2325),
.Y(n_2371)
);

INVxp67_ASAP7_75t_L g2372 ( 
.A(n_2351),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2346),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2344),
.Y(n_2374)
);

NAND3xp33_ASAP7_75t_L g2375 ( 
.A(n_2350),
.B(n_164),
.C(n_165),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2317),
.Y(n_2376)
);

NOR2x1_ASAP7_75t_L g2377 ( 
.A(n_2338),
.B(n_166),
.Y(n_2377)
);

AOI22xp5_ASAP7_75t_L g2378 ( 
.A1(n_2332),
.A2(n_2148),
.B1(n_2133),
.B2(n_2146),
.Y(n_2378)
);

O2A1O1Ixp33_ASAP7_75t_SL g2379 ( 
.A1(n_2333),
.A2(n_168),
.B(n_166),
.C(n_167),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2321),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2337),
.B(n_169),
.Y(n_2381)
);

AOI22xp5_ASAP7_75t_L g2382 ( 
.A1(n_2334),
.A2(n_2133),
.B1(n_2146),
.B2(n_2135),
.Y(n_2382)
);

NOR3x1_ASAP7_75t_L g2383 ( 
.A(n_2335),
.B(n_169),
.C(n_170),
.Y(n_2383)
);

NAND3x1_ASAP7_75t_L g2384 ( 
.A(n_2336),
.B(n_171),
.C(n_172),
.Y(n_2384)
);

OR2x2_ASAP7_75t_L g2385 ( 
.A(n_2328),
.B(n_171),
.Y(n_2385)
);

NOR2xp33_ASAP7_75t_L g2386 ( 
.A(n_2322),
.B(n_173),
.Y(n_2386)
);

O2A1O1Ixp33_ASAP7_75t_L g2387 ( 
.A1(n_2331),
.A2(n_175),
.B(n_173),
.C(n_174),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2347),
.B(n_174),
.Y(n_2388)
);

OR2x2_ASAP7_75t_L g2389 ( 
.A(n_2319),
.B(n_175),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2340),
.B(n_176),
.Y(n_2390)
);

AOI22xp5_ASAP7_75t_SL g2391 ( 
.A1(n_2363),
.A2(n_2133),
.B1(n_2075),
.B2(n_2079),
.Y(n_2391)
);

OR2x2_ASAP7_75t_L g2392 ( 
.A(n_2368),
.B(n_176),
.Y(n_2392)
);

CKINVDCx20_ASAP7_75t_R g2393 ( 
.A(n_2362),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2370),
.Y(n_2394)
);

AOI322xp5_ASAP7_75t_L g2395 ( 
.A1(n_2374),
.A2(n_2105),
.A3(n_2135),
.B1(n_2103),
.B2(n_2168),
.C1(n_2171),
.C2(n_2165),
.Y(n_2395)
);

AOI22xp5_ASAP7_75t_SL g2396 ( 
.A1(n_2372),
.A2(n_2075),
.B1(n_2079),
.B2(n_2077),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2355),
.B(n_2360),
.Y(n_2397)
);

OAI21xp5_ASAP7_75t_L g2398 ( 
.A1(n_2384),
.A2(n_2149),
.B(n_2153),
.Y(n_2398)
);

A2O1A1Ixp33_ASAP7_75t_L g2399 ( 
.A1(n_2361),
.A2(n_179),
.B(n_177),
.C(n_178),
.Y(n_2399)
);

AOI21xp33_ASAP7_75t_SL g2400 ( 
.A1(n_2385),
.A2(n_178),
.B(n_179),
.Y(n_2400)
);

A2O1A1Ixp33_ASAP7_75t_SL g2401 ( 
.A1(n_2354),
.A2(n_182),
.B(n_180),
.C(n_181),
.Y(n_2401)
);

OAI321xp33_ASAP7_75t_L g2402 ( 
.A1(n_2380),
.A2(n_183),
.A3(n_185),
.B1(n_180),
.B2(n_181),
.C(n_184),
.Y(n_2402)
);

AOI22x1_ASAP7_75t_L g2403 ( 
.A1(n_2355),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.Y(n_2403)
);

AOI22xp33_ASAP7_75t_L g2404 ( 
.A1(n_2355),
.A2(n_2135),
.B1(n_2065),
.B2(n_2077),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2379),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2358),
.B(n_2088),
.Y(n_2406)
);

AND2x2_ASAP7_75t_L g2407 ( 
.A(n_2357),
.B(n_2105),
.Y(n_2407)
);

XNOR2x1_ASAP7_75t_L g2408 ( 
.A(n_2377),
.B(n_186),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2390),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_SL g2410 ( 
.A(n_2364),
.B(n_2117),
.Y(n_2410)
);

NAND2x1p5_ASAP7_75t_L g2411 ( 
.A(n_2353),
.B(n_2065),
.Y(n_2411)
);

OAI211xp5_ASAP7_75t_SL g2412 ( 
.A1(n_2366),
.A2(n_188),
.B(n_186),
.C(n_187),
.Y(n_2412)
);

NAND3xp33_ASAP7_75t_SL g2413 ( 
.A(n_2369),
.B(n_187),
.C(n_188),
.Y(n_2413)
);

INVxp67_ASAP7_75t_L g2414 ( 
.A(n_2381),
.Y(n_2414)
);

NOR2x1_ASAP7_75t_L g2415 ( 
.A(n_2367),
.B(n_189),
.Y(n_2415)
);

INVx2_ASAP7_75t_SL g2416 ( 
.A(n_2389),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2375),
.Y(n_2417)
);

NOR2xp67_ASAP7_75t_L g2418 ( 
.A(n_2373),
.B(n_189),
.Y(n_2418)
);

OAI221xp5_ASAP7_75t_L g2419 ( 
.A1(n_2376),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.C(n_193),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2386),
.B(n_190),
.Y(n_2420)
);

OAI21xp5_ASAP7_75t_L g2421 ( 
.A1(n_2387),
.A2(n_2388),
.B(n_2382),
.Y(n_2421)
);

AOI211xp5_ASAP7_75t_L g2422 ( 
.A1(n_2371),
.A2(n_194),
.B(n_191),
.C(n_193),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2383),
.Y(n_2423)
);

OA22x2_ASAP7_75t_L g2424 ( 
.A1(n_2378),
.A2(n_2157),
.B1(n_2158),
.B2(n_2085),
.Y(n_2424)
);

AND2x2_ASAP7_75t_L g2425 ( 
.A(n_2359),
.B(n_2163),
.Y(n_2425)
);

A2O1A1Ixp33_ASAP7_75t_L g2426 ( 
.A1(n_2356),
.A2(n_2365),
.B(n_198),
.C(n_195),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2370),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2355),
.B(n_195),
.Y(n_2428)
);

NAND3xp33_ASAP7_75t_L g2429 ( 
.A(n_2361),
.B(n_196),
.C(n_198),
.Y(n_2429)
);

HB1xp67_ASAP7_75t_L g2430 ( 
.A(n_2355),
.Y(n_2430)
);

NOR2xp67_ASAP7_75t_L g2431 ( 
.A(n_2361),
.B(n_196),
.Y(n_2431)
);

INVxp67_ASAP7_75t_L g2432 ( 
.A(n_2363),
.Y(n_2432)
);

OAI21xp33_ASAP7_75t_L g2433 ( 
.A1(n_2374),
.A2(n_199),
.B(n_200),
.Y(n_2433)
);

AOI211xp5_ASAP7_75t_L g2434 ( 
.A1(n_2361),
.A2(n_203),
.B(n_200),
.C(n_202),
.Y(n_2434)
);

NOR2xp33_ASAP7_75t_L g2435 ( 
.A(n_2355),
.B(n_202),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_SL g2436 ( 
.A(n_2355),
.B(n_2117),
.Y(n_2436)
);

OAI22xp5_ASAP7_75t_L g2437 ( 
.A1(n_2378),
.A2(n_2062),
.B1(n_2068),
.B2(n_2114),
.Y(n_2437)
);

AOI21xp5_ASAP7_75t_L g2438 ( 
.A1(n_2379),
.A2(n_204),
.B(n_205),
.Y(n_2438)
);

NOR4xp75_ASAP7_75t_L g2439 ( 
.A(n_2384),
.B(n_207),
.C(n_204),
.D(n_206),
.Y(n_2439)
);

AOI22xp5_ASAP7_75t_L g2440 ( 
.A1(n_2374),
.A2(n_2101),
.B1(n_2114),
.B2(n_2136),
.Y(n_2440)
);

AOI221xp5_ASAP7_75t_L g2441 ( 
.A1(n_2372),
.A2(n_210),
.B1(n_208),
.B2(n_209),
.C(n_211),
.Y(n_2441)
);

HB1xp67_ASAP7_75t_L g2442 ( 
.A(n_2355),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2370),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2355),
.B(n_208),
.Y(n_2444)
);

AOI22xp33_ASAP7_75t_L g2445 ( 
.A1(n_2355),
.A2(n_2136),
.B1(n_2085),
.B2(n_2159),
.Y(n_2445)
);

INVx1_ASAP7_75t_SL g2446 ( 
.A(n_2370),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2370),
.Y(n_2447)
);

NAND5xp2_ASAP7_75t_L g2448 ( 
.A(n_2362),
.B(n_212),
.C(n_209),
.D(n_210),
.E(n_213),
.Y(n_2448)
);

AOI22xp5_ASAP7_75t_L g2449 ( 
.A1(n_2374),
.A2(n_2101),
.B1(n_2136),
.B2(n_2157),
.Y(n_2449)
);

AOI321xp33_ASAP7_75t_L g2450 ( 
.A1(n_2362),
.A2(n_212),
.A3(n_213),
.B1(n_214),
.B2(n_215),
.C(n_216),
.Y(n_2450)
);

AOI21xp33_ASAP7_75t_L g2451 ( 
.A1(n_2374),
.A2(n_214),
.B(n_215),
.Y(n_2451)
);

INVxp67_ASAP7_75t_L g2452 ( 
.A(n_2363),
.Y(n_2452)
);

INVxp67_ASAP7_75t_L g2453 ( 
.A(n_2363),
.Y(n_2453)
);

AOI21xp5_ASAP7_75t_L g2454 ( 
.A1(n_2379),
.A2(n_217),
.B(n_218),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2403),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2418),
.B(n_2435),
.Y(n_2456)
);

AOI22xp5_ASAP7_75t_L g2457 ( 
.A1(n_2393),
.A2(n_2101),
.B1(n_2158),
.B2(n_2160),
.Y(n_2457)
);

OA22x2_ASAP7_75t_L g2458 ( 
.A1(n_2405),
.A2(n_2085),
.B1(n_221),
.B2(n_218),
.Y(n_2458)
);

NOR2x1_ASAP7_75t_L g2459 ( 
.A(n_2428),
.B(n_220),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2444),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2411),
.Y(n_2461)
);

AO22x2_ASAP7_75t_L g2462 ( 
.A1(n_2408),
.A2(n_223),
.B1(n_220),
.B2(n_222),
.Y(n_2462)
);

HB1xp67_ASAP7_75t_L g2463 ( 
.A(n_2439),
.Y(n_2463)
);

NOR4xp25_ASAP7_75t_L g2464 ( 
.A(n_2413),
.B(n_224),
.C(n_222),
.D(n_223),
.Y(n_2464)
);

OAI22xp5_ASAP7_75t_L g2465 ( 
.A1(n_2404),
.A2(n_2066),
.B1(n_2163),
.B2(n_2160),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2431),
.B(n_225),
.Y(n_2466)
);

OAI22xp5_ASAP7_75t_L g2467 ( 
.A1(n_2429),
.A2(n_2066),
.B1(n_2107),
.B2(n_2049),
.Y(n_2467)
);

OA22x2_ASAP7_75t_SL g2468 ( 
.A1(n_2423),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.Y(n_2468)
);

AOI211xp5_ASAP7_75t_L g2469 ( 
.A1(n_2400),
.A2(n_228),
.B(n_226),
.C(n_227),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2430),
.Y(n_2470)
);

AOI22xp5_ASAP7_75t_L g2471 ( 
.A1(n_2410),
.A2(n_2049),
.B1(n_2090),
.B2(n_2087),
.Y(n_2471)
);

NOR4xp25_ASAP7_75t_L g2472 ( 
.A(n_2397),
.B(n_230),
.C(n_228),
.D(n_229),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_SL g2473 ( 
.A(n_2450),
.B(n_229),
.Y(n_2473)
);

NOR4xp25_ASAP7_75t_L g2474 ( 
.A(n_2417),
.B(n_232),
.C(n_230),
.D(n_231),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2392),
.Y(n_2475)
);

AOI221xp5_ASAP7_75t_L g2476 ( 
.A1(n_2436),
.A2(n_234),
.B1(n_231),
.B2(n_233),
.C(n_235),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2442),
.Y(n_2477)
);

AO22x2_ASAP7_75t_L g2478 ( 
.A1(n_2416),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2407),
.Y(n_2479)
);

AOI22xp5_ASAP7_75t_L g2480 ( 
.A1(n_2415),
.A2(n_2066),
.B1(n_2153),
.B2(n_1860),
.Y(n_2480)
);

AOI22xp5_ASAP7_75t_L g2481 ( 
.A1(n_2412),
.A2(n_2066),
.B1(n_1887),
.B2(n_1903),
.Y(n_2481)
);

OR2x2_ASAP7_75t_L g2482 ( 
.A(n_2448),
.B(n_236),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2399),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2433),
.Y(n_2484)
);

AOI22xp5_ASAP7_75t_L g2485 ( 
.A1(n_2432),
.A2(n_2066),
.B1(n_1939),
.B2(n_1858),
.Y(n_2485)
);

NOR2x1_ASAP7_75t_L g2486 ( 
.A(n_2419),
.B(n_237),
.Y(n_2486)
);

AO22x2_ASAP7_75t_L g2487 ( 
.A1(n_2446),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.Y(n_2487)
);

NOR2x1_ASAP7_75t_L g2488 ( 
.A(n_2433),
.B(n_238),
.Y(n_2488)
);

AOI22xp5_ASAP7_75t_L g2489 ( 
.A1(n_2452),
.A2(n_2071),
.B1(n_2061),
.B2(n_2055),
.Y(n_2489)
);

AO22x2_ASAP7_75t_L g2490 ( 
.A1(n_2394),
.A2(n_2427),
.B1(n_2447),
.B2(n_2443),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2420),
.Y(n_2491)
);

AOI22xp5_ASAP7_75t_L g2492 ( 
.A1(n_2453),
.A2(n_2061),
.B1(n_2055),
.B2(n_2156),
.Y(n_2492)
);

NOR2x1_ASAP7_75t_L g2493 ( 
.A(n_2438),
.B(n_239),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2422),
.B(n_241),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2391),
.Y(n_2495)
);

INVxp67_ASAP7_75t_L g2496 ( 
.A(n_2454),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2434),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2409),
.Y(n_2498)
);

NOR4xp25_ASAP7_75t_L g2499 ( 
.A(n_2414),
.B(n_244),
.C(n_241),
.D(n_242),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2406),
.B(n_242),
.Y(n_2500)
);

AO22x2_ASAP7_75t_L g2501 ( 
.A1(n_2421),
.A2(n_2401),
.B1(n_2437),
.B2(n_2402),
.Y(n_2501)
);

NOR2x1_ASAP7_75t_L g2502 ( 
.A(n_2426),
.B(n_245),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2451),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2424),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2425),
.Y(n_2505)
);

NOR2x1_ASAP7_75t_L g2506 ( 
.A(n_2441),
.B(n_245),
.Y(n_2506)
);

NOR2xp33_ASAP7_75t_L g2507 ( 
.A(n_2396),
.B(n_247),
.Y(n_2507)
);

A2O1A1Ixp33_ASAP7_75t_L g2508 ( 
.A1(n_2398),
.A2(n_250),
.B(n_248),
.C(n_249),
.Y(n_2508)
);

A2O1A1Ixp33_ASAP7_75t_L g2509 ( 
.A1(n_2445),
.A2(n_250),
.B(n_248),
.C(n_249),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2449),
.Y(n_2510)
);

AOI22xp33_ASAP7_75t_L g2511 ( 
.A1(n_2440),
.A2(n_2107),
.B1(n_2069),
.B2(n_2156),
.Y(n_2511)
);

OA22x2_ASAP7_75t_L g2512 ( 
.A1(n_2395),
.A2(n_253),
.B1(n_251),
.B2(n_252),
.Y(n_2512)
);

INVxp67_ASAP7_75t_SL g2513 ( 
.A(n_2418),
.Y(n_2513)
);

INVxp67_ASAP7_75t_L g2514 ( 
.A(n_2448),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2428),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2418),
.B(n_251),
.Y(n_2516)
);

AOI22xp5_ASAP7_75t_L g2517 ( 
.A1(n_2393),
.A2(n_2069),
.B1(n_254),
.B2(n_252),
.Y(n_2517)
);

NOR4xp25_ASAP7_75t_L g2518 ( 
.A(n_2413),
.B(n_255),
.C(n_253),
.D(n_254),
.Y(n_2518)
);

AOI22xp5_ASAP7_75t_L g2519 ( 
.A1(n_2393),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2428),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2428),
.Y(n_2521)
);

AOI22xp5_ASAP7_75t_L g2522 ( 
.A1(n_2393),
.A2(n_259),
.B1(n_256),
.B2(n_258),
.Y(n_2522)
);

OAI22xp5_ASAP7_75t_SL g2523 ( 
.A1(n_2393),
.A2(n_261),
.B1(n_259),
.B2(n_260),
.Y(n_2523)
);

AOI322xp5_ASAP7_75t_L g2524 ( 
.A1(n_2470),
.A2(n_260),
.A3(n_262),
.B1(n_263),
.B2(n_264),
.C1(n_265),
.C2(n_266),
.Y(n_2524)
);

NOR2x1p5_ASAP7_75t_L g2525 ( 
.A(n_2482),
.B(n_263),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2462),
.B(n_264),
.Y(n_2526)
);

NAND3xp33_ASAP7_75t_L g2527 ( 
.A(n_2469),
.B(n_265),
.C(n_266),
.Y(n_2527)
);

NOR3xp33_ASAP7_75t_L g2528 ( 
.A(n_2466),
.B(n_2477),
.C(n_2513),
.Y(n_2528)
);

NAND3xp33_ASAP7_75t_L g2529 ( 
.A(n_2507),
.B(n_267),
.C(n_268),
.Y(n_2529)
);

NAND3xp33_ASAP7_75t_L g2530 ( 
.A(n_2459),
.B(n_268),
.C(n_269),
.Y(n_2530)
);

AND2x2_ASAP7_75t_L g2531 ( 
.A(n_2463),
.B(n_2138),
.Y(n_2531)
);

OAI21xp5_ASAP7_75t_SL g2532 ( 
.A1(n_2514),
.A2(n_269),
.B(n_270),
.Y(n_2532)
);

AOI22xp5_ASAP7_75t_L g2533 ( 
.A1(n_2473),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.Y(n_2533)
);

OAI31xp33_ASAP7_75t_L g2534 ( 
.A1(n_2508),
.A2(n_274),
.A3(n_272),
.B(n_273),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2462),
.Y(n_2535)
);

AND2x2_ASAP7_75t_L g2536 ( 
.A(n_2472),
.B(n_2138),
.Y(n_2536)
);

NAND2x1p5_ASAP7_75t_L g2537 ( 
.A(n_2493),
.B(n_273),
.Y(n_2537)
);

AND2x4_ASAP7_75t_L g2538 ( 
.A(n_2488),
.B(n_274),
.Y(n_2538)
);

NAND3xp33_ASAP7_75t_L g2539 ( 
.A(n_2476),
.B(n_275),
.C(n_276),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2468),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2474),
.B(n_2138),
.Y(n_2541)
);

NOR4xp75_ASAP7_75t_L g2542 ( 
.A(n_2456),
.B(n_277),
.C(n_275),
.D(n_276),
.Y(n_2542)
);

AND2x2_ASAP7_75t_L g2543 ( 
.A(n_2499),
.B(n_2138),
.Y(n_2543)
);

O2A1O1Ixp5_ASAP7_75t_L g2544 ( 
.A1(n_2461),
.A2(n_279),
.B(n_277),
.C(n_278),
.Y(n_2544)
);

INVx2_ASAP7_75t_SL g2545 ( 
.A(n_2458),
.Y(n_2545)
);

INVx3_ASAP7_75t_L g2546 ( 
.A(n_2455),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_2464),
.B(n_2518),
.Y(n_2547)
);

XOR2xp5_ASAP7_75t_L g2548 ( 
.A(n_2501),
.B(n_279),
.Y(n_2548)
);

AOI21xp33_ASAP7_75t_L g2549 ( 
.A1(n_2516),
.A2(n_280),
.B(n_281),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2484),
.B(n_280),
.Y(n_2550)
);

NAND3xp33_ASAP7_75t_L g2551 ( 
.A(n_2495),
.B(n_281),
.C(n_282),
.Y(n_2551)
);

INVxp67_ASAP7_75t_L g2552 ( 
.A(n_2500),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2494),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2512),
.Y(n_2554)
);

NOR3xp33_ASAP7_75t_L g2555 ( 
.A(n_2496),
.B(n_283),
.C(n_284),
.Y(n_2555)
);

NOR3xp33_ASAP7_75t_L g2556 ( 
.A(n_2498),
.B(n_2483),
.C(n_2497),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_L g2557 ( 
.A(n_2509),
.B(n_283),
.Y(n_2557)
);

INVx1_ASAP7_75t_SL g2558 ( 
.A(n_2523),
.Y(n_2558)
);

INVxp67_ASAP7_75t_L g2559 ( 
.A(n_2487),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2487),
.Y(n_2560)
);

AOI22xp5_ASAP7_75t_L g2561 ( 
.A1(n_2479),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.Y(n_2561)
);

OAI211xp5_ASAP7_75t_L g2562 ( 
.A1(n_2486),
.A2(n_287),
.B(n_285),
.C(n_286),
.Y(n_2562)
);

OAI22xp5_ASAP7_75t_L g2563 ( 
.A1(n_2517),
.A2(n_2107),
.B1(n_289),
.B2(n_287),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2501),
.B(n_2138),
.Y(n_2564)
);

OR2x2_ASAP7_75t_L g2565 ( 
.A(n_2505),
.B(n_288),
.Y(n_2565)
);

AND2x4_ASAP7_75t_SL g2566 ( 
.A(n_2475),
.B(n_288),
.Y(n_2566)
);

AOI221xp5_ASAP7_75t_L g2567 ( 
.A1(n_2504),
.A2(n_290),
.B1(n_291),
.B2(n_292),
.C(n_293),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2478),
.Y(n_2568)
);

AND2x2_ASAP7_75t_L g2569 ( 
.A(n_2502),
.B(n_2506),
.Y(n_2569)
);

OR2x2_ASAP7_75t_L g2570 ( 
.A(n_2503),
.B(n_2460),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2478),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2519),
.B(n_290),
.Y(n_2572)
);

OR2x2_ASAP7_75t_L g2573 ( 
.A(n_2515),
.B(n_293),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2522),
.B(n_294),
.Y(n_2574)
);

NOR2x1_ASAP7_75t_L g2575 ( 
.A(n_2520),
.B(n_294),
.Y(n_2575)
);

AND3x2_ASAP7_75t_L g2576 ( 
.A(n_2521),
.B(n_295),
.C(n_296),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2490),
.B(n_297),
.Y(n_2577)
);

NOR2x1_ASAP7_75t_L g2578 ( 
.A(n_2491),
.B(n_298),
.Y(n_2578)
);

AOI221xp5_ASAP7_75t_L g2579 ( 
.A1(n_2510),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.C(n_301),
.Y(n_2579)
);

AND2x4_ASAP7_75t_L g2580 ( 
.A(n_2481),
.B(n_299),
.Y(n_2580)
);

AND2x4_ASAP7_75t_L g2581 ( 
.A(n_2480),
.B(n_300),
.Y(n_2581)
);

NAND3xp33_ASAP7_75t_L g2582 ( 
.A(n_2467),
.B(n_302),
.C(n_304),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_SL g2583 ( 
.A(n_2465),
.B(n_304),
.Y(n_2583)
);

NAND3xp33_ASAP7_75t_L g2584 ( 
.A(n_2485),
.B(n_305),
.C(n_307),
.Y(n_2584)
);

INVxp67_ASAP7_75t_L g2585 ( 
.A(n_2490),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2457),
.B(n_305),
.Y(n_2586)
);

XOR2x2_ASAP7_75t_L g2587 ( 
.A(n_2471),
.B(n_2489),
.Y(n_2587)
);

AND2x4_ASAP7_75t_L g2588 ( 
.A(n_2511),
.B(n_307),
.Y(n_2588)
);

NOR3xp33_ASAP7_75t_L g2589 ( 
.A(n_2585),
.B(n_2492),
.C(n_309),
.Y(n_2589)
);

OR2x2_ASAP7_75t_L g2590 ( 
.A(n_2537),
.B(n_309),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2577),
.Y(n_2591)
);

NAND4xp75_ASAP7_75t_L g2592 ( 
.A(n_2575),
.B(n_310),
.C(n_311),
.D(n_312),
.Y(n_2592)
);

NAND4xp25_ASAP7_75t_L g2593 ( 
.A(n_2556),
.B(n_310),
.C(n_312),
.D(n_313),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_L g2594 ( 
.A(n_2566),
.B(n_313),
.Y(n_2594)
);

AOI211xp5_ASAP7_75t_L g2595 ( 
.A1(n_2562),
.A2(n_2551),
.B(n_2529),
.C(n_2530),
.Y(n_2595)
);

NOR2xp33_ASAP7_75t_L g2596 ( 
.A(n_2548),
.B(n_314),
.Y(n_2596)
);

NOR3xp33_ASAP7_75t_L g2597 ( 
.A(n_2546),
.B(n_314),
.C(n_315),
.Y(n_2597)
);

AOI21xp5_ASAP7_75t_L g2598 ( 
.A1(n_2547),
.A2(n_316),
.B(n_317),
.Y(n_2598)
);

NOR3xp33_ASAP7_75t_L g2599 ( 
.A(n_2528),
.B(n_316),
.C(n_317),
.Y(n_2599)
);

NAND4xp25_ASAP7_75t_L g2600 ( 
.A(n_2533),
.B(n_2534),
.C(n_2527),
.D(n_2554),
.Y(n_2600)
);

NAND4xp25_ASAP7_75t_L g2601 ( 
.A(n_2539),
.B(n_318),
.C(n_320),
.D(n_321),
.Y(n_2601)
);

AOI22xp5_ASAP7_75t_L g2602 ( 
.A1(n_2525),
.A2(n_318),
.B1(n_320),
.B2(n_321),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2576),
.Y(n_2603)
);

NOR2xp67_ASAP7_75t_SL g2604 ( 
.A(n_2535),
.B(n_323),
.Y(n_2604)
);

NAND4xp25_ASAP7_75t_L g2605 ( 
.A(n_2582),
.B(n_323),
.C(n_324),
.D(n_325),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2578),
.Y(n_2606)
);

AOI21xp5_ASAP7_75t_L g2607 ( 
.A1(n_2526),
.A2(n_324),
.B(n_326),
.Y(n_2607)
);

NOR2xp67_ASAP7_75t_L g2608 ( 
.A(n_2559),
.B(n_326),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2573),
.Y(n_2609)
);

NAND4xp25_ASAP7_75t_L g2610 ( 
.A(n_2558),
.B(n_327),
.C(n_328),
.D(n_331),
.Y(n_2610)
);

NOR3xp33_ASAP7_75t_L g2611 ( 
.A(n_2545),
.B(n_327),
.C(n_332),
.Y(n_2611)
);

NOR3xp33_ASAP7_75t_L g2612 ( 
.A(n_2569),
.B(n_333),
.C(n_334),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2538),
.B(n_333),
.Y(n_2613)
);

NOR3xp33_ASAP7_75t_L g2614 ( 
.A(n_2552),
.B(n_334),
.C(n_335),
.Y(n_2614)
);

NOR2x1p5_ASAP7_75t_L g2615 ( 
.A(n_2540),
.B(n_335),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2538),
.B(n_336),
.Y(n_2616)
);

AND4x1_ASAP7_75t_L g2617 ( 
.A(n_2544),
.B(n_336),
.C(n_338),
.D(n_339),
.Y(n_2617)
);

AND2x2_ASAP7_75t_L g2618 ( 
.A(n_2555),
.B(n_339),
.Y(n_2618)
);

AOI22xp33_ASAP7_75t_L g2619 ( 
.A1(n_2564),
.A2(n_340),
.B1(n_341),
.B2(n_342),
.Y(n_2619)
);

OR2x6_ASAP7_75t_L g2620 ( 
.A(n_2571),
.B(n_341),
.Y(n_2620)
);

CKINVDCx5p33_ASAP7_75t_R g2621 ( 
.A(n_2560),
.Y(n_2621)
);

CKINVDCx16_ASAP7_75t_R g2622 ( 
.A(n_2570),
.Y(n_2622)
);

NOR3xp33_ASAP7_75t_L g2623 ( 
.A(n_2553),
.B(n_342),
.C(n_343),
.Y(n_2623)
);

NAND4xp25_ASAP7_75t_L g2624 ( 
.A(n_2572),
.B(n_343),
.C(n_344),
.D(n_345),
.Y(n_2624)
);

AND2x4_ASAP7_75t_L g2625 ( 
.A(n_2542),
.B(n_344),
.Y(n_2625)
);

NOR3xp33_ASAP7_75t_L g2626 ( 
.A(n_2549),
.B(n_345),
.C(n_346),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2532),
.B(n_346),
.Y(n_2627)
);

NAND3xp33_ASAP7_75t_L g2628 ( 
.A(n_2567),
.B(n_347),
.C(n_348),
.Y(n_2628)
);

OAI221xp5_ASAP7_75t_L g2629 ( 
.A1(n_2568),
.A2(n_348),
.B1(n_349),
.B2(n_350),
.C(n_351),
.Y(n_2629)
);

NAND3xp33_ASAP7_75t_L g2630 ( 
.A(n_2579),
.B(n_350),
.C(n_351),
.Y(n_2630)
);

AOI21x1_ASAP7_75t_L g2631 ( 
.A1(n_2550),
.A2(n_352),
.B(n_353),
.Y(n_2631)
);

NOR2xp67_ASAP7_75t_L g2632 ( 
.A(n_2561),
.B(n_352),
.Y(n_2632)
);

INVx4_ASAP7_75t_L g2633 ( 
.A(n_2565),
.Y(n_2633)
);

NOR3x1_ASAP7_75t_L g2634 ( 
.A(n_2574),
.B(n_353),
.C(n_354),
.Y(n_2634)
);

NAND4xp25_ASAP7_75t_L g2635 ( 
.A(n_2557),
.B(n_354),
.C(n_355),
.D(n_356),
.Y(n_2635)
);

OAI21xp5_ASAP7_75t_L g2636 ( 
.A1(n_2563),
.A2(n_355),
.B(n_357),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2604),
.Y(n_2637)
);

OAI21xp33_ASAP7_75t_SL g2638 ( 
.A1(n_2619),
.A2(n_2536),
.B(n_2543),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2613),
.Y(n_2639)
);

NAND4xp75_ASAP7_75t_L g2640 ( 
.A(n_2608),
.B(n_2586),
.C(n_2583),
.D(n_2541),
.Y(n_2640)
);

NOR3x2_ASAP7_75t_L g2641 ( 
.A(n_2592),
.B(n_2584),
.C(n_2524),
.Y(n_2641)
);

NOR3x1_ASAP7_75t_L g2642 ( 
.A(n_2635),
.B(n_2587),
.C(n_2588),
.Y(n_2642)
);

AOI221xp5_ASAP7_75t_L g2643 ( 
.A1(n_2596),
.A2(n_2581),
.B1(n_2580),
.B2(n_2531),
.C(n_361),
.Y(n_2643)
);

NAND4xp75_ASAP7_75t_L g2644 ( 
.A(n_2634),
.B(n_2581),
.C(n_359),
.D(n_360),
.Y(n_2644)
);

NOR3xp33_ASAP7_75t_L g2645 ( 
.A(n_2622),
.B(n_358),
.C(n_359),
.Y(n_2645)
);

NAND4xp25_ASAP7_75t_L g2646 ( 
.A(n_2595),
.B(n_358),
.C(n_360),
.D(n_362),
.Y(n_2646)
);

AO22x2_ASAP7_75t_L g2647 ( 
.A1(n_2591),
.A2(n_362),
.B1(n_363),
.B2(n_364),
.Y(n_2647)
);

NOR3x1_ASAP7_75t_L g2648 ( 
.A(n_2616),
.B(n_363),
.C(n_364),
.Y(n_2648)
);

AND2x2_ASAP7_75t_L g2649 ( 
.A(n_2625),
.B(n_365),
.Y(n_2649)
);

NOR3xp33_ASAP7_75t_L g2650 ( 
.A(n_2633),
.B(n_365),
.C(n_366),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_2602),
.B(n_368),
.Y(n_2651)
);

INVxp67_ASAP7_75t_L g2652 ( 
.A(n_2620),
.Y(n_2652)
);

OR2x2_ASAP7_75t_L g2653 ( 
.A(n_2605),
.B(n_368),
.Y(n_2653)
);

NOR3xp33_ASAP7_75t_L g2654 ( 
.A(n_2633),
.B(n_369),
.C(n_370),
.Y(n_2654)
);

NOR2xp67_ASAP7_75t_L g2655 ( 
.A(n_2610),
.B(n_369),
.Y(n_2655)
);

NOR2xp33_ASAP7_75t_L g2656 ( 
.A(n_2594),
.B(n_370),
.Y(n_2656)
);

XOR2xp5_ASAP7_75t_L g2657 ( 
.A(n_2624),
.B(n_371),
.Y(n_2657)
);

AOI21xp5_ASAP7_75t_L g2658 ( 
.A1(n_2606),
.A2(n_2603),
.B(n_2627),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2611),
.B(n_371),
.Y(n_2659)
);

OR2x2_ASAP7_75t_L g2660 ( 
.A(n_2590),
.B(n_372),
.Y(n_2660)
);

BUFx2_ASAP7_75t_L g2661 ( 
.A(n_2620),
.Y(n_2661)
);

NAND3xp33_ASAP7_75t_L g2662 ( 
.A(n_2599),
.B(n_373),
.C(n_374),
.Y(n_2662)
);

NAND4xp25_ASAP7_75t_L g2663 ( 
.A(n_2600),
.B(n_373),
.C(n_374),
.D(n_375),
.Y(n_2663)
);

NAND4xp75_ASAP7_75t_L g2664 ( 
.A(n_2607),
.B(n_375),
.C(n_376),
.D(n_377),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_L g2665 ( 
.A(n_2625),
.B(n_377),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2631),
.Y(n_2666)
);

NAND3xp33_ASAP7_75t_SL g2667 ( 
.A(n_2621),
.B(n_2617),
.C(n_2626),
.Y(n_2667)
);

OR2x2_ASAP7_75t_L g2668 ( 
.A(n_2601),
.B(n_378),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2615),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2618),
.Y(n_2670)
);

OAI22xp33_ASAP7_75t_L g2671 ( 
.A1(n_2628),
.A2(n_378),
.B1(n_380),
.B2(n_381),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2636),
.Y(n_2672)
);

AND3x4_ASAP7_75t_L g2673 ( 
.A(n_2632),
.B(n_380),
.C(n_381),
.Y(n_2673)
);

INVx3_ASAP7_75t_L g2674 ( 
.A(n_2609),
.Y(n_2674)
);

NOR2xp33_ASAP7_75t_L g2675 ( 
.A(n_2660),
.B(n_2665),
.Y(n_2675)
);

AND2x4_ASAP7_75t_L g2676 ( 
.A(n_2674),
.B(n_2649),
.Y(n_2676)
);

INVx3_ASAP7_75t_L g2677 ( 
.A(n_2666),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2647),
.Y(n_2678)
);

NAND3xp33_ASAP7_75t_SL g2679 ( 
.A(n_2673),
.B(n_2643),
.C(n_2661),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2648),
.Y(n_2680)
);

OAI22xp5_ASAP7_75t_L g2681 ( 
.A1(n_2657),
.A2(n_2653),
.B1(n_2668),
.B2(n_2662),
.Y(n_2681)
);

INVx3_ASAP7_75t_L g2682 ( 
.A(n_2641),
.Y(n_2682)
);

NOR2x1_ASAP7_75t_L g2683 ( 
.A(n_2664),
.B(n_2593),
.Y(n_2683)
);

NOR2x1_ASAP7_75t_L g2684 ( 
.A(n_2644),
.B(n_2598),
.Y(n_2684)
);

NOR3xp33_ASAP7_75t_L g2685 ( 
.A(n_2667),
.B(n_2630),
.C(n_2597),
.Y(n_2685)
);

NAND3xp33_ASAP7_75t_L g2686 ( 
.A(n_2638),
.B(n_2612),
.C(n_2623),
.Y(n_2686)
);

AND2x2_ASAP7_75t_L g2687 ( 
.A(n_2637),
.B(n_2589),
.Y(n_2687)
);

NOR2x1_ASAP7_75t_L g2688 ( 
.A(n_2663),
.B(n_2629),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2659),
.Y(n_2689)
);

NOR3x2_ASAP7_75t_L g2690 ( 
.A(n_2640),
.B(n_2614),
.C(n_383),
.Y(n_2690)
);

OR3x1_ASAP7_75t_L g2691 ( 
.A(n_2646),
.B(n_382),
.C(n_385),
.Y(n_2691)
);

NAND3x1_ASAP7_75t_L g2692 ( 
.A(n_2669),
.B(n_385),
.C(n_386),
.Y(n_2692)
);

AND2x2_ASAP7_75t_L g2693 ( 
.A(n_2655),
.B(n_386),
.Y(n_2693)
);

NOR3xp33_ASAP7_75t_L g2694 ( 
.A(n_2652),
.B(n_387),
.C(n_388),
.Y(n_2694)
);

NOR3xp33_ASAP7_75t_L g2695 ( 
.A(n_2658),
.B(n_387),
.C(n_388),
.Y(n_2695)
);

NOR3xp33_ASAP7_75t_L g2696 ( 
.A(n_2672),
.B(n_389),
.C(n_390),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2656),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2647),
.Y(n_2698)
);

NOR3xp33_ASAP7_75t_SL g2699 ( 
.A(n_2671),
.B(n_389),
.C(n_390),
.Y(n_2699)
);

XOR2xp5_ASAP7_75t_L g2700 ( 
.A(n_2651),
.B(n_391),
.Y(n_2700)
);

NOR3xp33_ASAP7_75t_L g2701 ( 
.A(n_2639),
.B(n_392),
.C(n_393),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_2695),
.B(n_2645),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2693),
.B(n_2650),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2700),
.Y(n_2704)
);

XOR2x2_ASAP7_75t_L g2705 ( 
.A(n_2683),
.B(n_2692),
.Y(n_2705)
);

AOI22xp5_ASAP7_75t_L g2706 ( 
.A1(n_2691),
.A2(n_2670),
.B1(n_2654),
.B2(n_2642),
.Y(n_2706)
);

INVx2_ASAP7_75t_SL g2707 ( 
.A(n_2678),
.Y(n_2707)
);

AND2x2_ASAP7_75t_L g2708 ( 
.A(n_2699),
.B(n_392),
.Y(n_2708)
);

INVx1_ASAP7_75t_SL g2709 ( 
.A(n_2690),
.Y(n_2709)
);

NOR2x1_ASAP7_75t_L g2710 ( 
.A(n_2698),
.B(n_393),
.Y(n_2710)
);

O2A1O1Ixp33_ASAP7_75t_L g2711 ( 
.A1(n_2682),
.A2(n_2677),
.B(n_2679),
.C(n_2681),
.Y(n_2711)
);

NAND3xp33_ASAP7_75t_SL g2712 ( 
.A(n_2685),
.B(n_394),
.C(n_395),
.Y(n_2712)
);

AND2x4_ASAP7_75t_L g2713 ( 
.A(n_2676),
.B(n_394),
.Y(n_2713)
);

AOI22xp5_ASAP7_75t_L g2714 ( 
.A1(n_2680),
.A2(n_2687),
.B1(n_2686),
.B2(n_2688),
.Y(n_2714)
);

OA21x2_ASAP7_75t_L g2715 ( 
.A1(n_2675),
.A2(n_395),
.B(n_396),
.Y(n_2715)
);

AOI21xp5_ASAP7_75t_L g2716 ( 
.A1(n_2684),
.A2(n_396),
.B(n_397),
.Y(n_2716)
);

XNOR2xp5_ASAP7_75t_L g2717 ( 
.A(n_2697),
.B(n_397),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2689),
.Y(n_2718)
);

HB1xp67_ASAP7_75t_L g2719 ( 
.A(n_2694),
.Y(n_2719)
);

INVx3_ASAP7_75t_L g2720 ( 
.A(n_2696),
.Y(n_2720)
);

CKINVDCx16_ASAP7_75t_R g2721 ( 
.A(n_2701),
.Y(n_2721)
);

XNOR2x1_ASAP7_75t_L g2722 ( 
.A(n_2683),
.B(n_398),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2700),
.Y(n_2723)
);

AOI22xp5_ASAP7_75t_L g2724 ( 
.A1(n_2691),
.A2(n_398),
.B1(n_399),
.B2(n_400),
.Y(n_2724)
);

INVx3_ASAP7_75t_L g2725 ( 
.A(n_2692),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2695),
.B(n_400),
.Y(n_2726)
);

AOI21xp5_ASAP7_75t_L g2727 ( 
.A1(n_2678),
.A2(n_401),
.B(n_402),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_2715),
.Y(n_2728)
);

OAI22xp5_ASAP7_75t_L g2729 ( 
.A1(n_2724),
.A2(n_401),
.B1(n_403),
.B2(n_404),
.Y(n_2729)
);

BUFx2_ASAP7_75t_L g2730 ( 
.A(n_2710),
.Y(n_2730)
);

AO22x2_ASAP7_75t_L g2731 ( 
.A1(n_2722),
.A2(n_403),
.B1(n_404),
.B2(n_405),
.Y(n_2731)
);

XOR2xp5_ASAP7_75t_L g2732 ( 
.A(n_2714),
.B(n_405),
.Y(n_2732)
);

OAI22xp5_ASAP7_75t_L g2733 ( 
.A1(n_2707),
.A2(n_2706),
.B1(n_2726),
.B2(n_2709),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2708),
.Y(n_2734)
);

INVxp67_ASAP7_75t_L g2735 ( 
.A(n_2712),
.Y(n_2735)
);

AOI22x1_ASAP7_75t_L g2736 ( 
.A1(n_2725),
.A2(n_406),
.B1(n_407),
.B2(n_408),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2705),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2703),
.Y(n_2738)
);

OA22x2_ASAP7_75t_L g2739 ( 
.A1(n_2719),
.A2(n_406),
.B1(n_408),
.B2(n_409),
.Y(n_2739)
);

INVx2_ASAP7_75t_L g2740 ( 
.A(n_2713),
.Y(n_2740)
);

OA22x2_ASAP7_75t_L g2741 ( 
.A1(n_2718),
.A2(n_409),
.B1(n_410),
.B2(n_411),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2717),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2702),
.Y(n_2743)
);

OAI22xp5_ASAP7_75t_L g2744 ( 
.A1(n_2732),
.A2(n_2737),
.B1(n_2735),
.B2(n_2731),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2741),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2739),
.Y(n_2746)
);

AOI22x1_ASAP7_75t_SL g2747 ( 
.A1(n_2740),
.A2(n_2723),
.B1(n_2704),
.B2(n_2720),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2730),
.Y(n_2748)
);

AOI221xp5_ASAP7_75t_L g2749 ( 
.A1(n_2733),
.A2(n_2711),
.B1(n_2729),
.B2(n_2728),
.C(n_2716),
.Y(n_2749)
);

HB1xp67_ASAP7_75t_L g2750 ( 
.A(n_2736),
.Y(n_2750)
);

NOR2xp33_ASAP7_75t_L g2751 ( 
.A(n_2738),
.B(n_2721),
.Y(n_2751)
);

OAI22xp5_ASAP7_75t_L g2752 ( 
.A1(n_2742),
.A2(n_2727),
.B1(n_411),
.B2(n_412),
.Y(n_2752)
);

HB1xp67_ASAP7_75t_L g2753 ( 
.A(n_2734),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2752),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2750),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2746),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2745),
.Y(n_2757)
);

INVxp33_ASAP7_75t_L g2758 ( 
.A(n_2751),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2748),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2753),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2747),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2760),
.Y(n_2762)
);

AOI21xp5_ASAP7_75t_L g2763 ( 
.A1(n_2759),
.A2(n_2761),
.B(n_2744),
.Y(n_2763)
);

OAI22xp5_ASAP7_75t_SL g2764 ( 
.A1(n_2756),
.A2(n_2743),
.B1(n_2749),
.B2(n_413),
.Y(n_2764)
);

AOI22xp33_ASAP7_75t_L g2765 ( 
.A1(n_2757),
.A2(n_410),
.B1(n_412),
.B2(n_414),
.Y(n_2765)
);

AOI22xp33_ASAP7_75t_SL g2766 ( 
.A1(n_2755),
.A2(n_414),
.B1(n_415),
.B2(n_416),
.Y(n_2766)
);

AO22x1_ASAP7_75t_L g2767 ( 
.A1(n_2758),
.A2(n_417),
.B1(n_418),
.B2(n_419),
.Y(n_2767)
);

OAI22xp5_ASAP7_75t_L g2768 ( 
.A1(n_2762),
.A2(n_2754),
.B1(n_419),
.B2(n_420),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2764),
.Y(n_2769)
);

OAI21xp33_ASAP7_75t_L g2770 ( 
.A1(n_2763),
.A2(n_417),
.B(n_420),
.Y(n_2770)
);

OR2x6_ASAP7_75t_L g2771 ( 
.A(n_2767),
.B(n_421),
.Y(n_2771)
);

NAND2xp33_ASAP7_75t_SL g2772 ( 
.A(n_2769),
.B(n_2765),
.Y(n_2772)
);

AOI22xp5_ASAP7_75t_L g2773 ( 
.A1(n_2771),
.A2(n_2766),
.B1(n_422),
.B2(n_423),
.Y(n_2773)
);

AOI22xp5_ASAP7_75t_L g2774 ( 
.A1(n_2770),
.A2(n_421),
.B1(n_422),
.B2(n_424),
.Y(n_2774)
);

AOI21xp5_ASAP7_75t_L g2775 ( 
.A1(n_2768),
.A2(n_425),
.B(n_426),
.Y(n_2775)
);

OAI22xp5_ASAP7_75t_L g2776 ( 
.A1(n_2773),
.A2(n_425),
.B1(n_427),
.B2(n_428),
.Y(n_2776)
);

AOI22xp5_ASAP7_75t_L g2777 ( 
.A1(n_2772),
.A2(n_427),
.B1(n_428),
.B2(n_429),
.Y(n_2777)
);

AOI22xp33_ASAP7_75t_SL g2778 ( 
.A1(n_2776),
.A2(n_2775),
.B1(n_2774),
.B2(n_433),
.Y(n_2778)
);

AOI21xp5_ASAP7_75t_L g2779 ( 
.A1(n_2778),
.A2(n_2777),
.B(n_431),
.Y(n_2779)
);

OAI22xp5_ASAP7_75t_L g2780 ( 
.A1(n_2779),
.A2(n_430),
.B1(n_431),
.B2(n_433),
.Y(n_2780)
);

OAI221xp5_ASAP7_75t_R g2781 ( 
.A1(n_2780),
.A2(n_430),
.B1(n_434),
.B2(n_435),
.C(n_436),
.Y(n_2781)
);

AOI22xp33_ASAP7_75t_L g2782 ( 
.A1(n_2781),
.A2(n_434),
.B1(n_435),
.B2(n_436),
.Y(n_2782)
);

AOI211xp5_ASAP7_75t_L g2783 ( 
.A1(n_2782),
.A2(n_437),
.B(n_438),
.C(n_439),
.Y(n_2783)
);


endmodule