module fake_jpeg_31426_n_516 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_516);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_516;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_19),
.B(n_17),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_52),
.B(n_43),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_55),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_25),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_57),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_16),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_25),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_58),
.B(n_60),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_70),
.Y(n_112)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_69),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_71),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_74),
.Y(n_122)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_32),
.B(n_14),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_76),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_31),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_77),
.B(n_80),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_31),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

INVx6_ASAP7_75t_SL g83 ( 
.A(n_47),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_83),
.Y(n_105)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_31),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_85),
.B(n_90),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

BUFx10_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_23),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_34),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_95),
.B(n_21),
.Y(n_152)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_18),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_18),
.Y(n_98)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_18),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_97),
.A2(n_43),
.B(n_32),
.C(n_28),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_104),
.B(n_152),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_L g118 ( 
.A1(n_67),
.A2(n_20),
.B1(n_49),
.B2(n_39),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_118),
.A2(n_96),
.B1(n_61),
.B2(n_82),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_121),
.B(n_146),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_66),
.A2(n_48),
.B1(n_49),
.B2(n_20),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_125),
.A2(n_71),
.B1(n_75),
.B2(n_78),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_128),
.Y(n_174)
);

BUFx12_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

CKINVDCx12_ASAP7_75t_R g181 ( 
.A(n_130),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_89),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_134),
.B(n_145),
.Y(n_218)
);

A2O1A1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_90),
.A2(n_50),
.B(n_29),
.C(n_23),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_140),
.B(n_37),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_51),
.Y(n_142)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_142),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_53),
.Y(n_144)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_144),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_70),
.B(n_29),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_89),
.B(n_22),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_59),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_155),
.Y(n_167)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_55),
.Y(n_158)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_161),
.A2(n_202),
.B1(n_205),
.B2(n_210),
.Y(n_220)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_162),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_164),
.Y(n_245)
);

NAND3xp33_ASAP7_75t_L g238 ( 
.A(n_166),
.B(n_171),
.C(n_187),
.Y(n_238)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_168),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_36),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_169),
.B(n_178),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_143),
.B(n_37),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_172),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_102),
.B(n_122),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_173),
.B(n_176),
.Y(n_239)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_106),
.Y(n_175)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_175),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_102),
.B(n_21),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_177),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_36),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_122),
.B(n_21),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_179),
.B(n_180),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_111),
.B(n_21),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_111),
.B(n_62),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_182),
.B(n_184),
.Y(n_259)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_183),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_132),
.B(n_68),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_185),
.A2(n_117),
.B1(n_155),
.B2(n_144),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_112),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_195),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_152),
.B(n_28),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_119),
.A2(n_91),
.B1(n_64),
.B2(n_69),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_188),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_105),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_189),
.B(n_215),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_112),
.A2(n_101),
.B(n_76),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_190),
.Y(n_264)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_103),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_191),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_109),
.B(n_40),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_213),
.Y(n_235)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_108),
.Y(n_193)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_135),
.Y(n_194)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_194),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_127),
.B(n_72),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_110),
.Y(n_196)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_196),
.Y(n_246)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_115),
.Y(n_197)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_154),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_199),
.B(n_201),
.Y(n_249)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_150),
.Y(n_200)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_200),
.Y(n_254)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_139),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_125),
.A2(n_79),
.B1(n_87),
.B2(n_86),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_127),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_203),
.B(n_204),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_128),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_L g205 ( 
.A1(n_120),
.A2(n_94),
.B1(n_20),
.B2(n_49),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_128),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_206),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_124),
.B(n_22),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_207),
.B(n_127),
.Y(n_228)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_133),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_209),
.A2(n_157),
.B1(n_114),
.B2(n_107),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_118),
.A2(n_39),
.B1(n_33),
.B2(n_40),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_131),
.B(n_93),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_123),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g212 ( 
.A(n_157),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_212),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_148),
.B(n_33),
.Y(n_213)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_153),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_214),
.Y(n_253)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_119),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_151),
.B(n_72),
.C(n_39),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_217),
.B(n_190),
.C(n_211),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_161),
.A2(n_149),
.B1(n_141),
.B2(n_129),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_221),
.A2(n_222),
.B1(n_224),
.B2(n_194),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_163),
.A2(n_159),
.B1(n_136),
.B2(n_113),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_156),
.B1(n_103),
.B2(n_117),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_225),
.A2(n_257),
.B1(n_203),
.B2(n_167),
.Y(n_274)
);

OA22x2_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_155),
.B1(n_144),
.B2(n_142),
.Y(n_227)
);

AO22x1_ASAP7_75t_L g300 ( 
.A1(n_227),
.A2(n_266),
.B1(n_6),
.B2(n_7),
.Y(n_300)
);

NAND3xp33_ASAP7_75t_L g278 ( 
.A(n_228),
.B(n_181),
.C(n_216),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_192),
.A2(n_116),
.B1(n_129),
.B2(n_142),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_231),
.A2(n_258),
.B1(n_164),
.B2(n_174),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_169),
.B(n_9),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_236),
.B(n_8),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_237),
.Y(n_275)
);

A2O1A1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_178),
.A2(n_14),
.B(n_13),
.C(n_12),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_240),
.A2(n_3),
.B(n_4),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_242),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_212),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_265),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_208),
.B(n_12),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_256),
.B(n_1),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_209),
.A2(n_130),
.B1(n_10),
.B2(n_9),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_213),
.A2(n_10),
.B1(n_9),
.B2(n_2),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_216),
.C(n_198),
.Y(n_286)
);

AOI22x1_ASAP7_75t_SL g262 ( 
.A1(n_218),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_262)
);

NOR2x1_ASAP7_75t_R g294 ( 
.A(n_262),
.B(n_165),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_212),
.Y(n_265)
);

NOR2x1_ASAP7_75t_L g266 ( 
.A(n_211),
.B(n_0),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_267),
.Y(n_339)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_252),
.Y(n_268)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_268),
.Y(n_318)
);

AND2x6_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_189),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_269),
.B(n_278),
.Y(n_328)
);

INVx13_ASAP7_75t_L g270 ( 
.A(n_245),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_270),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_271),
.Y(n_316)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_272),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_273),
.B(n_284),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_274),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_261),
.A2(n_191),
.B1(n_170),
.B2(n_168),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_276),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_264),
.A2(n_175),
.B1(n_196),
.B2(n_193),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_279),
.A2(n_287),
.B1(n_289),
.B2(n_221),
.Y(n_311)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_254),
.Y(n_281)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_281),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_220),
.A2(n_217),
.B1(n_172),
.B2(n_162),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_282),
.A2(n_285),
.B1(n_249),
.B2(n_223),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_233),
.B(n_214),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_283),
.B(n_290),
.Y(n_343)
);

AND2x6_ASAP7_75t_L g284 ( 
.A(n_238),
.B(n_201),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_286),
.B(n_227),
.C(n_242),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_220),
.A2(n_198),
.B1(n_206),
.B2(n_165),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_297),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_231),
.A2(n_261),
.B1(n_235),
.B2(n_239),
.Y(n_289)
);

INVx11_ASAP7_75t_L g291 ( 
.A(n_241),
.Y(n_291)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_291),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_239),
.B(n_206),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_292),
.B(n_298),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_260),
.A2(n_165),
.B(n_212),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_293),
.A2(n_309),
.B(n_227),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_294),
.A2(n_300),
.B(n_303),
.Y(n_320)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_219),
.Y(n_295)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_295),
.Y(n_337)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_243),
.Y(n_296)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_296),
.Y(n_345)
);

INVx6_ASAP7_75t_SL g297 ( 
.A(n_251),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_248),
.B(n_5),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_245),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_299),
.A2(n_243),
.B1(n_265),
.B2(n_241),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_248),
.B(n_6),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_301),
.B(n_302),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_259),
.B(n_228),
.Y(n_302)
);

OR2x2_ASAP7_75t_SL g303 ( 
.A(n_262),
.B(n_6),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_235),
.B(n_6),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_305),
.Y(n_321)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_219),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_308),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_259),
.A2(n_8),
.B(n_244),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_307),
.A2(n_240),
.B(n_256),
.Y(n_326)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_223),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_242),
.A2(n_8),
.B1(n_266),
.B2(n_225),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_233),
.B(n_263),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_310),
.B(n_236),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_311),
.A2(n_312),
.B1(n_324),
.B2(n_336),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_289),
.A2(n_244),
.B1(n_263),
.B2(n_232),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_317),
.B(n_348),
.C(n_349),
.Y(n_361)
);

AO22x1_ASAP7_75t_SL g322 ( 
.A1(n_300),
.A2(n_227),
.B1(n_266),
.B2(n_263),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_322),
.B(n_331),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_323),
.A2(n_325),
.B1(n_276),
.B2(n_275),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_273),
.A2(n_310),
.B1(n_294),
.B2(n_309),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_SL g382 ( 
.A(n_326),
.B(n_270),
.C(n_8),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_304),
.B(n_280),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_333),
.B(n_347),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_334),
.A2(n_275),
.B(n_277),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_300),
.A2(n_226),
.B1(n_255),
.B2(n_253),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_307),
.A2(n_250),
.B(n_229),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_338),
.A2(n_315),
.B(n_313),
.Y(n_350)
);

AOI22x1_ASAP7_75t_SL g341 ( 
.A1(n_269),
.A2(n_226),
.B1(n_253),
.B2(n_247),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_341),
.B(n_234),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_271),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_344),
.B(n_297),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_303),
.A2(n_246),
.B1(n_229),
.B2(n_230),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_346),
.A2(n_285),
.B1(n_291),
.B2(n_272),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_283),
.B(n_246),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_286),
.B(n_230),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_293),
.B(n_234),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_350),
.A2(n_358),
.B(n_374),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_319),
.B(n_306),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_351),
.B(n_371),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_352),
.Y(n_385)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_318),
.Y(n_355)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_355),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_314),
.A2(n_340),
.B1(n_323),
.B2(n_341),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_356),
.A2(n_365),
.B1(n_379),
.B2(n_342),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_330),
.B(n_288),
.Y(n_359)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_359),
.Y(n_393)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_318),
.Y(n_360)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_360),
.Y(n_397)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_327),
.Y(n_362)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_362),
.Y(n_409)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_327),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_363),
.B(n_366),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_330),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_364),
.B(n_372),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_349),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_348),
.B(n_277),
.C(n_305),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_367),
.B(n_361),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_368),
.B(n_369),
.Y(n_394)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_329),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_321),
.B(n_281),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_370),
.B(n_373),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_315),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_333),
.B(n_247),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_329),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_334),
.A2(n_290),
.B(n_267),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_312),
.B(n_296),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_375),
.B(n_376),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_336),
.Y(n_376)
);

AND2x6_ASAP7_75t_L g377 ( 
.A(n_328),
.B(n_284),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_377),
.A2(n_381),
.B(n_382),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_321),
.B(n_268),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_378),
.B(n_337),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_340),
.A2(n_295),
.B1(n_308),
.B2(n_299),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_335),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_380),
.B(n_337),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_324),
.A2(n_311),
.B1(n_342),
.B2(n_346),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_383),
.A2(n_338),
.B1(n_322),
.B2(n_320),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_382),
.Y(n_387)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_387),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_388),
.B(n_404),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_389),
.B(n_392),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_364),
.B(n_331),
.Y(n_390)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_390),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_356),
.A2(n_335),
.B1(n_317),
.B2(n_320),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_353),
.B(n_326),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_399),
.Y(n_416)
);

OA21x2_ASAP7_75t_L g401 ( 
.A1(n_353),
.A2(n_322),
.B(n_347),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_401),
.A2(n_362),
.B(n_369),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_402),
.A2(n_376),
.B1(n_357),
.B2(n_383),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_403),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_361),
.B(n_343),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_381),
.A2(n_316),
.B(n_343),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_406),
.B(n_412),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_410),
.Y(n_422)
);

NOR4xp25_ASAP7_75t_L g408 ( 
.A(n_354),
.B(n_339),
.C(n_332),
.D(n_345),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_408),
.B(n_368),
.Y(n_430)
);

NOR2x1_ASAP7_75t_L g410 ( 
.A(n_381),
.B(n_332),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_354),
.B(n_359),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_411),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_370),
.B(n_316),
.Y(n_412)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_395),
.Y(n_415)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_415),
.Y(n_438)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_395),
.Y(n_417)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_417),
.Y(n_441)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_407),
.Y(n_419)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_419),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_388),
.B(n_366),
.C(n_367),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_420),
.B(n_423),
.C(n_435),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_404),
.B(n_350),
.C(n_378),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_390),
.B(n_380),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_424),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_405),
.B(n_377),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_426),
.B(n_428),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_399),
.B(n_385),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_427),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_430),
.B(n_431),
.Y(n_448)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_384),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_385),
.B(n_357),
.Y(n_432)
);

INVxp33_ASAP7_75t_L g451 ( 
.A(n_432),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_402),
.A2(n_398),
.B1(n_410),
.B2(n_391),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_433),
.A2(n_401),
.B1(n_408),
.B2(n_400),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_386),
.B(n_358),
.C(n_374),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_392),
.B(n_379),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_436),
.B(n_400),
.C(n_386),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_437),
.B(n_394),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_422),
.B(n_416),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_440),
.B(n_452),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_414),
.A2(n_391),
.B1(n_389),
.B2(n_393),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_443),
.B(n_449),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_434),
.A2(n_387),
.B1(n_393),
.B2(n_396),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_447),
.B(n_454),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_418),
.B(n_420),
.C(n_423),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_450),
.B(n_421),
.C(n_436),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_418),
.B(n_406),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_457),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_425),
.A2(n_387),
.B1(n_410),
.B2(n_384),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_414),
.A2(n_409),
.B1(n_397),
.B2(n_355),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_455),
.B(n_431),
.Y(n_459)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_456),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_435),
.B(n_394),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_439),
.B(n_424),
.Y(n_458)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_458),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_459),
.B(n_462),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_461),
.B(n_472),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_442),
.B(n_429),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_445),
.A2(n_419),
.B1(n_415),
.B2(n_417),
.Y(n_463)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_463),
.Y(n_485)
);

INVx13_ASAP7_75t_L g464 ( 
.A(n_440),
.Y(n_464)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_464),
.Y(n_486)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_438),
.Y(n_467)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_467),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_429),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_470),
.B(n_422),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_446),
.B(n_421),
.C(n_433),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_471),
.B(n_473),
.C(n_457),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_448),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_446),
.B(n_428),
.C(n_413),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_469),
.A2(n_442),
.B1(n_441),
.B2(n_449),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_474),
.B(n_478),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_475),
.B(n_480),
.Y(n_489)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_477),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_460),
.B(n_453),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_460),
.B(n_450),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_482),
.C(n_478),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_458),
.B(n_409),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_469),
.A2(n_456),
.B1(n_444),
.B2(n_443),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_481),
.B(n_466),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_452),
.C(n_437),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_474),
.A2(n_465),
.B1(n_473),
.B2(n_461),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_488),
.B(n_491),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_484),
.B(n_451),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_492),
.B(n_493),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_475),
.B(n_482),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_483),
.A2(n_464),
.B(n_401),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_495),
.A2(n_496),
.B(n_477),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_476),
.B(n_466),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_497),
.B(n_479),
.C(n_490),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_498),
.B(n_499),
.Y(n_506)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_489),
.A2(n_480),
.B(n_481),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_501),
.A2(n_502),
.B(n_495),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_497),
.B(n_486),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_503),
.B(n_494),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_504),
.B(n_505),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_500),
.B(n_488),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_507),
.B(n_490),
.Y(n_509)
);

AOI322xp5_ASAP7_75t_L g511 ( 
.A1(n_509),
.A2(n_487),
.A3(n_345),
.B1(n_397),
.B2(n_363),
.C1(n_373),
.C2(n_360),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_508),
.A2(n_506),
.B(n_485),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_510),
.B(n_511),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_512),
.A2(n_316),
.B(n_468),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_513),
.A2(n_468),
.B(n_430),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_514),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_515),
.Y(n_516)
);


endmodule