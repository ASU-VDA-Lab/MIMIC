module fake_jpeg_29643_n_389 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_389);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_389;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_SL g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_19),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_27),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_54),
.B(n_81),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_35),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_58),
.A2(n_25),
.B1(n_49),
.B2(n_47),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_33),
.B(n_21),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_28),
.Y(n_84)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_33),
.B(n_20),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_42),
.Y(n_89)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_30),
.B(n_1),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_56),
.A2(n_30),
.B1(n_49),
.B2(n_48),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_83),
.B(n_92),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_95),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_89),
.B(n_107),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_35),
.B1(n_48),
.B2(n_47),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_90),
.A2(n_102),
.B1(n_65),
.B2(n_79),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_35),
.C(n_51),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_26),
.C(n_46),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_68),
.A2(n_38),
.B1(n_30),
.B2(n_34),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_105),
.B(n_40),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_59),
.A2(n_34),
.B1(n_36),
.B2(n_32),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_106),
.A2(n_36),
.B1(n_57),
.B2(n_62),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_42),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_32),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_117),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_L g117 ( 
.A1(n_52),
.A2(n_40),
.B(n_51),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_70),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_61),
.Y(n_135)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_125),
.Y(n_162)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_129),
.Y(n_180)
);

OAI22x1_ASAP7_75t_L g170 ( 
.A1(n_131),
.A2(n_136),
.B1(n_144),
.B2(n_120),
.Y(n_170)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_135),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_69),
.B1(n_71),
.B2(n_53),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_147),
.B1(n_120),
.B2(n_55),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_115),
.A2(n_63),
.B1(n_46),
.B2(n_44),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_137),
.A2(n_142),
.B1(n_156),
.B2(n_115),
.Y(n_161)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_141),
.Y(n_164)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_25),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_146),
.Y(n_169)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_148),
.Y(n_176)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_151),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_85),
.B(n_44),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_24),
.C(n_99),
.Y(n_168)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_86),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_153),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_89),
.B(n_41),
.Y(n_153)
);

AOI32xp33_ASAP7_75t_L g155 ( 
.A1(n_113),
.A2(n_41),
.A3(n_26),
.B1(n_29),
.B2(n_31),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_155),
.B(n_31),
.Y(n_165)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_157),
.A2(n_119),
.B1(n_122),
.B2(n_112),
.Y(n_181)
);

AOI222xp33_ASAP7_75t_L g159 ( 
.A1(n_130),
.A2(n_109),
.B1(n_82),
.B2(n_102),
.C1(n_106),
.C2(n_74),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_159),
.A2(n_167),
.B(n_145),
.C(n_37),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_165),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_24),
.B(n_29),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_174),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_170),
.A2(n_159),
.B1(n_177),
.B2(n_174),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_128),
.B(n_3),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_171),
.B(n_4),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_111),
.B1(n_110),
.B2(n_98),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_101),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_140),
.C(n_154),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_139),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_164),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_183),
.B(n_184),
.Y(n_201)
);

AOI22x1_ASAP7_75t_SL g185 ( 
.A1(n_170),
.A2(n_151),
.B1(n_134),
.B2(n_126),
.Y(n_185)
);

INVxp33_ASAP7_75t_SL g204 ( 
.A(n_185),
.Y(n_204)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_197),
.B1(n_190),
.B2(n_194),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_189),
.B(n_190),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_158),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_198),
.B(n_179),
.Y(n_216)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_160),
.Y(n_200)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_187),
.A2(n_158),
.B(n_165),
.Y(n_203)
);

A2O1A1Ixp33_ASAP7_75t_SL g227 ( 
.A1(n_203),
.A2(n_211),
.B(n_217),
.C(n_184),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_195),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_183),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_182),
.A2(n_170),
.B(n_167),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_185),
.A2(n_163),
.B1(n_169),
.B2(n_168),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_212),
.A2(n_215),
.B1(n_220),
.B2(n_186),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_185),
.A2(n_177),
.B1(n_169),
.B2(n_179),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_162),
.B1(n_180),
.B2(n_176),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_198),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_194),
.A2(n_177),
.B(n_175),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_188),
.A2(n_181),
.B1(n_110),
.B2(n_98),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_221),
.A2(n_209),
.B1(n_208),
.B2(n_210),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_222),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_223),
.B(n_232),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_206),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_224),
.Y(n_256)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_204),
.A2(n_189),
.B1(n_188),
.B2(n_199),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_226),
.A2(n_231),
.B(n_180),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_219),
.Y(n_249)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

AND2x2_ASAP7_75t_SL g230 ( 
.A(n_205),
.B(n_217),
.Y(n_230)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_230),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_211),
.A2(n_175),
.B(n_197),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_171),
.Y(n_232)
);

NOR2xp67_ASAP7_75t_R g233 ( 
.A(n_203),
.B(n_196),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_233),
.B(n_241),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_173),
.C(n_166),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_235),
.C(n_236),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_193),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_192),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_213),
.Y(n_237)
);

BUFx5_ASAP7_75t_L g247 ( 
.A(n_237),
.Y(n_247)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_242),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_239),
.A2(n_209),
.B1(n_208),
.B2(n_210),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_191),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_132),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_176),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_172),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_244),
.A2(n_255),
.B1(n_228),
.B2(n_243),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_246),
.A2(n_248),
.B1(n_262),
.B2(n_229),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_219),
.B1(n_200),
.B2(n_160),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_249),
.B(n_259),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_250),
.A2(n_254),
.B(n_260),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_172),
.C(n_129),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_236),
.C(n_240),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_231),
.A2(n_172),
.B(n_180),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_239),
.A2(n_200),
.B1(n_160),
.B2(n_133),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_180),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_226),
.A2(n_142),
.B1(n_94),
.B2(n_67),
.Y(n_262)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_263),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_253),
.A2(n_250),
.B1(n_254),
.B2(n_222),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_265),
.A2(n_271),
.B1(n_99),
.B2(n_87),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_249),
.A2(n_224),
.B(n_234),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_266),
.B(n_270),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_264),
.B(n_225),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_275),
.Y(n_291)
);

INVx13_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

BUFx12f_ASAP7_75t_L g295 ( 
.A(n_268),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_230),
.B(n_241),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_288),
.C(n_289),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_238),
.Y(n_274)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_257),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_276),
.A2(n_282),
.B1(n_255),
.B2(n_244),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_230),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_280),
.Y(n_300)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_278),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_227),
.Y(n_279)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_247),
.B(n_261),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_257),
.A2(n_227),
.B(n_146),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_281),
.B(n_284),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_248),
.A2(n_227),
.B1(n_94),
.B2(n_125),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_283),
.Y(n_307)
);

NOR3xp33_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_227),
.C(n_141),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_251),
.Y(n_286)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_286),
.Y(n_309)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_258),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_287),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_245),
.B(n_127),
.C(n_138),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_245),
.B(n_252),
.C(n_259),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_290),
.A2(n_271),
.B1(n_302),
.B2(n_294),
.Y(n_314)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_293),
.Y(n_312)
);

NAND4xp25_ASAP7_75t_SL g296 ( 
.A(n_268),
.B(n_148),
.C(n_149),
.D(n_152),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_296),
.B(n_287),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_246),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_303),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_262),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_273),
.B(n_263),
.C(n_258),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_279),
.C(n_288),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_305),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_265),
.A2(n_114),
.B1(n_104),
.B2(n_75),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_308),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_266),
.B(n_114),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_285),
.Y(n_315)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_300),
.Y(n_313)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_313),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_314),
.A2(n_282),
.B1(n_305),
.B2(n_276),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_315),
.B(n_308),
.Y(n_341)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_292),
.Y(n_316)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_316),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_317),
.B(n_319),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_281),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_299),
.Y(n_320)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_320),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_291),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_325),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_298),
.B(n_283),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_303),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_304),
.B(n_270),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_309),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_328),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_301),
.A2(n_307),
.B(n_310),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_327),
.A2(n_311),
.B(n_278),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_297),
.C(n_318),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_329),
.B(n_332),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_331),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_334),
.B(n_341),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_324),
.B(n_290),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_338),
.B(n_321),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_315),
.B(n_269),
.C(n_306),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_339),
.B(n_312),
.C(n_323),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_330),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_343),
.B(n_346),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_344),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_333),
.A2(n_323),
.B1(n_295),
.B2(n_321),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_345),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_338),
.A2(n_269),
.B(n_286),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_349),
.A2(n_5),
.B(n_6),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_336),
.B(n_337),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_350),
.B(n_351),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_341),
.A2(n_272),
.B1(n_296),
.B2(n_295),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_329),
.A2(n_295),
.B(n_87),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_352),
.A2(n_5),
.B(n_6),
.Y(n_363)
);

INVx11_ASAP7_75t_L g353 ( 
.A(n_335),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_353),
.B(n_5),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_343),
.B(n_339),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_355),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_348),
.A2(n_340),
.B1(n_334),
.B2(n_66),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_347),
.B(n_4),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_360),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_345),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_361),
.B(n_7),
.Y(n_368)
);

NAND3xp33_ASAP7_75t_L g370 ( 
.A(n_362),
.B(n_9),
.C(n_10),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_363),
.B(n_364),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_342),
.B(n_7),
.C(n_8),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_365),
.B(n_353),
.C(n_349),
.Y(n_366)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_366),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_368),
.B(n_370),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_359),
.A2(n_10),
.B(n_12),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_372),
.B(n_373),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_356),
.A2(n_14),
.B(n_15),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_369),
.B(n_358),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_376),
.A2(n_15),
.B(n_17),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_367),
.A2(n_364),
.B1(n_358),
.B2(n_16),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_378),
.B(n_379),
.C(n_14),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_371),
.B(n_37),
.C(n_15),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_380),
.Y(n_384)
);

AO21x1_ASAP7_75t_L g383 ( 
.A1(n_381),
.A2(n_382),
.B(n_375),
.Y(n_383)
);

AO21x1_ASAP7_75t_L g382 ( 
.A1(n_377),
.A2(n_17),
.B(n_18),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_383),
.A2(n_374),
.B(n_379),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_385),
.A2(n_384),
.B(n_18),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_386),
.B(n_17),
.C(n_19),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_387),
.A2(n_37),
.B(n_386),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_388),
.B(n_37),
.Y(n_389)
);


endmodule