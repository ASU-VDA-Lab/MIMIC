module fake_netlist_1_7894_n_737 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_737);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_737;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g82 ( .A(n_26), .Y(n_82) );
BUFx3_ASAP7_75t_L g83 ( .A(n_43), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_64), .Y(n_84) );
BUFx2_ASAP7_75t_SL g85 ( .A(n_80), .Y(n_85) );
HB1xp67_ASAP7_75t_L g86 ( .A(n_0), .Y(n_86) );
INVx1_ASAP7_75t_SL g87 ( .A(n_30), .Y(n_87) );
CKINVDCx20_ASAP7_75t_R g88 ( .A(n_77), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_36), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_14), .Y(n_90) );
INVxp67_ASAP7_75t_L g91 ( .A(n_9), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_41), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_45), .Y(n_93) );
INVxp67_ASAP7_75t_SL g94 ( .A(n_24), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_22), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_46), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_78), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_34), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_67), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_61), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_56), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_18), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_69), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_60), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_32), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_72), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_35), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_55), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_20), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_71), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_44), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_57), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_33), .Y(n_113) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_1), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_25), .Y(n_115) );
INVxp33_ASAP7_75t_L g116 ( .A(n_79), .Y(n_116) );
INVxp33_ASAP7_75t_L g117 ( .A(n_76), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_31), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_37), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_11), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_1), .Y(n_121) );
INVx1_ASAP7_75t_SL g122 ( .A(n_23), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_74), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_52), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_27), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_38), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_39), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_5), .Y(n_128) );
INVxp33_ASAP7_75t_L g129 ( .A(n_59), .Y(n_129) );
INVxp67_ASAP7_75t_L g130 ( .A(n_62), .Y(n_130) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_51), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_86), .B(n_0), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_121), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_92), .Y(n_134) );
BUFx2_ASAP7_75t_L g135 ( .A(n_114), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_92), .Y(n_136) );
OA21x2_ASAP7_75t_L g137 ( .A1(n_93), .A2(n_28), .B(n_75), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_131), .B(n_2), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_99), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_93), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_96), .Y(n_141) );
CKINVDCx16_ASAP7_75t_R g142 ( .A(n_88), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_116), .B(n_2), .Y(n_143) );
AOI22x1_ASAP7_75t_L g144 ( .A1(n_99), .A2(n_103), .B1(n_89), .B2(n_123), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_91), .B(n_3), .Y(n_145) );
INVxp67_ASAP7_75t_L g146 ( .A(n_90), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_99), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_121), .Y(n_148) );
INVx6_ASAP7_75t_L g149 ( .A(n_83), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_82), .Y(n_150) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_90), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_82), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_82), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_96), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_97), .B(n_3), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_89), .B(n_4), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_82), .B(n_4), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_97), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_83), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_82), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_83), .B(n_5), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_82), .Y(n_162) );
NOR2xp67_ASAP7_75t_L g163 ( .A(n_130), .B(n_6), .Y(n_163) );
OAI22xp5_ASAP7_75t_L g164 ( .A1(n_120), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_120), .B(n_7), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_95), .Y(n_166) );
BUFx12f_ASAP7_75t_L g167 ( .A(n_106), .Y(n_167) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_128), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_98), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_98), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_100), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_95), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_115), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_100), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_101), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_101), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_165), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_165), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_135), .B(n_129), .Y(n_179) );
AO22x2_ASAP7_75t_L g180 ( .A1(n_161), .A2(n_128), .B1(n_85), .B2(n_124), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_139), .Y(n_181) );
AND2x2_ASAP7_75t_SL g182 ( .A(n_165), .B(n_127), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_135), .A2(n_117), .B1(n_84), .B2(n_94), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_161), .B(n_123), .Y(n_184) );
INVx2_ASAP7_75t_SL g185 ( .A(n_161), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_161), .B(n_103), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_139), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_165), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_176), .Y(n_189) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_143), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_146), .B(n_111), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_151), .B(n_127), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_168), .B(n_85), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_176), .Y(n_194) );
AND2x6_ASAP7_75t_L g195 ( .A(n_159), .B(n_102), .Y(n_195) );
NOR2xp33_ASAP7_75t_SL g196 ( .A(n_167), .B(n_126), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_139), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_176), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_134), .B(n_110), .Y(n_199) );
INVx3_ASAP7_75t_L g200 ( .A(n_176), .Y(n_200) );
BUFx3_ASAP7_75t_L g201 ( .A(n_149), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_134), .B(n_110), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_136), .B(n_109), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_143), .B(n_112), .Y(n_204) );
INVx6_ASAP7_75t_L g205 ( .A(n_167), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_147), .Y(n_206) );
CKINVDCx6p67_ASAP7_75t_R g207 ( .A(n_167), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_136), .Y(n_208) );
XNOR2x2_ASAP7_75t_SL g209 ( .A(n_173), .B(n_102), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_140), .Y(n_210) );
NAND2x1p5_ASAP7_75t_L g211 ( .A(n_140), .B(n_109), .Y(n_211) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_132), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_142), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_141), .B(n_125), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_141), .B(n_119), .Y(n_215) );
INVx1_ASAP7_75t_SL g216 ( .A(n_142), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_159), .B(n_124), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_154), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_154), .B(n_107), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_158), .Y(n_220) );
INVxp67_ASAP7_75t_SL g221 ( .A(n_159), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_158), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_169), .B(n_107), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_169), .B(n_118), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_175), .B(n_118), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_170), .B(n_113), .Y(n_226) );
BUFx10_ASAP7_75t_L g227 ( .A(n_138), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_170), .B(n_113), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_171), .B(n_108), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_150), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_171), .B(n_108), .Y(n_231) );
BUFx6f_ASAP7_75t_SL g232 ( .A(n_174), .Y(n_232) );
INVx4_ASAP7_75t_L g233 ( .A(n_159), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_174), .B(n_105), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_175), .B(n_105), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_133), .B(n_104), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_166), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_145), .Y(n_238) );
OR2x2_ASAP7_75t_L g239 ( .A(n_133), .B(n_104), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_147), .Y(n_240) );
INVxp33_ASAP7_75t_L g241 ( .A(n_163), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_241), .B(n_156), .Y(n_242) );
BUFx3_ASAP7_75t_L g243 ( .A(n_201), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_200), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_207), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_192), .B(n_163), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_200), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_200), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_211), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_179), .B(n_148), .Y(n_250) );
BUFx2_ASAP7_75t_L g251 ( .A(n_207), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_233), .Y(n_252) );
NOR2x1p5_ASAP7_75t_L g253 ( .A(n_213), .B(n_148), .Y(n_253) );
INVx3_ASAP7_75t_L g254 ( .A(n_232), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_211), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_239), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_182), .A2(n_155), .B1(n_164), .B2(n_157), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_233), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_193), .B(n_192), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_233), .Y(n_260) );
BUFx3_ASAP7_75t_L g261 ( .A(n_201), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_213), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_189), .Y(n_263) );
O2A1O1Ixp5_ASAP7_75t_L g264 ( .A1(n_184), .A2(n_172), .B(n_166), .C(n_147), .Y(n_264) );
INVx2_ASAP7_75t_SL g265 ( .A(n_205), .Y(n_265) );
AO22x2_ASAP7_75t_L g266 ( .A1(n_209), .A2(n_172), .B1(n_166), .B2(n_148), .Y(n_266) );
INVx1_ASAP7_75t_SL g267 ( .A(n_216), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_180), .A2(n_144), .B1(n_172), .B2(n_133), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_182), .B(n_144), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_194), .Y(n_270) );
O2A1O1Ixp5_ASAP7_75t_L g271 ( .A1(n_184), .A2(n_133), .B(n_148), .C(n_152), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_198), .Y(n_272) );
A2O1A1Ixp33_ASAP7_75t_L g273 ( .A1(n_177), .A2(n_160), .B(n_152), .C(n_122), .Y(n_273) );
OR2x2_ASAP7_75t_L g274 ( .A(n_212), .B(n_193), .Y(n_274) );
OAI22xp5_ASAP7_75t_L g275 ( .A1(n_178), .A2(n_149), .B1(n_87), .B2(n_137), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_192), .B(n_149), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_191), .B(n_149), .Y(n_277) );
AOI22xp5_ASAP7_75t_L g278 ( .A1(n_180), .A2(n_149), .B1(n_137), .B2(n_152), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_190), .B(n_137), .Y(n_279) );
INVx5_ASAP7_75t_L g280 ( .A(n_195), .Y(n_280) );
INVx2_ASAP7_75t_SL g281 ( .A(n_205), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_199), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_199), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_199), .B(n_137), .Y(n_284) );
BUFx12f_ASAP7_75t_L g285 ( .A(n_205), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_188), .B(n_162), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_185), .B(n_162), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_238), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_181), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_203), .B(n_160), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g291 ( .A1(n_180), .A2(n_160), .B1(n_153), .B2(n_150), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_185), .B(n_162), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_181), .Y(n_293) );
BUFx6f_ASAP7_75t_L g294 ( .A(n_195), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_187), .Y(n_295) );
INVx2_ASAP7_75t_SL g296 ( .A(n_203), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_203), .B(n_225), .Y(n_297) );
BUFx3_ASAP7_75t_L g298 ( .A(n_195), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_225), .Y(n_299) );
INVxp67_ASAP7_75t_L g300 ( .A(n_204), .Y(n_300) );
INVx5_ASAP7_75t_L g301 ( .A(n_195), .Y(n_301) );
INVx2_ASAP7_75t_SL g302 ( .A(n_225), .Y(n_302) );
NOR2xp33_ASAP7_75t_R g303 ( .A(n_232), .B(n_196), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g304 ( .A1(n_208), .A2(n_162), .B1(n_153), .B2(n_150), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_241), .B(n_48), .Y(n_305) );
INVx2_ASAP7_75t_SL g306 ( .A(n_238), .Y(n_306) );
NOR3xp33_ASAP7_75t_SL g307 ( .A(n_224), .B(n_8), .C(n_9), .Y(n_307) );
NAND2xp33_ASAP7_75t_L g308 ( .A(n_195), .B(n_162), .Y(n_308) );
AND2x6_ASAP7_75t_L g309 ( .A(n_217), .B(n_162), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_210), .B(n_153), .Y(n_310) );
INVx3_ASAP7_75t_L g311 ( .A(n_232), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_256), .B(n_222), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_274), .B(n_227), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_282), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_284), .A2(n_186), .B(n_221), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_247), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_283), .Y(n_317) );
NOR2x1_ASAP7_75t_L g318 ( .A(n_251), .B(n_215), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_247), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_259), .A2(n_183), .B1(n_227), .B2(n_220), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g321 ( .A1(n_259), .A2(n_227), .B1(n_218), .B2(n_186), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_269), .A2(n_214), .B(n_202), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_299), .Y(n_323) );
INVx5_ASAP7_75t_L g324 ( .A(n_294), .Y(n_324) );
NAND2xp5_ASAP7_75t_R g325 ( .A(n_306), .B(n_226), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_296), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_302), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_285), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_300), .A2(n_226), .B1(n_228), .B2(n_195), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_289), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_297), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_289), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_263), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_272), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_268), .A2(n_223), .B1(n_228), .B2(n_229), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_254), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_250), .Y(n_337) );
INVx4_ASAP7_75t_L g338 ( .A(n_285), .Y(n_338) );
CKINVDCx16_ASAP7_75t_R g339 ( .A(n_267), .Y(n_339) );
A2O1A1Ixp33_ASAP7_75t_L g340 ( .A1(n_279), .A2(n_234), .B(n_202), .C(n_231), .Y(n_340) );
A2O1A1Ixp33_ASAP7_75t_L g341 ( .A1(n_242), .A2(n_219), .B(n_231), .C(n_235), .Y(n_341) );
INVx3_ASAP7_75t_L g342 ( .A(n_254), .Y(n_342) );
INVx3_ASAP7_75t_L g343 ( .A(n_311), .Y(n_343) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_294), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_293), .Y(n_345) );
INVxp67_ASAP7_75t_L g346 ( .A(n_249), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_266), .A2(n_219), .B1(n_235), .B2(n_240), .Y(n_347) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_288), .A2(n_237), .B1(n_236), .B2(n_240), .Y(n_348) );
INVx2_ASAP7_75t_SL g349 ( .A(n_255), .Y(n_349) );
BUFx2_ASAP7_75t_L g350 ( .A(n_266), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_276), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_270), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_266), .Y(n_353) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_242), .A2(n_240), .B1(n_206), .B2(n_197), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_293), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_294), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_269), .A2(n_206), .B(n_197), .Y(n_357) );
AND2x4_ASAP7_75t_L g358 ( .A(n_311), .B(n_253), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_268), .A2(n_187), .B1(n_153), .B2(n_150), .Y(n_359) );
OR2x6_ASAP7_75t_L g360 ( .A(n_265), .B(n_150), .Y(n_360) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_294), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_291), .A2(n_150), .B1(n_153), .B2(n_12), .Y(n_362) );
AOI21x1_ASAP7_75t_L g363 ( .A1(n_275), .A2(n_230), .B(n_153), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_257), .B(n_10), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_309), .A2(n_230), .B1(n_11), .B2(n_12), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_270), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_339), .B(n_262), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_331), .B(n_295), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_333), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_313), .B(n_245), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_363), .A2(n_278), .B(n_264), .Y(n_371) );
O2A1O1Ixp33_ASAP7_75t_L g372 ( .A1(n_364), .A2(n_246), .B(n_273), .C(n_307), .Y(n_372) );
OAI21x1_ASAP7_75t_L g373 ( .A1(n_357), .A2(n_271), .B(n_310), .Y(n_373) );
BUFx12f_ASAP7_75t_L g374 ( .A(n_338), .Y(n_374) );
AOI22x1_ASAP7_75t_L g375 ( .A1(n_322), .A2(n_295), .B1(n_248), .B2(n_244), .Y(n_375) );
CKINVDCx20_ASAP7_75t_R g376 ( .A(n_328), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_334), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_352), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g379 ( .A1(n_322), .A2(n_287), .B(n_292), .Y(n_379) );
INVx2_ASAP7_75t_SL g380 ( .A(n_324), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_312), .B(n_281), .Y(n_381) );
OAI21x1_ASAP7_75t_L g382 ( .A1(n_357), .A2(n_310), .B(n_287), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_344), .Y(n_383) );
INVx2_ASAP7_75t_SL g384 ( .A(n_324), .Y(n_384) );
OAI21x1_ASAP7_75t_L g385 ( .A1(n_359), .A2(n_292), .B(n_277), .Y(n_385) );
OAI21x1_ASAP7_75t_L g386 ( .A1(n_359), .A2(n_286), .B(n_305), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_366), .Y(n_387) );
OAI21x1_ASAP7_75t_SL g388 ( .A1(n_364), .A2(n_290), .B(n_258), .Y(n_388) );
NAND3xp33_ASAP7_75t_SL g389 ( .A(n_320), .B(n_303), .C(n_273), .Y(n_389) );
INVxp67_ASAP7_75t_L g390 ( .A(n_349), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_315), .A2(n_286), .B(n_258), .Y(n_391) );
OA21x2_ASAP7_75t_L g392 ( .A1(n_347), .A2(n_305), .B(n_304), .Y(n_392) );
AND2x4_ASAP7_75t_L g393 ( .A(n_346), .B(n_298), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_330), .Y(n_394) );
OAI21x1_ASAP7_75t_L g395 ( .A1(n_315), .A2(n_304), .B(n_252), .Y(n_395) );
INVx3_ASAP7_75t_L g396 ( .A(n_324), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_312), .B(n_252), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_332), .Y(n_398) );
OAI21x1_ASAP7_75t_L g399 ( .A1(n_347), .A2(n_260), .B(n_309), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_350), .A2(n_298), .B1(n_280), .B2(n_301), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_345), .Y(n_401) );
OAI22xp33_ASAP7_75t_L g402 ( .A1(n_381), .A2(n_353), .B1(n_329), .B2(n_348), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_368), .B(n_346), .Y(n_403) );
NAND3xp33_ASAP7_75t_L g404 ( .A(n_372), .B(n_365), .C(n_321), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_389), .A2(n_337), .B1(n_351), .B2(n_327), .Y(n_405) );
INVx3_ASAP7_75t_L g406 ( .A(n_396), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_370), .A2(n_327), .B1(n_303), .B2(n_335), .Y(n_407) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_381), .A2(n_318), .B1(n_326), .B2(n_335), .C(n_341), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_369), .A2(n_317), .B1(n_314), .B2(n_323), .C(n_340), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_379), .A2(n_355), .B(n_316), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_367), .A2(n_358), .B1(n_309), .B2(n_336), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_368), .B(n_354), .Y(n_412) );
OAI22xp33_ASAP7_75t_L g413 ( .A1(n_367), .A2(n_397), .B1(n_338), .B2(n_376), .Y(n_413) );
INVx3_ASAP7_75t_L g414 ( .A(n_396), .Y(n_414) );
OAI21xp5_ASAP7_75t_L g415 ( .A1(n_391), .A2(n_362), .B(n_309), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_397), .B(n_319), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_369), .A2(n_358), .B1(n_309), .B2(n_336), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_388), .A2(n_362), .B(n_360), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_377), .A2(n_342), .B1(n_343), .B2(n_365), .Y(n_419) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_377), .A2(n_325), .B1(n_343), .B2(n_342), .C(n_308), .Y(n_420) );
INVx3_ASAP7_75t_L g421 ( .A(n_396), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_378), .A2(n_360), .B1(n_324), .B2(n_361), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_378), .A2(n_360), .B1(n_260), .B2(n_243), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_387), .Y(n_424) );
INVx4_ASAP7_75t_L g425 ( .A(n_396), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_387), .Y(n_426) );
OAI22xp33_ASAP7_75t_L g427 ( .A1(n_390), .A2(n_301), .B1(n_280), .B2(n_344), .Y(n_427) );
AOI222xp33_ASAP7_75t_L g428 ( .A1(n_374), .A2(n_261), .B1(n_243), .B2(n_301), .C1(n_280), .C2(n_344), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_401), .B(n_361), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_401), .B(n_361), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_393), .B(n_261), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_424), .B(n_388), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_416), .B(n_401), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_424), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_416), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_426), .B(n_398), .Y(n_436) );
INVx3_ASAP7_75t_L g437 ( .A(n_425), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_426), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_403), .B(n_398), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_403), .B(n_394), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_429), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_412), .B(n_394), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_429), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_412), .Y(n_444) );
AO21x2_ASAP7_75t_L g445 ( .A1(n_418), .A2(n_371), .B(n_399), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_430), .Y(n_446) );
INVx2_ASAP7_75t_SL g447 ( .A(n_425), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_413), .B(n_374), .Y(n_448) );
NAND2x1p5_ASAP7_75t_SL g449 ( .A(n_430), .B(n_375), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_425), .B(n_380), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_407), .B(n_402), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_406), .Y(n_452) );
INVx5_ASAP7_75t_L g453 ( .A(n_406), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_408), .A2(n_393), .B1(n_392), .B2(n_375), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_406), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_414), .B(n_384), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_414), .B(n_380), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_414), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_421), .B(n_384), .Y(n_459) );
AND2x4_ASAP7_75t_L g460 ( .A(n_421), .B(n_399), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_421), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_431), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_422), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_405), .B(n_393), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_409), .B(n_392), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_423), .Y(n_466) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_404), .Y(n_467) );
BUFx2_ASAP7_75t_L g468 ( .A(n_437), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_435), .B(n_411), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_444), .B(n_415), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_435), .B(n_417), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_433), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_444), .B(n_371), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_446), .B(n_10), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_434), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_460), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_460), .B(n_410), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_446), .B(n_13), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_434), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_438), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_446), .B(n_13), .Y(n_481) );
NAND2x1p5_ASAP7_75t_L g482 ( .A(n_437), .B(n_383), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_442), .B(n_14), .Y(n_483) );
AOI221xp5_ASAP7_75t_L g484 ( .A1(n_451), .A2(n_420), .B1(n_419), .B2(n_393), .C(n_423), .Y(n_484) );
BUFx2_ASAP7_75t_L g485 ( .A(n_437), .Y(n_485) );
OAI31xp33_ASAP7_75t_L g486 ( .A1(n_448), .A2(n_427), .A3(n_400), .B(n_383), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_438), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_432), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_442), .B(n_15), .Y(n_489) );
BUFx2_ASAP7_75t_L g490 ( .A(n_437), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_432), .Y(n_491) );
OAI221xp5_ASAP7_75t_L g492 ( .A1(n_454), .A2(n_464), .B1(n_467), .B2(n_463), .C(n_450), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_436), .Y(n_493) );
BUFx2_ASAP7_75t_L g494 ( .A(n_447), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_442), .A2(n_392), .B1(n_386), .B2(n_428), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_443), .B(n_15), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_460), .Y(n_497) );
OA332x1_ASAP7_75t_L g498 ( .A1(n_439), .A2(n_16), .A3(n_17), .B1(n_440), .B2(n_467), .B3(n_464), .C1(n_449), .C2(n_443), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_460), .B(n_383), .Y(n_499) );
AND2x4_ASAP7_75t_L g500 ( .A(n_458), .B(n_382), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_433), .B(n_16), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_439), .A2(n_392), .B1(n_386), .B2(n_385), .Y(n_502) );
AOI221xp5_ASAP7_75t_L g503 ( .A1(n_467), .A2(n_230), .B1(n_17), .B2(n_356), .C(n_301), .Y(n_503) );
INVx3_ASAP7_75t_L g504 ( .A(n_447), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_441), .B(n_395), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_441), .B(n_395), .Y(n_506) );
INVx4_ASAP7_75t_L g507 ( .A(n_453), .Y(n_507) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_439), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_440), .B(n_373), .Y(n_509) );
NOR2xp67_ASAP7_75t_L g510 ( .A(n_447), .B(n_19), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_453), .B(n_356), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_440), .B(n_373), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_441), .B(n_382), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_436), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_462), .B(n_385), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_445), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_436), .B(n_21), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_462), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_509), .B(n_512), .Y(n_519) );
NOR3xp33_ASAP7_75t_L g520 ( .A(n_501), .B(n_459), .C(n_456), .Y(n_520) );
AOI22xp33_ASAP7_75t_SL g521 ( .A1(n_494), .A2(n_463), .B1(n_453), .B2(n_456), .Y(n_521) );
INVx3_ASAP7_75t_L g522 ( .A(n_507), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_475), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_475), .Y(n_524) );
INVxp67_ASAP7_75t_SL g525 ( .A(n_494), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_509), .B(n_445), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_507), .B(n_504), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_512), .B(n_445), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_473), .B(n_445), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_479), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_472), .B(n_462), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_473), .B(n_466), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_470), .B(n_466), .Y(n_533) );
AOI221xp5_ASAP7_75t_L g534 ( .A1(n_492), .A2(n_467), .B1(n_465), .B2(n_455), .C(n_461), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_470), .B(n_466), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_508), .B(n_452), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_468), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_513), .B(n_467), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_483), .B(n_452), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_483), .B(n_461), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_516), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_488), .B(n_465), .Y(n_542) );
NOR2x1p5_ASAP7_75t_L g543 ( .A(n_507), .B(n_450), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_516), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_513), .B(n_467), .Y(n_545) );
AND2x4_ASAP7_75t_L g546 ( .A(n_476), .B(n_458), .Y(n_546) );
BUFx2_ASAP7_75t_L g547 ( .A(n_468), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_488), .B(n_458), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_491), .B(n_455), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_516), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_489), .B(n_459), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_479), .Y(n_552) );
OAI21xp5_ASAP7_75t_SL g553 ( .A1(n_498), .A2(n_457), .B(n_453), .Y(n_553) );
OAI21xp5_ASAP7_75t_L g554 ( .A1(n_510), .A2(n_501), .B(n_489), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_493), .B(n_457), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_518), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_480), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_491), .B(n_453), .Y(n_558) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_485), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_480), .Y(n_560) );
AND3x1_ASAP7_75t_L g561 ( .A(n_504), .B(n_453), .C(n_449), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_493), .B(n_453), .Y(n_562) );
AND2x4_ASAP7_75t_SL g563 ( .A(n_507), .B(n_449), .Y(n_563) );
INVx3_ASAP7_75t_L g564 ( .A(n_504), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_514), .B(n_29), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_487), .Y(n_566) );
AOI31xp33_ASAP7_75t_SL g567 ( .A1(n_496), .A2(n_40), .A3(n_42), .B(n_47), .Y(n_567) );
BUFx2_ASAP7_75t_L g568 ( .A(n_485), .Y(n_568) );
INVxp67_ASAP7_75t_R g569 ( .A(n_517), .Y(n_569) );
AOI211x1_ASAP7_75t_SL g570 ( .A1(n_469), .A2(n_230), .B(n_50), .C(n_53), .Y(n_570) );
NOR2x1_ASAP7_75t_R g571 ( .A(n_490), .B(n_504), .Y(n_571) );
NOR2xp67_ASAP7_75t_L g572 ( .A(n_510), .B(n_49), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_518), .Y(n_573) );
OAI21xp5_ASAP7_75t_SL g574 ( .A1(n_490), .A2(n_356), .B(n_58), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_514), .B(n_54), .Y(n_575) );
INVx3_ASAP7_75t_L g576 ( .A(n_477), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_487), .Y(n_577) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_474), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_519), .B(n_474), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_519), .B(n_481), .Y(n_580) );
INVx2_ASAP7_75t_SL g581 ( .A(n_543), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_541), .Y(n_582) );
NOR2x1_ASAP7_75t_L g583 ( .A(n_574), .B(n_496), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_523), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_569), .B(n_499), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_523), .Y(n_586) );
INVxp67_ASAP7_75t_L g587 ( .A(n_547), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_524), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_524), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_569), .B(n_499), .Y(n_590) );
AND2x4_ASAP7_75t_L g591 ( .A(n_543), .B(n_476), .Y(n_591) );
OR2x6_ASAP7_75t_L g592 ( .A(n_554), .B(n_497), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_547), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_530), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_530), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_578), .B(n_562), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_520), .B(n_478), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_531), .B(n_497), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_549), .B(n_478), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_549), .B(n_481), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_552), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_552), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_551), .B(n_497), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_541), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_557), .B(n_471), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_557), .B(n_505), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_541), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_560), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_544), .Y(n_609) );
AOI21xp33_ASAP7_75t_L g610 ( .A1(n_553), .A2(n_486), .B(n_517), .Y(n_610) );
NAND3xp33_ASAP7_75t_L g611 ( .A(n_534), .B(n_486), .C(n_484), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_560), .B(n_505), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_562), .B(n_499), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_542), .B(n_539), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_566), .B(n_506), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_533), .B(n_499), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_544), .Y(n_617) );
AND2x4_ASAP7_75t_SL g618 ( .A(n_522), .B(n_476), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_542), .B(n_506), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_536), .B(n_515), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_540), .B(n_515), .Y(n_621) );
INVx2_ASAP7_75t_SL g622 ( .A(n_522), .Y(n_622) );
INVxp67_ASAP7_75t_L g623 ( .A(n_568), .Y(n_623) );
INVx1_ASAP7_75t_SL g624 ( .A(n_568), .Y(n_624) );
NOR4xp25_ASAP7_75t_L g625 ( .A(n_567), .B(n_495), .C(n_502), .D(n_503), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_566), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_544), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_577), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_577), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_556), .Y(n_630) );
BUFx2_ASAP7_75t_L g631 ( .A(n_571), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_533), .B(n_477), .Y(n_632) );
AND2x4_ASAP7_75t_L g633 ( .A(n_576), .B(n_477), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_596), .B(n_526), .Y(n_634) );
OAI22xp33_ASAP7_75t_L g635 ( .A1(n_597), .A2(n_522), .B1(n_525), .B2(n_537), .Y(n_635) );
NOR2xp33_ASAP7_75t_SL g636 ( .A(n_581), .B(n_571), .Y(n_636) );
OAI21xp33_ASAP7_75t_L g637 ( .A1(n_625), .A2(n_583), .B(n_610), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_582), .Y(n_638) );
AOI222xp33_ASAP7_75t_L g639 ( .A1(n_611), .A2(n_526), .B1(n_528), .B2(n_529), .C1(n_555), .C2(n_535), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_584), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_586), .Y(n_641) );
AOI211xp5_ASAP7_75t_SL g642 ( .A1(n_587), .A2(n_522), .B(n_572), .C(n_559), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_616), .B(n_528), .Y(n_643) );
INVx1_ASAP7_75t_SL g644 ( .A(n_593), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_588), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_589), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_594), .Y(n_647) );
INVxp67_ASAP7_75t_L g648 ( .A(n_614), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_595), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_632), .B(n_545), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_614), .B(n_529), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_601), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_582), .Y(n_653) );
AOI32xp33_ASAP7_75t_L g654 ( .A1(n_581), .A2(n_561), .A3(n_521), .B1(n_563), .B2(n_576), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_602), .Y(n_655) );
O2A1O1Ixp33_ASAP7_75t_L g656 ( .A1(n_587), .A2(n_527), .B(n_575), .C(n_565), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_624), .B(n_564), .Y(n_657) );
OAI21xp33_ASAP7_75t_L g658 ( .A1(n_592), .A2(n_563), .B(n_576), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_619), .B(n_535), .Y(n_659) );
INVxp67_ASAP7_75t_L g660 ( .A(n_622), .Y(n_660) );
O2A1O1Ixp33_ASAP7_75t_L g661 ( .A1(n_623), .A2(n_575), .B(n_565), .C(n_576), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_608), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_613), .B(n_538), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_592), .A2(n_561), .B1(n_572), .B2(n_563), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_592), .A2(n_558), .B1(n_538), .B2(n_545), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_631), .A2(n_558), .B1(n_477), .B2(n_548), .Y(n_666) );
OAI21xp5_ASAP7_75t_SL g667 ( .A1(n_585), .A2(n_570), .B(n_564), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_604), .Y(n_668) );
OAI22xp33_ASAP7_75t_L g669 ( .A1(n_579), .A2(n_564), .B1(n_573), .B2(n_556), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_590), .B(n_532), .Y(n_670) );
AND2x4_ASAP7_75t_L g671 ( .A(n_622), .B(n_564), .Y(n_671) );
NOR2xp33_ASAP7_75t_R g672 ( .A(n_591), .B(n_548), .Y(n_672) );
OAI21xp33_ASAP7_75t_L g673 ( .A1(n_637), .A2(n_623), .B(n_619), .Y(n_673) );
XNOR2xp5_ASAP7_75t_L g674 ( .A(n_644), .B(n_580), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_665), .A2(n_591), .B1(n_603), .B2(n_618), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_640), .Y(n_676) );
OAI221xp5_ASAP7_75t_L g677 ( .A1(n_654), .A2(n_605), .B1(n_620), .B2(n_621), .C(n_598), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_665), .A2(n_591), .B1(n_600), .B2(n_599), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_639), .B(n_629), .Y(n_679) );
NAND5xp2_ASAP7_75t_L g680 ( .A(n_636), .B(n_482), .C(n_532), .D(n_628), .E(n_626), .Y(n_680) );
INVx1_ASAP7_75t_SL g681 ( .A(n_672), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_648), .A2(n_618), .B1(n_633), .B2(n_630), .Y(n_682) );
A2O1A1Ixp33_ASAP7_75t_L g683 ( .A1(n_658), .A2(n_633), .B(n_615), .C(n_556), .Y(n_683) );
INVxp67_ASAP7_75t_SL g684 ( .A(n_635), .Y(n_684) );
NOR2x1_ASAP7_75t_L g685 ( .A(n_635), .B(n_633), .Y(n_685) );
OR2x2_ASAP7_75t_L g686 ( .A(n_659), .B(n_606), .Y(n_686) );
OR2x2_ASAP7_75t_L g687 ( .A(n_651), .B(n_612), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g688 ( .A(n_664), .B(n_627), .Y(n_688) );
AOI211xp5_ASAP7_75t_L g689 ( .A1(n_669), .A2(n_627), .B(n_617), .C(n_609), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_641), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_634), .B(n_617), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_666), .A2(n_609), .B1(n_607), .B2(n_604), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_645), .Y(n_693) );
AO22x1_ASAP7_75t_L g694 ( .A1(n_671), .A2(n_573), .B1(n_607), .B2(n_546), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_669), .B(n_573), .Y(n_695) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_672), .Y(n_696) );
NOR2x1_ASAP7_75t_L g697 ( .A(n_656), .B(n_550), .Y(n_697) );
NAND2xp5_ASAP7_75t_SL g698 ( .A(n_685), .B(n_671), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_679), .B(n_643), .Y(n_699) );
NAND2xp33_ASAP7_75t_SL g700 ( .A(n_696), .B(n_666), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_681), .A2(n_642), .B(n_661), .Y(n_701) );
OAI21xp33_ASAP7_75t_SL g702 ( .A1(n_684), .A2(n_660), .B(n_657), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_676), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_690), .Y(n_704) );
A2O1A1Ixp33_ASAP7_75t_L g705 ( .A1(n_673), .A2(n_667), .B(n_657), .C(n_670), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g706 ( .A1(n_694), .A2(n_511), .B(n_653), .Y(n_706) );
AOI22xp5_ASAP7_75t_SL g707 ( .A1(n_680), .A2(n_663), .B1(n_650), .B2(n_662), .Y(n_707) );
O2A1O1Ixp5_ASAP7_75t_SL g708 ( .A1(n_688), .A2(n_647), .B(n_655), .C(n_652), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_693), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g710 ( .A1(n_677), .A2(n_649), .B1(n_646), .B2(n_668), .C(n_653), .Y(n_710) );
NOR2xp67_ASAP7_75t_L g711 ( .A(n_682), .B(n_668), .Y(n_711) );
XNOR2xp5_ASAP7_75t_L g712 ( .A(n_674), .B(n_638), .Y(n_712) );
INVx1_ASAP7_75t_SL g713 ( .A(n_700), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_707), .A2(n_675), .B1(n_683), .B2(n_678), .Y(n_714) );
NAND4xp25_ASAP7_75t_SL g715 ( .A(n_702), .B(n_697), .C(n_689), .D(n_692), .Y(n_715) );
XNOR2x2_ASAP7_75t_L g716 ( .A(n_698), .B(n_682), .Y(n_716) );
AOI211xp5_ASAP7_75t_L g717 ( .A1(n_705), .A2(n_678), .B(n_695), .C(n_687), .Y(n_717) );
AOI221xp5_ASAP7_75t_L g718 ( .A1(n_710), .A2(n_699), .B1(n_701), .B2(n_709), .C(n_703), .Y(n_718) );
AOI211xp5_ASAP7_75t_SL g719 ( .A1(n_711), .A2(n_686), .B(n_691), .C(n_638), .Y(n_719) );
A2O1A1Ixp33_ASAP7_75t_L g720 ( .A1(n_706), .A2(n_546), .B(n_550), .C(n_500), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_704), .Y(n_721) );
BUFx2_ASAP7_75t_L g722 ( .A(n_716), .Y(n_722) );
AND4x1_ASAP7_75t_L g723 ( .A(n_717), .B(n_706), .C(n_570), .D(n_708), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_721), .Y(n_724) );
NOR3xp33_ASAP7_75t_L g725 ( .A(n_715), .B(n_550), .C(n_712), .Y(n_725) );
NAND3xp33_ASAP7_75t_L g726 ( .A(n_718), .B(n_500), .C(n_546), .Y(n_726) );
NOR2x1_ASAP7_75t_L g727 ( .A(n_722), .B(n_713), .Y(n_727) );
OR4x2_ASAP7_75t_L g728 ( .A(n_725), .B(n_720), .C(n_714), .D(n_719), .Y(n_728) );
OR4x2_ASAP7_75t_L g729 ( .A(n_723), .B(n_482), .C(n_546), .D(n_500), .Y(n_729) );
INVx3_ASAP7_75t_L g730 ( .A(n_728), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_727), .B(n_724), .Y(n_731) );
OAI22x1_ASAP7_75t_L g732 ( .A1(n_730), .A2(n_729), .B1(n_726), .B2(n_482), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_731), .Y(n_733) );
AND2x4_ASAP7_75t_L g734 ( .A(n_733), .B(n_500), .Y(n_734) );
AOI222xp33_ASAP7_75t_L g735 ( .A1(n_734), .A2(n_732), .B1(n_280), .B2(n_66), .C1(n_68), .C2(n_63), .Y(n_735) );
OAI22xp33_ASAP7_75t_L g736 ( .A1(n_735), .A2(n_734), .B1(n_70), .B2(n_73), .Y(n_736) );
AOI21xp5_ASAP7_75t_L g737 ( .A1(n_736), .A2(n_65), .B(n_81), .Y(n_737) );
endmodule