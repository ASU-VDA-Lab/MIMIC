module fake_netlist_6_2877_n_453 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_453);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_453;

wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_209;
wire n_367;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_161;
wire n_208;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_350;
wire n_392;
wire n_442;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_443;
wire n_246;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_230;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_372;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_375;
wire n_338;
wire n_360;
wire n_235;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_428;
wire n_432;
wire n_167;
wire n_174;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_294;
wire n_302;
wire n_380;
wire n_197;
wire n_343;
wire n_448;
wire n_397;
wire n_445;
wire n_425;
wire n_218;
wire n_234;
wire n_381;
wire n_236;
wire n_172;
wire n_270;
wire n_239;
wire n_414;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_417;
wire n_446;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_293;
wire n_334;
wire n_370;
wire n_232;
wire n_163;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_321;
wire n_331;
wire n_227;
wire n_406;
wire n_204;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_164;
wire n_292;
wire n_307;
wire n_433;
wire n_291;
wire n_219;
wire n_357;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_282;
wire n_436;
wire n_211;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_240;
wire n_319;
wire n_273;
wire n_311;
wire n_403;
wire n_253;
wire n_249;
wire n_201;
wire n_386;
wire n_159;
wire n_162;
wire n_241;
wire n_275;
wire n_276;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_318;
wire n_303;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_277;
wire n_418;
wire n_199;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_431;
wire n_347;
wire n_328;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_205;
wire n_251;
wire n_301;
wire n_274;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_288;
wire n_427;
wire n_422;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_391;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_187;
wire n_361;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_13),
.B(n_150),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_16),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_34),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_69),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_117),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_12),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_60),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_63),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_67),
.Y(n_168)
);

INVxp33_ASAP7_75t_SL g169 ( 
.A(n_45),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_84),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_36),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_74),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_31),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_92),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_134),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_28),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_151),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_39),
.B(n_5),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_138),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_81),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_38),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_24),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_102),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_42),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_26),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_132),
.Y(n_186)
);

INVxp33_ASAP7_75t_SL g187 ( 
.A(n_20),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_40),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_87),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_68),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_142),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_89),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_147),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_6),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_30),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_7),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_156),
.Y(n_198)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_133),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_1),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_65),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_96),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_18),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_101),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_155),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_93),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_48),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_127),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_104),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_125),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_64),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_91),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_106),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_8),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_76),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_29),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_57),
.B(n_140),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_88),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_32),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_157),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_21),
.Y(n_221)
);

BUFx2_ASAP7_75t_SL g222 ( 
.A(n_44),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_124),
.B(n_43),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_23),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_95),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_54),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_70),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_53),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_2),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_9),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_137),
.Y(n_231)
);

INVxp67_ASAP7_75t_SL g232 ( 
.A(n_58),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_15),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_14),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_62),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_33),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_118),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_46),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_77),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_3),
.Y(n_240)
);

INVxp67_ASAP7_75t_SL g241 ( 
.A(n_139),
.Y(n_241)
);

BUFx6f_ASAP7_75t_SL g242 ( 
.A(n_94),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_25),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_152),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_131),
.B(n_154),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_61),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_113),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_83),
.Y(n_248)
);

NOR2xp67_ASAP7_75t_L g249 ( 
.A(n_116),
.B(n_153),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_51),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_115),
.Y(n_251)
);

INVxp67_ASAP7_75t_SL g252 ( 
.A(n_130),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_97),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_78),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_49),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_86),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_111),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_80),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_103),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_72),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_82),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_50),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_110),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_143),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_27),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_71),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_120),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_85),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_R g269 ( 
.A(n_112),
.B(n_17),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_75),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_121),
.Y(n_271)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_136),
.Y(n_272)
);

INVxp67_ASAP7_75t_SL g273 ( 
.A(n_22),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_4),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_52),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_55),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_119),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_123),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_202),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_196),
.B(n_0),
.Y(n_280)
);

INVxp67_ASAP7_75t_SL g281 ( 
.A(n_182),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_225),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_160),
.Y(n_283)
);

BUFx4f_ASAP7_75t_L g284 ( 
.A(n_159),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_161),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_183),
.B(n_0),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_162),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_163),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_185),
.A2(n_10),
.B1(n_11),
.B2(n_19),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_165),
.Y(n_290)
);

BUFx10_ASAP7_75t_L g291 ( 
.A(n_242),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_220),
.B(n_35),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_238),
.B(n_37),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_214),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_242),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_251),
.B(n_41),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_169),
.B(n_47),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_167),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_164),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_166),
.Y(n_300)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_204),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_187),
.B(n_56),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_176),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_260),
.B(n_262),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_170),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_168),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_171),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_173),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_248),
.B(n_59),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_175),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_244),
.B(n_66),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_188),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_172),
.Y(n_313)
);

AND2x6_ASAP7_75t_L g314 ( 
.A(n_158),
.B(n_73),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_191),
.Y(n_315)
);

AND2x6_ASAP7_75t_L g316 ( 
.A(n_178),
.B(n_79),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_192),
.Y(n_317)
);

AND2x4_ASAP7_75t_L g318 ( 
.A(n_194),
.B(n_90),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_198),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_203),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_210),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_212),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_221),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_174),
.Y(n_324)
);

BUFx10_ASAP7_75t_L g325 ( 
.A(n_223),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_228),
.B(n_98),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_231),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_233),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_236),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_222),
.A2(n_99),
.B1(n_100),
.B2(n_105),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_239),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_240),
.B(n_107),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_250),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_253),
.B(n_108),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_255),
.B(n_109),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_257),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_282),
.B(n_177),
.Y(n_337)
);

NAND2xp33_ASAP7_75t_SL g338 ( 
.A(n_286),
.B(n_190),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_325),
.B(n_179),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_324),
.B(n_259),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_301),
.B(n_180),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_295),
.B(n_181),
.Y(n_342)
);

NAND2xp33_ASAP7_75t_SL g343 ( 
.A(n_296),
.B(n_197),
.Y(n_343)
);

NAND2xp33_ASAP7_75t_SL g344 ( 
.A(n_304),
.B(n_205),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_291),
.B(n_184),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_283),
.B(n_186),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_299),
.B(n_189),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_280),
.B(n_193),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_306),
.B(n_263),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_313),
.B(n_267),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_279),
.B(n_207),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_300),
.B(n_271),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_279),
.B(n_235),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_292),
.B(n_227),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_309),
.B(n_201),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_284),
.B(n_318),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_332),
.B(n_237),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_335),
.B(n_293),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_281),
.B(n_294),
.Y(n_359)
);

NAND2xp33_ASAP7_75t_SL g360 ( 
.A(n_336),
.B(n_229),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_329),
.B(n_275),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_297),
.B(n_226),
.Y(n_362)
);

NAND2xp33_ASAP7_75t_SL g363 ( 
.A(n_330),
.B(n_234),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_331),
.B(n_278),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_302),
.B(n_219),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_326),
.B(n_224),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_285),
.B(n_277),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_334),
.B(n_218),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_305),
.B(n_276),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_311),
.B(n_274),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_305),
.B(n_195),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_307),
.B(n_320),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_308),
.B(n_247),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_341),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_358),
.A2(n_363),
.B1(n_314),
.B2(n_316),
.Y(n_375)
);

OA21x2_ASAP7_75t_L g376 ( 
.A1(n_350),
.A2(n_217),
.B(n_333),
.Y(n_376)
);

OAI21x1_ASAP7_75t_L g377 ( 
.A1(n_356),
.A2(n_289),
.B(n_328),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_373),
.Y(n_378)
);

OAI21x1_ASAP7_75t_L g379 ( 
.A1(n_340),
.A2(n_312),
.B(n_322),
.Y(n_379)
);

BUFx8_ASAP7_75t_SL g380 ( 
.A(n_349),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_355),
.A2(n_314),
.B(n_316),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_367),
.Y(n_382)
);

OAI22xp33_ASAP7_75t_L g383 ( 
.A1(n_361),
.A2(n_364),
.B1(n_339),
.B2(n_258),
.Y(n_383)
);

OAI21x1_ASAP7_75t_L g384 ( 
.A1(n_366),
.A2(n_327),
.B(n_323),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_L g385 ( 
.A1(n_370),
.A2(n_321),
.B1(n_287),
.B2(n_319),
.Y(n_385)
);

AOI22x1_ASAP7_75t_L g386 ( 
.A1(n_338),
.A2(n_288),
.B1(n_317),
.B2(n_315),
.Y(n_386)
);

AO31x2_ASAP7_75t_L g387 ( 
.A1(n_352),
.A2(n_310),
.A3(n_298),
.B(n_290),
.Y(n_387)
);

OAI21x1_ASAP7_75t_L g388 ( 
.A1(n_368),
.A2(n_241),
.B(n_232),
.Y(n_388)
);

OAI21x1_ASAP7_75t_L g389 ( 
.A1(n_354),
.A2(n_252),
.B(n_273),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_357),
.A2(n_199),
.B(n_272),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_359),
.B(n_320),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_372),
.Y(n_392)
);

NAND2x1p5_ASAP7_75t_L g393 ( 
.A(n_346),
.B(n_249),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_369),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_351),
.B(n_266),
.Y(n_395)
);

OA21x2_ASAP7_75t_L g396 ( 
.A1(n_348),
.A2(n_245),
.B(n_270),
.Y(n_396)
);

OAI21x1_ASAP7_75t_L g397 ( 
.A1(n_342),
.A2(n_269),
.B(n_209),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_353),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_371),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_391),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_374),
.B(n_360),
.Y(n_401)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_391),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_380),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_378),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_392),
.B(n_303),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_384),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_378),
.B(n_347),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_R g408 ( 
.A(n_399),
.B(n_344),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_382),
.B(n_365),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_394),
.B(n_345),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_387),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_379),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_376),
.B(n_362),
.Y(n_413)
);

BUFx8_ASAP7_75t_SL g414 ( 
.A(n_395),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_386),
.B(n_337),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_398),
.B(n_206),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_377),
.B(n_216),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_402),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_400),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_404),
.B(n_385),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_411),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_SL g422 ( 
.A1(n_409),
.A2(n_393),
.B1(n_381),
.B2(n_390),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_417),
.B(n_383),
.Y(n_423)
);

OAI31xp33_ASAP7_75t_L g424 ( 
.A1(n_415),
.A2(n_343),
.A3(n_375),
.B(n_261),
.Y(n_424)
);

AO21x2_ASAP7_75t_L g425 ( 
.A1(n_413),
.A2(n_389),
.B(n_388),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_405),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_406),
.Y(n_427)
);

OAI31xp33_ASAP7_75t_SL g428 ( 
.A1(n_422),
.A2(n_407),
.A3(n_410),
.B(n_397),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_423),
.B(n_408),
.Y(n_429)
);

NOR2x1_ASAP7_75t_L g430 ( 
.A(n_426),
.B(n_401),
.Y(n_430)
);

OAI221xp5_ASAP7_75t_L g431 ( 
.A1(n_424),
.A2(n_401),
.B1(n_403),
.B2(n_396),
.C(n_414),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_418),
.B(n_416),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_420),
.B(n_230),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_419),
.B(n_387),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_421),
.B(n_412),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_427),
.B(n_307),
.Y(n_436)
);

NAND3xp33_ASAP7_75t_L g437 ( 
.A(n_433),
.B(n_200),
.C(n_268),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_435),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_429),
.A2(n_427),
.B1(n_246),
.B2(n_265),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_432),
.B(n_430),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_436),
.B(n_425),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_438),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_440),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_439),
.Y(n_444)
);

XNOR2x1_ASAP7_75t_L g445 ( 
.A(n_442),
.B(n_437),
.Y(n_445)
);

AOI322xp5_ASAP7_75t_L g446 ( 
.A1(n_444),
.A2(n_443),
.A3(n_431),
.B1(n_208),
.B2(n_211),
.C1(n_213),
.C2(n_215),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_446),
.B(n_428),
.Y(n_447)
);

NAND2xp33_ASAP7_75t_SL g448 ( 
.A(n_445),
.B(n_434),
.Y(n_448)
);

OAI221xp5_ASAP7_75t_L g449 ( 
.A1(n_448),
.A2(n_264),
.B1(n_256),
.B2(n_254),
.C(n_243),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_447),
.Y(n_450)
);

AOI31xp33_ASAP7_75t_L g451 ( 
.A1(n_450),
.A2(n_449),
.A3(n_441),
.B(n_126),
.Y(n_451)
);

AO221x1_ASAP7_75t_L g452 ( 
.A1(n_451),
.A2(n_114),
.B1(n_122),
.B2(n_129),
.C(n_141),
.Y(n_452)
);

AOI221xp5_ASAP7_75t_L g453 ( 
.A1(n_452),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.C(n_148),
.Y(n_453)
);


endmodule