module fake_netlist_5_853_n_151 (n_29, n_16, n_0, n_12, n_9, n_36, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_40, n_34, n_38, n_4, n_32, n_35, n_41, n_11, n_17, n_19, n_7, n_37, n_15, n_26, n_30, n_20, n_5, n_33, n_14, n_2, n_31, n_23, n_13, n_3, n_6, n_39, n_151);

input n_29;
input n_16;
input n_0;
input n_12;
input n_9;
input n_36;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_40;
input n_34;
input n_38;
input n_4;
input n_32;
input n_35;
input n_41;
input n_11;
input n_17;
input n_19;
input n_7;
input n_37;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_33;
input n_14;
input n_2;
input n_31;
input n_23;
input n_13;
input n_3;
input n_6;
input n_39;

output n_151;

wire n_137;
wire n_91;
wire n_82;
wire n_122;
wire n_142;
wire n_140;
wire n_124;
wire n_86;
wire n_136;
wire n_146;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_111;
wire n_108;
wire n_129;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_123;
wire n_139;
wire n_105;
wire n_80;
wire n_125;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_126;
wire n_84;
wire n_130;
wire n_79;
wire n_131;
wire n_47;
wire n_53;
wire n_44;
wire n_100;
wire n_62;
wire n_138;
wire n_148;
wire n_71;
wire n_109;
wire n_112;
wire n_85;
wire n_95;
wire n_119;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_49;
wire n_54;
wire n_147;
wire n_67;
wire n_121;
wire n_76;
wire n_87;
wire n_150;
wire n_64;
wire n_77;
wire n_102;
wire n_106;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_134;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_97;
wire n_63;
wire n_141;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_16),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_2),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_1),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_58),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_2),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

AOI21x1_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_5),
.B(n_6),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_49),
.Y(n_87)
);

OR2x6_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_68),
.Y(n_88)
);

AND2x4_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_65),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

NAND3xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_49),
.C(n_57),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_81),
.B(n_85),
.C(n_82),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_69),
.B1(n_70),
.B2(n_73),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

AOI31xp67_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_86),
.A3(n_62),
.B(n_73),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_76),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

OAI21x1_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_84),
.B(n_83),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_67),
.B(n_63),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_83),
.Y(n_110)
);

OA21x2_ASAP7_75t_L g111 ( 
.A1(n_107),
.A2(n_100),
.B(n_105),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_109),
.A2(n_54),
.B(n_47),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_98),
.Y(n_114)
);

INVx3_ASAP7_75t_SL g115 ( 
.A(n_101),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_78),
.Y(n_116)
);

AOI31xp33_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_44),
.A3(n_18),
.B(n_19),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_90),
.B1(n_21),
.B2(n_22),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

AND2x4_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_110),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_115),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_90),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_8),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_23),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

NOR2x1_ASAP7_75t_SL g128 ( 
.A(n_119),
.B(n_90),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_27),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_121),
.B(n_117),
.Y(n_131)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

NAND3xp33_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_103),
.C(n_32),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_123),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_SL g137 ( 
.A1(n_131),
.A2(n_122),
.B(n_124),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_135),
.B(n_122),
.Y(n_139)
);

OR2x6_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_136),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_132),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_140),
.A2(n_134),
.B1(n_129),
.B2(n_130),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_141),
.B(n_137),
.Y(n_143)
);

INVxp67_ASAP7_75t_SL g144 ( 
.A(n_142),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_145),
.Y(n_146)
);

OAI221xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_143),
.B1(n_138),
.B2(n_130),
.C(n_37),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_28),
.B(n_33),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_35),
.B1(n_38),
.B2(n_40),
.Y(n_151)
);


endmodule