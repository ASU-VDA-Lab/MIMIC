module real_jpeg_29766_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_70;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_0),
.A2(n_36),
.B1(n_37),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_0),
.A2(n_22),
.B1(n_27),
.B2(n_44),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_0),
.A2(n_44),
.B1(n_67),
.B2(n_68),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_0),
.A2(n_44),
.B1(n_62),
.B2(n_65),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_SL g90 ( 
.A1(n_0),
.A2(n_62),
.B(n_64),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_SL g124 ( 
.A1(n_0),
.A2(n_37),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_0),
.B(n_61),
.Y(n_135)
);

AOI21xp33_ASAP7_75t_L g150 ( 
.A1(n_0),
.A2(n_22),
.B(n_38),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_0),
.B(n_76),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_4),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_6),
.A2(n_22),
.B1(n_27),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_8),
.A2(n_22),
.B1(n_27),
.B2(n_39),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_9),
.A2(n_42),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_9),
.A2(n_22),
.B1(n_27),
.B2(n_42),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_9),
.A2(n_42),
.B1(n_62),
.B2(n_65),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_10),
.A2(n_62),
.B1(n_65),
.B2(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_10),
.Y(n_80)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_11),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_114),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_113),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_99),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_16),
.B(n_99),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_84),
.B2(n_98),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_46),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_32),
.B1(n_33),
.B2(n_45),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_21),
.A2(n_29),
.B1(n_52),
.B2(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_21),
.B(n_24),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_26),
.A2(n_29),
.B(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_27),
.B(n_164),
.Y(n_163)
);

INVx11_ASAP7_75t_L g139 ( 
.A(n_29),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_29),
.B(n_44),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_32),
.A2(n_33),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_32),
.A2(n_33),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_33),
.B(n_91),
.C(n_154),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_33),
.B(n_131),
.C(n_144),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_34),
.B(n_40),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_40),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_37),
.A2(n_39),
.B(n_44),
.C(n_150),
.Y(n_149)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_40),
.B(n_44),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_44),
.A2(n_63),
.B(n_68),
.C(n_90),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_44),
.A2(n_62),
.B(n_77),
.C(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_58),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_53),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_48),
.A2(n_53),
.B1(n_54),
.B2(n_104),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_48),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_49),
.A2(n_92),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_51),
.B(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_53),
.A2(n_54),
.B1(n_149),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_53),
.A2(n_54),
.B1(n_107),
.B2(n_121),
.Y(n_173)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_54),
.B(n_121),
.C(n_122),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_54),
.B(n_149),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B(n_57),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_73),
.B1(n_74),
.B2(n_83),
.Y(n_58)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_59),
.B(n_107),
.C(n_109),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_59),
.A2(n_83),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_66),
.B(n_69),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_70),
.B1(n_71),
.B2(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_61)
);

INVx5_ASAP7_75t_SL g65 ( 
.A(n_62),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_72)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_81),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_82),
.Y(n_108)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_81),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_94)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_84),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_87),
.C(n_93),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_85),
.A2(n_93),
.B1(n_94),
.B2(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_87),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_88),
.A2(n_89),
.B1(n_91),
.B2(n_155),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_91),
.A2(n_152),
.B1(n_155),
.B2(n_156),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_91),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_91),
.B(n_166),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_93),
.A2(n_94),
.B1(n_133),
.B2(n_140),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_94),
.B(n_134),
.C(n_137),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_97),
.B(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.C(n_105),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_100),
.B(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_103),
.A2(n_105),
.B1(n_106),
.B2(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_103),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_107),
.A2(n_109),
.B1(n_110),
.B2(n_121),
.Y(n_183)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_191),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_186),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_176),
.B(n_185),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_145),
.B(n_175),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_130),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_120),
.B(n_130),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_122),
.B(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_126),
.B1(n_127),
.B2(n_129),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_123),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_129),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_141),
.B2(n_142),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_133),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_136),
.B(n_159),
.Y(n_168)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_137),
.B(n_163),
.Y(n_162)
);

INVx5_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_143),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_170),
.B(n_174),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_157),
.B(n_169),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_151),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_149),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_152),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_153),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_161),
.B(n_168),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_165),
.B(n_167),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_172),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_178),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_182),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_181),
.C(n_182),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_183),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_188),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);


endmodule