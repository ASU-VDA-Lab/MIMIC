module fake_jpeg_13736_n_160 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_160);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_4),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_27),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_8),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_24),
.B(n_7),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_6),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_0),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_73),
.Y(n_83)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_0),
.Y(n_73)
);

BUFx4f_ASAP7_75t_SL g74 ( 
.A(n_56),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_62),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_68),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_64),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_77),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_80)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_50),
.B(n_6),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_75),
.A2(n_65),
.B1(n_66),
.B2(n_49),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_81),
.A2(n_26),
.B1(n_43),
.B2(n_42),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_57),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_87),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_69),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_74),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_57),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_93),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_74),
.B(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_95),
.B(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_91),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_96),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_55),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_98),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_61),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_58),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_99),
.B(n_100),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_1),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_86),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_53),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_103),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_4),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_105),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_50),
.C(n_53),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_109),
.B(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_28),
.C(n_45),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_113),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_13),
.B1(n_16),
.B2(n_18),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_5),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_105),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_115),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_109),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_119),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_122),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_103),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_124),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_107),
.A2(n_23),
.B(n_29),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_30),
.B(n_32),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_41),
.B(n_46),
.Y(n_136)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_34),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_129),
.B(n_123),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_SL g131 ( 
.A(n_109),
.B(n_35),
.C(n_36),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_38),
.C(n_39),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_133),
.B(n_137),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_136),
.A2(n_122),
.B(n_133),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_129),
.Y(n_137)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_126),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_142),
.C(n_145),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_125),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_141),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_117),
.A2(n_130),
.B1(n_132),
.B2(n_124),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_144),
.A2(n_143),
.B1(n_135),
.B2(n_138),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_132),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_151),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_134),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_153),
.B(n_154),
.Y(n_155)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_149),
.Y(n_154)
);

FAx1_ASAP7_75t_SL g156 ( 
.A(n_152),
.B(n_148),
.CI(n_144),
.CON(n_156),
.SN(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_143),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_155),
.C(n_156),
.Y(n_158)
);

BUFx4f_ASAP7_75t_SL g159 ( 
.A(n_158),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_147),
.Y(n_160)
);


endmodule