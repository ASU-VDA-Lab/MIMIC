module fake_netlist_1_5934_n_30 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_30);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NOR2xp33_ASAP7_75t_L g12 ( .A(n_8), .B(n_1), .Y(n_12) );
INVxp33_ASAP7_75t_SL g13 ( .A(n_0), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_9), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_8), .Y(n_15) );
OAI22xp5_ASAP7_75t_L g16 ( .A1(n_6), .A2(n_4), .B1(n_10), .B2(n_2), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_13), .B(n_0), .Y(n_17) );
AOI22xp33_ASAP7_75t_L g18 ( .A1(n_15), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_18) );
O2A1O1Ixp33_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_15), .B(n_16), .C(n_12), .Y(n_19) );
A2O1A1Ixp33_ASAP7_75t_L g20 ( .A1(n_18), .A2(n_16), .B(n_14), .C(n_5), .Y(n_20) );
BUFx6f_ASAP7_75t_L g21 ( .A(n_19), .Y(n_21) );
OR2x2_ASAP7_75t_L g22 ( .A(n_21), .B(n_20), .Y(n_22) );
AND2x4_ASAP7_75t_L g23 ( .A(n_22), .B(n_21), .Y(n_23) );
OAI221xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_21), .B1(n_4), .B2(n_5), .C(n_6), .Y(n_24) );
OAI22xp5_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_23), .B1(n_21), .B2(n_7), .Y(n_25) );
NOR2xp33_ASAP7_75t_L g26 ( .A(n_24), .B(n_23), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
INVx3_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
OAI22xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_25), .B1(n_23), .B2(n_7), .Y(n_29) );
OA22x2_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_28), .B1(n_3), .B2(n_11), .Y(n_30) );
endmodule