module fake_jpeg_8444_n_254 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_254);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_SL g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_39),
.Y(n_50)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_59),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_49),
.A2(n_51),
.B1(n_32),
.B2(n_17),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_22),
.B1(n_24),
.B2(n_29),
.Y(n_51)
);

CKINVDCx6p67_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

INVx5_ASAP7_75t_SL g77 ( 
.A(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_18),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_18),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_20),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_57),
.B(n_58),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_28),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_24),
.B1(n_22),
.B2(n_29),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_63),
.B1(n_68),
.B2(n_19),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_24),
.B1(n_22),
.B2(n_29),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_46),
.A2(n_35),
.B1(n_17),
.B2(n_21),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_31),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_19),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_71),
.A2(n_78),
.B1(n_91),
.B2(n_92),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_40),
.B1(n_39),
.B2(n_38),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_74),
.A2(n_83),
.B1(n_63),
.B2(n_62),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_79),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_65),
.A2(n_39),
.B1(n_28),
.B2(n_37),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_44),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_86),
.Y(n_103)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_85),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_44),
.C(n_28),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_79),
.C(n_87),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_39),
.B1(n_32),
.B2(n_19),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_84),
.Y(n_97)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_66),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_89),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_50),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_67),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_90),
.A2(n_93),
.B1(n_64),
.B2(n_59),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_48),
.A2(n_39),
.B1(n_31),
.B2(n_35),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_48),
.A2(n_31),
.B1(n_23),
.B2(n_27),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_70),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_99),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_98),
.A2(n_114),
.B1(n_90),
.B2(n_81),
.Y(n_136)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_81),
.B1(n_71),
.B2(n_83),
.Y(n_120)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_108),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_93),
.A2(n_62),
.B1(n_54),
.B2(n_53),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_107),
.B1(n_113),
.B2(n_82),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_56),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_116),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_54),
.B1(n_67),
.B2(n_58),
.Y(n_107)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_80),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_109),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_110),
.Y(n_124)
);

AND2x6_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_58),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_111),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_57),
.C(n_50),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_115),
.C(n_84),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_70),
.A2(n_32),
.B1(n_57),
.B2(n_27),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_75),
.B(n_45),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_26),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_117),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_118),
.B1(n_112),
.B2(n_111),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_120),
.A2(n_139),
.B1(n_101),
.B2(n_99),
.Y(n_144)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_122),
.B(n_126),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_140),
.C(n_5),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_114),
.A2(n_108),
.B1(n_96),
.B2(n_102),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_77),
.B(n_73),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_130),
.A2(n_135),
.B(n_116),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_131),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_137),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_77),
.B(n_85),
.Y(n_135)
);

AO21x1_ASAP7_75t_L g145 ( 
.A1(n_136),
.A2(n_107),
.B(n_112),
.Y(n_145)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_18),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_142),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_100),
.A2(n_32),
.B1(n_55),
.B2(n_26),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_45),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_55),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_18),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_143),
.A2(n_149),
.B1(n_153),
.B2(n_154),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_145),
.B1(n_150),
.B2(n_126),
.Y(n_167)
);

XNOR2x1_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_158),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_109),
.B1(n_97),
.B2(n_108),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_128),
.A2(n_113),
.B1(n_21),
.B2(n_23),
.Y(n_150)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_55),
.B1(n_45),
.B2(n_41),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_45),
.B1(n_41),
.B2(n_34),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_41),
.B1(n_34),
.B2(n_33),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_156),
.A2(n_161),
.B1(n_162),
.B2(n_5),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_34),
.B(n_33),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_34),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_165),
.C(n_158),
.Y(n_173)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_160),
.B(n_164),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_120),
.A2(n_33),
.B1(n_16),
.B2(n_4),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_119),
.A2(n_16),
.B1(n_3),
.B2(n_4),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_127),
.A2(n_2),
.B(n_3),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_167),
.A2(n_171),
.B1(n_156),
.B2(n_162),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_147),
.A2(n_137),
.B1(n_122),
.B2(n_139),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_169),
.A2(n_170),
.B(n_145),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_147),
.A2(n_133),
.B1(n_124),
.B2(n_132),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_124),
.B1(n_141),
.B2(n_138),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_178),
.C(n_180),
.Y(n_197)
);

BUFx12_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_142),
.C(n_131),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_5),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_179),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_131),
.C(n_6),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_164),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_182),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_166),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_183),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_184),
.A2(n_149),
.B1(n_161),
.B2(n_165),
.Y(n_198)
);

INVx13_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_186),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_6),
.Y(n_187)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_183),
.A2(n_150),
.B1(n_145),
.B2(n_154),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_176),
.B1(n_185),
.B2(n_186),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_143),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_203),
.C(n_176),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_155),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_191),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_192),
.A2(n_169),
.B1(n_168),
.B2(n_180),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_168),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_163),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_204),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_198),
.B(n_9),
.Y(n_215)
);

NOR3xp33_ASAP7_75t_SL g201 ( 
.A(n_174),
.B(n_148),
.C(n_7),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_SL g210 ( 
.A(n_201),
.B(n_7),
.C(n_9),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_173),
.C(n_177),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_167),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_6),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_10),
.Y(n_217)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_211),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_196),
.A2(n_172),
.B(n_170),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_212),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_209),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_215),
.Y(n_225)
);

OA21x2_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_175),
.B(n_10),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_197),
.C(n_190),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_197),
.C(n_194),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_175),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_205),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_195),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_224),
.Y(n_234)
);

FAx1_ASAP7_75t_SL g222 ( 
.A(n_218),
.B(n_191),
.CI(n_189),
.CON(n_222),
.SN(n_222)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_213),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_226),
.Y(n_233)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_201),
.C(n_192),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_227),
.A2(n_188),
.B1(n_199),
.B2(n_212),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_223),
.A2(n_206),
.B(n_202),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_219),
.C(n_11),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_220),
.A2(n_207),
.B1(n_214),
.B2(n_216),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_230),
.A2(n_227),
.B1(n_224),
.B2(n_228),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_231),
.A2(n_236),
.B1(n_221),
.B2(n_233),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_193),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_235),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_212),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_241),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_239),
.A2(n_240),
.B1(n_234),
.B2(n_11),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_230),
.A2(n_199),
.B1(n_219),
.B2(n_193),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_200),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_10),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_243),
.A2(n_246),
.B(n_240),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_242),
.A2(n_234),
.B(n_12),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_244),
.A2(n_237),
.B(n_238),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_13),
.Y(n_250)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_248),
.A2(n_249),
.B(n_14),
.Y(n_251)
);

OAI21x1_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_15),
.B(n_13),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_250),
.B(n_251),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_14),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_15),
.Y(n_254)
);


endmodule