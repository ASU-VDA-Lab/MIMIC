module fake_jpeg_20310_n_164 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_0),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_0),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_41),
.Y(n_50)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_1),
.Y(n_41)
);

AO22x2_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_30),
.B1(n_28),
.B2(n_16),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_39),
.B1(n_31),
.B2(n_36),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_55),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_33),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_23),
.B1(n_29),
.B2(n_30),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_57),
.Y(n_60)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_62),
.B(n_64),
.Y(n_87)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_17),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_54),
.Y(n_66)
);

INVx5_ASAP7_75t_SL g93 ( 
.A(n_66),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_67),
.B(n_69),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_73),
.B1(n_84),
.B2(n_1),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_18),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_74),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_36),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_77),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_40),
.B(n_29),
.C(n_26),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_24),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_40),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_79),
.C(n_81),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_35),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_24),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_35),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_20),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_28),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_82),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_20),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_3),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_45),
.A2(n_15),
.B1(n_27),
.B2(n_25),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_15),
.B1(n_28),
.B2(n_25),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_68),
.Y(n_108)
);

MAJx2_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_58),
.C(n_59),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_100),
.C(n_66),
.Y(n_120)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_99),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_3),
.C(n_4),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_101),
.B(n_105),
.Y(n_113)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_84),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_76),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_82),
.Y(n_105)
);

OR2x2_ASAP7_75t_SL g107 ( 
.A(n_89),
.B(n_60),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_119),
.B(n_120),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_121),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_72),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_111),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_75),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_90),
.B(n_79),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_116),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_73),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_77),
.B(n_76),
.C(n_66),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_118),
.Y(n_130)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_65),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_107),
.A2(n_86),
.B(n_105),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_122),
.A2(n_93),
.B(n_103),
.C(n_106),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_92),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_127),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_86),
.B(n_88),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_92),
.C(n_96),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_93),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_87),
.B(n_91),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_132),
.A2(n_110),
.B(n_99),
.Y(n_135)
);

AOI322xp5_ASAP7_75t_SL g133 ( 
.A1(n_123),
.A2(n_113),
.A3(n_100),
.B1(n_7),
.B2(n_8),
.C1(n_11),
.C2(n_5),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_133),
.B(n_5),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_130),
.A2(n_121),
.B(n_115),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_134),
.A2(n_135),
.B(n_139),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_125),
.A2(n_112),
.B1(n_96),
.B2(n_106),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_138),
.Y(n_146)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_140),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_124),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_122),
.B(n_126),
.Y(n_144)
);

OAI21x1_ASAP7_75t_L g155 ( 
.A1(n_144),
.A2(n_65),
.B(n_97),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_148),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_134),
.A2(n_132),
.B(n_129),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_147),
.A2(n_139),
.B(n_137),
.Y(n_151)
);

AO21x1_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_139),
.B(n_140),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_152),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_153),
.B1(n_6),
.B2(n_8),
.Y(n_159)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_149),
.A2(n_146),
.B(n_139),
.Y(n_153)
);

NOR2x1_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_143),
.Y(n_156)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_156),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_97),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_158),
.A2(n_159),
.B(n_13),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_11),
.C(n_12),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_157),
.B(n_158),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_163),
.Y(n_164)
);


endmodule