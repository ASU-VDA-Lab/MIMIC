module fake_jpeg_4639_n_21 (n_0, n_3, n_2, n_1, n_21);

input n_0;
input n_3;
input n_2;
input n_1;

output n_21;

wire n_13;
wire n_10;
wire n_6;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_4;
wire n_16;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx8_ASAP7_75t_L g4 ( 
.A(n_2),
.Y(n_4)
);

BUFx3_ASAP7_75t_L g5 ( 
.A(n_3),
.Y(n_5)
);

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

INVx8_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_L g9 ( 
.A1(n_4),
.A2(n_3),
.B1(n_0),
.B2(n_1),
.Y(n_9)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_9),
.B(n_10),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_L g10 ( 
.A1(n_5),
.A2(n_0),
.B(n_1),
.Y(n_10)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_12),
.A2(n_10),
.B1(n_8),
.B2(n_4),
.Y(n_13)
);

XNOR2xp5_ASAP7_75t_SL g16 ( 
.A(n_13),
.B(n_6),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_12),
.B(n_0),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_14),
.B(n_1),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_16),
.C(n_13),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_17),
.A2(n_18),
.B(n_5),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_16),
.B(n_11),
.C(n_4),
.Y(n_18)
);

AO21x1_ASAP7_75t_L g20 ( 
.A1(n_19),
.A2(n_3),
.B(n_6),
.Y(n_20)
);

NAND3xp33_ASAP7_75t_SL g21 ( 
.A(n_20),
.B(n_7),
.C(n_0),
.Y(n_21)
);


endmodule