module fake_ariane_2432_n_1109 (n_295, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_294, n_197, n_176, n_34, n_172, n_183, n_299, n_12, n_133, n_66, n_205, n_71, n_109, n_245, n_96, n_49, n_20, n_283, n_50, n_187, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_214, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_77, n_15, n_23, n_87, n_279, n_207, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_239, n_35, n_272, n_54, n_8, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_115, n_267, n_291, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_227, n_48, n_188, n_11, n_129, n_126, n_282, n_277, n_248, n_301, n_293, n_228, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_238, n_136, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_16, n_273, n_305, n_233, n_56, n_60, n_221, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_26, n_246, n_0, n_159, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_101, n_243, n_134, n_185, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_22, n_241, n_29, n_191, n_80, n_211, n_97, n_251, n_116, n_39, n_155, n_127, n_1109);

input n_295;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_71;
input n_109;
input n_245;
input n_96;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_214;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_115;
input n_267;
input n_291;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_227;
input n_48;
input n_188;
input n_11;
input n_129;
input n_126;
input n_282;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_238;
input n_136;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_16;
input n_273;
input n_305;
input n_233;
input n_56;
input n_60;
input n_221;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_26;
input n_246;
input n_0;
input n_159;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_101;
input n_243;
input n_134;
input n_185;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_22;
input n_241;
input n_29;
input n_191;
input n_80;
input n_211;
input n_97;
input n_251;
input n_116;
input n_39;
input n_155;
input n_127;

output n_1109;

wire n_356;
wire n_556;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_908;
wire n_850;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_643;
wire n_679;
wire n_924;
wire n_927;
wire n_781;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_586;
wire n_443;
wire n_864;
wire n_952;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_528;
wire n_584;
wire n_424;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_349;
wire n_634;
wire n_391;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_1016;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_891;
wire n_737;
wire n_885;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_790;
wire n_898;
wire n_857;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_1064;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_1093;
wire n_473;
wire n_801;
wire n_733;
wire n_818;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_311;
wire n_402;
wire n_1052;
wire n_1068;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_835;
wire n_808;
wire n_953;
wire n_553;
wire n_446;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_1107;
wire n_858;
wire n_645;
wire n_989;
wire n_331;
wire n_320;
wire n_559;
wire n_485;
wire n_401;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_1090;
wire n_529;
wire n_502;
wire n_561;
wire n_821;
wire n_770;
wire n_839;
wire n_928;
wire n_1099;
wire n_465;
wire n_507;
wire n_486;
wire n_901;
wire n_759;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_971;
wire n_369;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_604;
wire n_439;
wire n_614;
wire n_677;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_997;
wire n_635;
wire n_707;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_983;
wire n_328;
wire n_368;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_644;
wire n_536;
wire n_823;
wire n_921;
wire n_620;
wire n_325;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_365;
wire n_429;
wire n_654;
wire n_455;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_539;
wire n_312;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_911;
wire n_458;
wire n_361;
wire n_383;
wire n_623;
wire n_838;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_705;
wire n_630;
wire n_658;
wire n_570;
wire n_1055;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_628;
wire n_809;
wire n_461;
wire n_490;
wire n_743;
wire n_907;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_534;
wire n_1108;
wire n_355;
wire n_609;
wire n_444;
wire n_851;
wire n_1043;
wire n_560;
wire n_450;
wire n_890;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_982;
wire n_915;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_862;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1100;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_697;
wire n_622;
wire n_967;
wire n_999;
wire n_998;
wire n_1083;
wire n_472;
wire n_937;
wire n_746;
wire n_456;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_704;
wire n_1060;
wire n_1044;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_580;
wire n_358;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_563;
wire n_394;
wire n_923;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_972;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_484;
wire n_411;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_54),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_287),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_116),
.Y(n_312)
);

INVxp33_ASAP7_75t_SL g313 ( 
.A(n_13),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_130),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_87),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_194),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_L g317 ( 
.A(n_167),
.B(n_235),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_284),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_51),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_106),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_296),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_23),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_L g323 ( 
.A(n_42),
.B(n_218),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_52),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_107),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_253),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_169),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_222),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_168),
.Y(n_329)
);

BUFx2_ASAP7_75t_SL g330 ( 
.A(n_189),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_226),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_248),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_204),
.Y(n_333)
);

BUFx5_ASAP7_75t_L g334 ( 
.A(n_209),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_173),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_212),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_202),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_164),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_238),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_196),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_20),
.B(n_102),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_108),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_86),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_243),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_271),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_90),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_4),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_260),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_71),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_104),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_309),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_220),
.Y(n_352)
);

INVxp33_ASAP7_75t_SL g353 ( 
.A(n_51),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_264),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_225),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_170),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_294),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_178),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_251),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_282),
.Y(n_360)
);

BUFx2_ASAP7_75t_SL g361 ( 
.A(n_115),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_231),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_125),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_24),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_233),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_67),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_109),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_180),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_191),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_106),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_278),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_262),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_279),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_265),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_207),
.B(n_308),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_129),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_123),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_299),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_261),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_72),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_234),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_126),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_49),
.Y(n_383)
);

BUFx10_ASAP7_75t_L g384 ( 
.A(n_70),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_14),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_165),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_183),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_273),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_132),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_182),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_276),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_297),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_105),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_188),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_137),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_141),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_54),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_181),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_163),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_229),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_L g401 ( 
.A(n_140),
.B(n_301),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_263),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_108),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_195),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_87),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_139),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_44),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_275),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_203),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_138),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_224),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_26),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_124),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_127),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_232),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_160),
.Y(n_416)
);

BUFx8_ASAP7_75t_SL g417 ( 
.A(n_110),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_286),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_185),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_280),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_48),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_7),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_119),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_187),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_34),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_154),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_208),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_64),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_144),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_166),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_205),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_99),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_32),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_157),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_258),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_268),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_153),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_88),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_285),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_122),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_95),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_84),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_131),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_128),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_85),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_283),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_175),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_133),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_45),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_103),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_94),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_155),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_72),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_17),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_147),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_242),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_136),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_199),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_198),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_107),
.Y(n_460)
);

NOR2xp67_ASAP7_75t_L g461 ( 
.A(n_239),
.B(n_277),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_206),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_241),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_3),
.Y(n_464)
);

BUFx5_ASAP7_75t_L g465 ( 
.A(n_36),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_310),
.A2(n_325),
.B1(n_432),
.B2(n_366),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_322),
.B(n_0),
.Y(n_467)
);

OAI21x1_ASAP7_75t_L g468 ( 
.A1(n_406),
.A2(n_434),
.B(n_365),
.Y(n_468)
);

OAI21x1_ASAP7_75t_L g469 ( 
.A1(n_406),
.A2(n_434),
.B(n_365),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_421),
.B(n_1),
.Y(n_470)
);

AND2x6_ASAP7_75t_L g471 ( 
.A(n_314),
.B(n_379),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_421),
.B(n_1),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_364),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_386),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_465),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_2),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_386),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_433),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_318),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_433),
.Y(n_480)
);

OAI22x1_ASAP7_75t_R g481 ( 
.A1(n_405),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_481)
);

NOR2x1_ASAP7_75t_L g482 ( 
.A(n_390),
.B(n_118),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_453),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_465),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_390),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_369),
.B(n_5),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_413),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_311),
.B(n_8),
.Y(n_488)
);

OA21x2_ASAP7_75t_L g489 ( 
.A1(n_316),
.A2(n_8),
.B(n_9),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_413),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_384),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_415),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_364),
.Y(n_493)
);

CKINVDCx6p67_ASAP7_75t_R g494 ( 
.A(n_368),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_458),
.B(n_9),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_384),
.B(n_10),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_328),
.B(n_10),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_312),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_326),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_499)
);

BUFx8_ASAP7_75t_SL g500 ( 
.A(n_417),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_329),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_458),
.Y(n_502)
);

OAI21x1_ASAP7_75t_L g503 ( 
.A1(n_314),
.A2(n_121),
.B(n_120),
.Y(n_503)
);

BUFx12f_ASAP7_75t_L g504 ( 
.A(n_324),
.Y(n_504)
);

OA21x2_ASAP7_75t_L g505 ( 
.A1(n_331),
.A2(n_11),
.B(n_12),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_315),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_393),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_319),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_320),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_350),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_403),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_346),
.B(n_14),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_333),
.B(n_15),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_403),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_403),
.Y(n_515)
);

OA21x2_ASAP7_75t_L g516 ( 
.A1(n_335),
.A2(n_15),
.B(n_16),
.Y(n_516)
);

OA21x2_ASAP7_75t_L g517 ( 
.A1(n_337),
.A2(n_16),
.B(n_17),
.Y(n_517)
);

BUFx12f_ASAP7_75t_L g518 ( 
.A(n_342),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_338),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_519)
);

INVx5_ASAP7_75t_L g520 ( 
.A(n_452),
.Y(n_520)
);

OA21x2_ASAP7_75t_L g521 ( 
.A1(n_340),
.A2(n_18),
.B(n_19),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_367),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_380),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_344),
.B(n_21),
.Y(n_524)
);

INVx5_ASAP7_75t_L g525 ( 
.A(n_382),
.Y(n_525)
);

OA21x2_ASAP7_75t_L g526 ( 
.A1(n_348),
.A2(n_21),
.B(n_22),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_383),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_385),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_382),
.Y(n_529)
);

OA21x2_ASAP7_75t_L g530 ( 
.A1(n_351),
.A2(n_22),
.B(n_23),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_397),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_414),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_422),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_352),
.B(n_24),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_428),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_438),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_414),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_345),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_354),
.Y(n_539)
);

BUFx10_ASAP7_75t_L g540 ( 
.A(n_501),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_507),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_494),
.A2(n_339),
.B1(n_436),
.B2(n_402),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_466),
.B(n_437),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_538),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_484),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_474),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_507),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_507),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_479),
.B(n_356),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_507),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_485),
.B(n_357),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_495),
.B(n_448),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_SL g553 ( 
.A(n_538),
.B(n_447),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_520),
.B(n_388),
.Y(n_554)
);

BUFx10_ASAP7_75t_L g555 ( 
.A(n_495),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_474),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_480),
.B(n_441),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_485),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_525),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_511),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_498),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_506),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_491),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_520),
.B(n_360),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_L g565 ( 
.A(n_471),
.B(n_334),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_511),
.Y(n_566)
);

NOR2x1p5_ASAP7_75t_L g567 ( 
.A(n_504),
.B(n_343),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_508),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_509),
.Y(n_569)
);

INVx8_ASAP7_75t_L g570 ( 
.A(n_520),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_474),
.Y(n_571)
);

AND3x2_ASAP7_75t_L g572 ( 
.A(n_496),
.B(n_388),
.C(n_341),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_520),
.B(n_362),
.Y(n_573)
);

NAND3xp33_ASAP7_75t_L g574 ( 
.A(n_486),
.B(n_370),
.C(n_347),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_473),
.B(n_442),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_511),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_514),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_510),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_531),
.Y(n_579)
);

BUFx6f_ASAP7_75t_SL g580 ( 
.A(n_467),
.Y(n_580)
);

OAI22xp33_ASAP7_75t_L g581 ( 
.A1(n_499),
.A2(n_349),
.B1(n_407),
.B2(n_353),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_518),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_477),
.Y(n_583)
);

NAND3xp33_ASAP7_75t_L g584 ( 
.A(n_486),
.B(n_425),
.C(n_412),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_514),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_467),
.B(n_448),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_533),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_466),
.B(n_313),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_478),
.B(n_371),
.Y(n_589)
);

OAI22xp33_ASAP7_75t_L g590 ( 
.A1(n_581),
.A2(n_519),
.B1(n_483),
.B2(n_523),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_552),
.B(n_525),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_545),
.B(n_525),
.Y(n_592)
);

A2O1A1Ixp33_ASAP7_75t_L g593 ( 
.A1(n_586),
.A2(n_513),
.B(n_534),
.C(n_476),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_586),
.B(n_539),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_553),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_558),
.B(n_539),
.Y(n_596)
);

NOR3xp33_ASAP7_75t_L g597 ( 
.A(n_581),
.B(n_483),
.C(n_488),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_554),
.B(n_477),
.Y(n_598)
);

A2O1A1Ixp33_ASAP7_75t_L g599 ( 
.A1(n_554),
.A2(n_513),
.B(n_534),
.C(n_476),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_546),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_546),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_582),
.B(n_481),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_561),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_549),
.B(n_555),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_544),
.B(n_470),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_562),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_568),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_556),
.B(n_477),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_556),
.B(n_477),
.Y(n_609)
);

NOR2xp67_ASAP7_75t_L g610 ( 
.A(n_544),
.B(n_473),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_571),
.B(n_487),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_565),
.A2(n_512),
.B1(n_471),
.B2(n_505),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_571),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_569),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_583),
.B(n_487),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_578),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_579),
.Y(n_617)
);

NOR2xp67_ASAP7_75t_L g618 ( 
.A(n_563),
.B(n_493),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_587),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_583),
.B(n_487),
.Y(n_620)
);

OAI22xp33_ASAP7_75t_L g621 ( 
.A1(n_542),
.A2(n_497),
.B1(n_524),
.B2(n_575),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_541),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_551),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_580),
.A2(n_472),
.B1(n_512),
.B2(n_460),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_557),
.Y(n_625)
);

OAI22xp33_ASAP7_75t_L g626 ( 
.A1(n_574),
.A2(n_493),
.B1(n_449),
.B2(n_450),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_589),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_572),
.B(n_472),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_570),
.B(n_487),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_580),
.B(n_584),
.Y(n_630)
);

OR2x2_ASAP7_75t_SL g631 ( 
.A(n_588),
.B(n_500),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_540),
.B(n_464),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_540),
.B(n_490),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_565),
.A2(n_471),
.B1(n_505),
.B2(n_489),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_547),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_572),
.B(n_490),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_564),
.B(n_573),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_547),
.Y(n_638)
);

AO22x1_ASAP7_75t_L g639 ( 
.A1(n_548),
.A2(n_471),
.B1(n_451),
.B2(n_454),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_567),
.B(n_522),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_559),
.B(n_492),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_559),
.B(n_527),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_585),
.B(n_528),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_550),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_576),
.B(n_502),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_560),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_566),
.B(n_502),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_637),
.A2(n_469),
.B(n_468),
.Y(n_648)
);

NAND3xp33_ASAP7_75t_L g649 ( 
.A(n_597),
.B(n_435),
.C(n_445),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_610),
.B(n_535),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_623),
.B(n_604),
.Y(n_651)
);

A2O1A1Ixp33_ASAP7_75t_L g652 ( 
.A1(n_599),
.A2(n_323),
.B(n_503),
.C(n_475),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_618),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_627),
.A2(n_482),
.B(n_489),
.Y(n_654)
);

BUFx8_ASAP7_75t_L g655 ( 
.A(n_628),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_598),
.A2(n_517),
.B(n_516),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_644),
.Y(n_657)
);

AOI22x1_ASAP7_75t_L g658 ( 
.A1(n_603),
.A2(n_361),
.B1(n_330),
.B2(n_577),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_593),
.A2(n_517),
.B1(n_521),
.B2(n_516),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_606),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_607),
.B(n_614),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_616),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_600),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_617),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_641),
.A2(n_530),
.B(n_526),
.Y(n_665)
);

BUFx4f_ASAP7_75t_L g666 ( 
.A(n_640),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_619),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_625),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_L g669 ( 
.A1(n_634),
.A2(n_375),
.B(n_530),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_628),
.B(n_321),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_608),
.Y(n_671)
);

AOI221xp5_ASAP7_75t_L g672 ( 
.A1(n_590),
.A2(n_536),
.B1(n_389),
.B2(n_391),
.C(n_381),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_633),
.A2(n_375),
.B(n_372),
.Y(n_673)
);

AO22x1_ASAP7_75t_L g674 ( 
.A1(n_597),
.A2(n_327),
.B1(n_378),
.B2(n_376),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_595),
.B(n_515),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_609),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_594),
.B(n_399),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_L g678 ( 
.A1(n_624),
.A2(n_605),
.B1(n_612),
.B2(n_632),
.Y(n_678)
);

OAI21xp33_ASAP7_75t_L g679 ( 
.A1(n_630),
.A2(n_626),
.B(n_590),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_642),
.Y(n_680)
);

BUFx12f_ASAP7_75t_L g681 ( 
.A(n_631),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_596),
.B(n_416),
.Y(n_682)
);

A2O1A1Ixp33_ASAP7_75t_L g683 ( 
.A1(n_612),
.A2(n_636),
.B(n_601),
.C(n_613),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_611),
.Y(n_684)
);

AOI22x1_ASAP7_75t_L g685 ( 
.A1(n_622),
.A2(n_396),
.B1(n_398),
.B2(n_395),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_595),
.B(n_400),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_592),
.A2(n_423),
.B(n_411),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_615),
.Y(n_688)
);

O2A1O1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_626),
.A2(n_621),
.B(n_620),
.C(n_645),
.Y(n_689)
);

CKINVDCx10_ASAP7_75t_R g690 ( 
.A(n_602),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_591),
.A2(n_429),
.B1(n_430),
.B2(n_427),
.Y(n_691)
);

NOR2x1p5_ASAP7_75t_SL g692 ( 
.A(n_638),
.B(n_334),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_629),
.A2(n_439),
.B(n_431),
.Y(n_693)
);

BUFx8_ASAP7_75t_SL g694 ( 
.A(n_602),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_602),
.B(n_529),
.Y(n_695)
);

AO21x2_ASAP7_75t_L g696 ( 
.A1(n_646),
.A2(n_401),
.B(n_317),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_647),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_635),
.Y(n_698)
);

O2A1O1Ixp5_ASAP7_75t_L g699 ( 
.A1(n_639),
.A2(n_459),
.B(n_457),
.C(n_463),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_L g700 ( 
.A(n_597),
.B(n_532),
.C(n_529),
.Y(n_700)
);

OAI21xp5_ASAP7_75t_L g701 ( 
.A1(n_599),
.A2(n_461),
.B(n_332),
.Y(n_701)
);

A2O1A1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_599),
.A2(n_537),
.B(n_532),
.C(n_336),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_628),
.B(n_532),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_610),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_643),
.Y(n_705)
);

INVxp67_ASAP7_75t_SL g706 ( 
.A(n_610),
.Y(n_706)
);

O2A1O1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_599),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_707)
);

A2O1A1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_599),
.A2(n_537),
.B(n_358),
.C(n_359),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_643),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_610),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_623),
.B(n_355),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_643),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_610),
.B(n_363),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_643),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_623),
.B(n_373),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_637),
.A2(n_377),
.B(n_374),
.Y(n_716)
);

INVx5_ASAP7_75t_L g717 ( 
.A(n_628),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_623),
.B(n_387),
.Y(n_718)
);

AO22x1_ASAP7_75t_L g719 ( 
.A1(n_597),
.A2(n_394),
.B1(n_404),
.B2(n_392),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_637),
.A2(n_409),
.B(n_408),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_623),
.B(n_410),
.Y(n_721)
);

BUFx2_ASAP7_75t_L g722 ( 
.A(n_628),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_643),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_644),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_644),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_610),
.B(n_418),
.Y(n_726)
);

AO32x1_ASAP7_75t_L g727 ( 
.A1(n_638),
.A2(n_334),
.A3(n_576),
.B1(n_514),
.B2(n_28),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_637),
.A2(n_420),
.B(n_419),
.Y(n_728)
);

AOI21x1_ASAP7_75t_L g729 ( 
.A1(n_665),
.A2(n_656),
.B(n_648),
.Y(n_729)
);

NOR2xp67_ASAP7_75t_SL g730 ( 
.A(n_717),
.B(n_424),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_660),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_651),
.B(n_426),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_711),
.B(n_718),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_650),
.B(n_440),
.Y(n_734)
);

OAI21x1_ASAP7_75t_L g735 ( 
.A1(n_669),
.A2(n_654),
.B(n_659),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_662),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_678),
.B(n_443),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_722),
.Y(n_738)
);

AOI21xp33_ASAP7_75t_L g739 ( 
.A1(n_686),
.A2(n_446),
.B(n_444),
.Y(n_739)
);

OR2x6_ASAP7_75t_L g740 ( 
.A(n_681),
.B(n_514),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_668),
.B(n_25),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_712),
.B(n_455),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_666),
.B(n_695),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_655),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_657),
.Y(n_745)
);

AO31x2_ASAP7_75t_L g746 ( 
.A1(n_652),
.A2(n_30),
.A3(n_28),
.B(n_29),
.Y(n_746)
);

OAI21xp5_ASAP7_75t_L g747 ( 
.A1(n_702),
.A2(n_462),
.B(n_456),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_675),
.B(n_29),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_661),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_664),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_667),
.A2(n_34),
.B1(n_31),
.B2(n_33),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_694),
.Y(n_752)
);

NAND3xp33_ASAP7_75t_SL g753 ( 
.A(n_672),
.B(n_649),
.C(n_701),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_724),
.Y(n_754)
);

AOI221xp5_ASAP7_75t_SL g755 ( 
.A1(n_708),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.C(n_38),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_724),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_715),
.B(n_37),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_725),
.Y(n_758)
);

NAND2x1p5_ASAP7_75t_L g759 ( 
.A(n_680),
.B(n_38),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_721),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_706),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_705),
.B(n_43),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_725),
.Y(n_763)
);

OAI21x1_ASAP7_75t_L g764 ( 
.A1(n_673),
.A2(n_135),
.B(n_134),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_725),
.B(n_46),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_709),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_714),
.B(n_46),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_723),
.B(n_47),
.Y(n_768)
);

AO31x2_ASAP7_75t_L g769 ( 
.A1(n_683),
.A2(n_49),
.A3(n_47),
.B(n_48),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_682),
.B(n_50),
.Y(n_770)
);

OAI21xp5_ASAP7_75t_SL g771 ( 
.A1(n_707),
.A2(n_50),
.B(n_52),
.Y(n_771)
);

OAI22x1_ASAP7_75t_L g772 ( 
.A1(n_670),
.A2(n_56),
.B1(n_53),
.B2(n_55),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_697),
.Y(n_773)
);

OAI21xp5_ASAP7_75t_L g774 ( 
.A1(n_671),
.A2(n_143),
.B(n_142),
.Y(n_774)
);

AO22x2_ASAP7_75t_L g775 ( 
.A1(n_674),
.A2(n_56),
.B1(n_53),
.B2(n_55),
.Y(n_775)
);

OAI21x1_ASAP7_75t_L g776 ( 
.A1(n_693),
.A2(n_146),
.B(n_145),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_676),
.A2(n_688),
.B(n_684),
.Y(n_777)
);

BUFx2_ASAP7_75t_L g778 ( 
.A(n_710),
.Y(n_778)
);

OA21x2_ASAP7_75t_L g779 ( 
.A1(n_700),
.A2(n_149),
.B(n_148),
.Y(n_779)
);

OAI222xp33_ASAP7_75t_L g780 ( 
.A1(n_691),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.C1(n_60),
.C2(n_61),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_704),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_677),
.B(n_60),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_719),
.B(n_61),
.Y(n_783)
);

INVxp67_ASAP7_75t_SL g784 ( 
.A(n_689),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_663),
.B(n_62),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_728),
.A2(n_151),
.B(n_150),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_653),
.B(n_63),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_698),
.Y(n_788)
);

INVxp67_ASAP7_75t_SL g789 ( 
.A(n_697),
.Y(n_789)
);

A2O1A1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_687),
.A2(n_66),
.B(n_64),
.C(n_65),
.Y(n_790)
);

OAI21x1_ASAP7_75t_L g791 ( 
.A1(n_699),
.A2(n_156),
.B(n_152),
.Y(n_791)
);

INVx1_ASAP7_75t_SL g792 ( 
.A(n_690),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_696),
.Y(n_793)
);

OAI21xp33_ASAP7_75t_L g794 ( 
.A1(n_713),
.A2(n_67),
.B(n_68),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_726),
.Y(n_795)
);

AO31x2_ASAP7_75t_L g796 ( 
.A1(n_727),
.A2(n_71),
.A3(n_69),
.B(n_70),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_L g797 ( 
.A1(n_716),
.A2(n_74),
.B1(n_69),
.B2(n_73),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_720),
.A2(n_159),
.B(n_158),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_727),
.A2(n_658),
.B(n_685),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_692),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_660),
.Y(n_801)
);

AO31x2_ASAP7_75t_L g802 ( 
.A1(n_659),
.A2(n_78),
.A3(n_76),
.B(n_77),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_660),
.Y(n_803)
);

NAND2x1p5_ASAP7_75t_L g804 ( 
.A(n_717),
.B(n_77),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_679),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_651),
.B(n_79),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_648),
.A2(n_162),
.B(n_161),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_660),
.Y(n_808)
);

OAI22x1_ASAP7_75t_L g809 ( 
.A1(n_649),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_809)
);

AO22x2_ASAP7_75t_L g810 ( 
.A1(n_678),
.A2(n_84),
.B1(n_86),
.B2(n_88),
.Y(n_810)
);

NAND2x1p5_ASAP7_75t_L g811 ( 
.A(n_717),
.B(n_89),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_648),
.A2(n_172),
.B(n_171),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_648),
.A2(n_176),
.B(n_174),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_648),
.A2(n_179),
.B(n_177),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_651),
.B(n_90),
.Y(n_815)
);

NAND2x1p5_ASAP7_75t_L g816 ( 
.A(n_717),
.B(n_91),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_651),
.B(n_92),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_722),
.B(n_92),
.Y(n_818)
);

AO32x2_ASAP7_75t_L g819 ( 
.A1(n_659),
.A2(n_93),
.A3(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_651),
.B(n_96),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_660),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_651),
.B(n_97),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_694),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_651),
.B(n_98),
.Y(n_824)
);

AO31x2_ASAP7_75t_L g825 ( 
.A1(n_659),
.A2(n_99),
.A3(n_100),
.B(n_101),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_679),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_651),
.B(n_103),
.Y(n_827)
);

AND2x6_ASAP7_75t_L g828 ( 
.A(n_703),
.B(n_184),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_648),
.A2(n_190),
.B(n_186),
.Y(n_829)
);

OAI21xp5_ASAP7_75t_L g830 ( 
.A1(n_648),
.A2(n_193),
.B(n_192),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_743),
.B(n_110),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_784),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_733),
.B(n_111),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_763),
.Y(n_834)
);

CKINVDCx11_ASAP7_75t_R g835 ( 
.A(n_752),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_731),
.Y(n_836)
);

INVx8_ASAP7_75t_L g837 ( 
.A(n_823),
.Y(n_837)
);

AO221x2_ASAP7_75t_L g838 ( 
.A1(n_780),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.C(n_114),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_753),
.A2(n_112),
.B(n_114),
.C(n_116),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_736),
.Y(n_840)
);

INVx8_ASAP7_75t_L g841 ( 
.A(n_740),
.Y(n_841)
);

NAND2x1p5_ASAP7_75t_L g842 ( 
.A(n_745),
.B(n_197),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_750),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_801),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_732),
.B(n_117),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_803),
.Y(n_846)
);

AO21x2_ASAP7_75t_L g847 ( 
.A1(n_729),
.A2(n_200),
.B(n_201),
.Y(n_847)
);

AO22x1_ASAP7_75t_L g848 ( 
.A1(n_744),
.A2(n_210),
.B1(n_211),
.B2(n_213),
.Y(n_848)
);

OAI22xp33_ASAP7_75t_L g849 ( 
.A1(n_815),
.A2(n_307),
.B1(n_214),
.B2(n_215),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_810),
.A2(n_216),
.B1(n_217),
.B2(n_219),
.Y(n_850)
);

INVxp67_ASAP7_75t_L g851 ( 
.A(n_738),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_810),
.A2(n_793),
.B1(n_766),
.B2(n_788),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_808),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_817),
.A2(n_221),
.B(n_223),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_756),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_822),
.A2(n_227),
.B1(n_228),
.B2(n_230),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_741),
.B(n_306),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_821),
.Y(n_858)
);

A2O1A1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_737),
.A2(n_236),
.B(n_237),
.C(n_240),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_818),
.B(n_305),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_758),
.Y(n_861)
);

INVx6_ASAP7_75t_L g862 ( 
.A(n_740),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_754),
.B(n_778),
.Y(n_863)
);

INVx3_ASAP7_75t_SL g864 ( 
.A(n_792),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_769),
.Y(n_865)
);

OA21x2_ASAP7_75t_L g866 ( 
.A1(n_830),
.A2(n_244),
.B(n_245),
.Y(n_866)
);

AO21x2_ASAP7_75t_L g867 ( 
.A1(n_774),
.A2(n_246),
.B(n_247),
.Y(n_867)
);

OAI221xp5_ASAP7_75t_SL g868 ( 
.A1(n_805),
.A2(n_249),
.B1(n_250),
.B2(n_252),
.C(n_254),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_795),
.B(n_255),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_757),
.A2(n_256),
.B1(n_257),
.B2(n_259),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_746),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_782),
.A2(n_770),
.B1(n_820),
.B2(n_827),
.Y(n_872)
);

BUFx2_ASAP7_75t_L g873 ( 
.A(n_765),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_746),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_748),
.B(n_734),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_824),
.A2(n_266),
.B1(n_267),
.B2(n_269),
.Y(n_876)
);

OR2x6_ASAP7_75t_L g877 ( 
.A(n_804),
.B(n_270),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_762),
.B(n_272),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_746),
.Y(n_879)
);

OAI21x1_ASAP7_75t_L g880 ( 
.A1(n_812),
.A2(n_829),
.B(n_813),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_739),
.B(n_274),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_828),
.Y(n_882)
);

OAI21x1_ASAP7_75t_L g883 ( 
.A1(n_814),
.A2(n_281),
.B(n_288),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_775),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_884)
);

OAI21x1_ASAP7_75t_SL g885 ( 
.A1(n_783),
.A2(n_292),
.B(n_293),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_787),
.B(n_304),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_767),
.B(n_295),
.Y(n_887)
);

OAI21xp5_ASAP7_75t_L g888 ( 
.A1(n_768),
.A2(n_298),
.B(n_300),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_811),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_816),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_773),
.Y(n_891)
);

AOI211xp5_ASAP7_75t_L g892 ( 
.A1(n_761),
.A2(n_302),
.B(n_303),
.C(n_781),
.Y(n_892)
);

CKINVDCx20_ASAP7_75t_R g893 ( 
.A(n_742),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_785),
.Y(n_894)
);

AO21x2_ASAP7_75t_L g895 ( 
.A1(n_747),
.A2(n_798),
.B(n_786),
.Y(n_895)
);

OR2x6_ASAP7_75t_L g896 ( 
.A(n_759),
.B(n_775),
.Y(n_896)
);

NAND2x1p5_ASAP7_75t_L g897 ( 
.A(n_730),
.B(n_779),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_809),
.Y(n_898)
);

OAI222xp33_ASAP7_75t_L g899 ( 
.A1(n_826),
.A2(n_751),
.B1(n_749),
.B2(n_760),
.C1(n_797),
.C2(n_800),
.Y(n_899)
);

OA21x2_ASAP7_75t_L g900 ( 
.A1(n_764),
.A2(n_791),
.B(n_776),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_789),
.B(n_771),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_794),
.A2(n_755),
.B(n_802),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_790),
.B(n_802),
.Y(n_903)
);

CKINVDCx16_ASAP7_75t_R g904 ( 
.A(n_772),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_819),
.B(n_825),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_819),
.A2(n_588),
.B1(n_679),
.B2(n_543),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_796),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_796),
.A2(n_588),
.B1(n_679),
.B2(n_543),
.Y(n_908)
);

AO21x2_ASAP7_75t_L g909 ( 
.A1(n_735),
.A2(n_669),
.B(n_729),
.Y(n_909)
);

OA21x2_ASAP7_75t_L g910 ( 
.A1(n_735),
.A2(n_799),
.B(n_729),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_SL g911 ( 
.A1(n_733),
.A2(n_602),
.B1(n_588),
.B2(n_543),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_733),
.A2(n_830),
.B(n_807),
.Y(n_912)
);

AND2x6_ASAP7_75t_L g913 ( 
.A(n_743),
.B(n_805),
.Y(n_913)
);

BUFx8_ASAP7_75t_L g914 ( 
.A(n_763),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_733),
.A2(n_830),
.B(n_807),
.Y(n_915)
);

OA21x2_ASAP7_75t_L g916 ( 
.A1(n_735),
.A2(n_799),
.B(n_729),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_733),
.A2(n_777),
.B(n_651),
.Y(n_917)
);

NAND2xp33_ASAP7_75t_SL g918 ( 
.A(n_733),
.B(n_806),
.Y(n_918)
);

OA21x2_ASAP7_75t_L g919 ( 
.A1(n_735),
.A2(n_799),
.B(n_729),
.Y(n_919)
);

AO21x2_ASAP7_75t_L g920 ( 
.A1(n_735),
.A2(n_669),
.B(n_729),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_861),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_906),
.B(n_908),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_836),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_835),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_840),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_873),
.B(n_831),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_832),
.B(n_917),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_912),
.A2(n_915),
.B(n_833),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_841),
.Y(n_929)
);

NOR2x1_ASAP7_75t_SL g930 ( 
.A(n_832),
.B(n_882),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_843),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_891),
.B(n_834),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_844),
.Y(n_933)
);

INVxp33_ASAP7_75t_L g934 ( 
.A(n_863),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_846),
.B(n_853),
.Y(n_935)
);

AOI221xp5_ASAP7_75t_L g936 ( 
.A1(n_899),
.A2(n_911),
.B1(n_898),
.B2(n_904),
.C(n_918),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_871),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_846),
.Y(n_938)
);

O2A1O1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_872),
.A2(n_839),
.B(n_845),
.C(n_875),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_851),
.B(n_855),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_858),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_871),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_874),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_874),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_914),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_SL g946 ( 
.A1(n_838),
.A2(n_913),
.B1(n_896),
.B2(n_857),
.Y(n_946)
);

BUFx2_ASAP7_75t_R g947 ( 
.A(n_864),
.Y(n_947)
);

CKINVDCx20_ASAP7_75t_R g948 ( 
.A(n_837),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_889),
.B(n_890),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_893),
.B(n_860),
.Y(n_950)
);

CKINVDCx14_ASAP7_75t_R g951 ( 
.A(n_862),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_852),
.B(n_877),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_894),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_837),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_877),
.B(n_886),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_880),
.A2(n_895),
.B(n_909),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_879),
.Y(n_957)
);

AND2x4_ASAP7_75t_SL g958 ( 
.A(n_901),
.B(n_869),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_865),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_902),
.A2(n_903),
.B(n_887),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_884),
.B(n_850),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_842),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_907),
.Y(n_963)
);

OR2x2_ASAP7_75t_L g964 ( 
.A(n_878),
.B(n_881),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_SL g965 ( 
.A1(n_892),
.A2(n_854),
.B(n_859),
.C(n_888),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_909),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_905),
.B(n_848),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_897),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_885),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_920),
.B(n_883),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_876),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_910),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_916),
.B(n_919),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_870),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_856),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_868),
.B(n_867),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_866),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_849),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_900),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_847),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_933),
.B(n_938),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_940),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_935),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_923),
.B(n_925),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_931),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_957),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_941),
.B(n_946),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_946),
.B(n_953),
.Y(n_988)
);

INVx3_ASAP7_75t_SL g989 ( 
.A(n_924),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_936),
.B(n_926),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_959),
.Y(n_991)
);

INVx2_ASAP7_75t_SL g992 ( 
.A(n_932),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_937),
.B(n_942),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_937),
.B(n_942),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_943),
.B(n_944),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_963),
.B(n_927),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_960),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_927),
.B(n_952),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_967),
.B(n_928),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_966),
.B(n_972),
.Y(n_1000)
);

NOR2x1_ASAP7_75t_L g1001 ( 
.A(n_945),
.B(n_962),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_928),
.B(n_930),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_960),
.B(n_961),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_934),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_958),
.B(n_934),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_922),
.B(n_966),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_979),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_950),
.B(n_951),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_955),
.B(n_973),
.Y(n_1009)
);

OR2x2_ASAP7_75t_L g1010 ( 
.A(n_964),
.B(n_976),
.Y(n_1010)
);

OR2x2_ASAP7_75t_L g1011 ( 
.A(n_977),
.B(n_968),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_921),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_921),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_947),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_1002),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_1009),
.B(n_980),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_1003),
.B(n_970),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_985),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_984),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_1002),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_999),
.B(n_978),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_999),
.B(n_956),
.Y(n_1022)
);

BUFx2_ASAP7_75t_SL g1023 ( 
.A(n_992),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_982),
.B(n_939),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_1014),
.B(n_947),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_1006),
.B(n_956),
.Y(n_1026)
);

OR2x2_ASAP7_75t_L g1027 ( 
.A(n_1010),
.B(n_993),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_998),
.B(n_975),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_993),
.B(n_974),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_981),
.B(n_991),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_998),
.B(n_994),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_994),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_995),
.B(n_997),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_986),
.Y(n_1034)
);

NAND4xp25_ASAP7_75t_L g1035 ( 
.A(n_990),
.B(n_965),
.C(n_971),
.D(n_969),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_991),
.Y(n_1036)
);

NOR2xp67_ASAP7_75t_L g1037 ( 
.A(n_992),
.B(n_954),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_1004),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_1031),
.B(n_1005),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_1030),
.B(n_1005),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1034),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_1025),
.B(n_989),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1028),
.B(n_1021),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1018),
.Y(n_1044)
);

INVxp67_ASAP7_75t_L g1045 ( 
.A(n_1038),
.Y(n_1045)
);

OR2x2_ASAP7_75t_L g1046 ( 
.A(n_1027),
.B(n_996),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_1027),
.B(n_1032),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_1032),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_1033),
.B(n_1008),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1028),
.B(n_983),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_1029),
.B(n_1019),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1036),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1022),
.B(n_1007),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_1029),
.B(n_1000),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_1015),
.B(n_987),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_1015),
.B(n_1011),
.Y(n_1056)
);

OAI21xp33_ASAP7_75t_L g1057 ( 
.A1(n_1048),
.A2(n_1035),
.B(n_1024),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_1048),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1044),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_1052),
.Y(n_1060)
);

OR2x2_ASAP7_75t_L g1061 ( 
.A(n_1047),
.B(n_1026),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_1041),
.Y(n_1062)
);

OR2x2_ASAP7_75t_L g1063 ( 
.A(n_1043),
.B(n_1026),
.Y(n_1063)
);

NAND2x1_ASAP7_75t_L g1064 ( 
.A(n_1056),
.B(n_1020),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1054),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1045),
.B(n_1022),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_1039),
.B(n_1017),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1051),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_1049),
.Y(n_1069)
);

OR2x2_ASAP7_75t_L g1070 ( 
.A(n_1043),
.B(n_1016),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_1056),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_1040),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1062),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1066),
.B(n_1050),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_1058),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_1072),
.B(n_1055),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1062),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1063),
.B(n_1050),
.Y(n_1078)
);

OR2x2_ASAP7_75t_L g1079 ( 
.A(n_1061),
.B(n_1046),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_1057),
.A2(n_988),
.B(n_1014),
.C(n_1037),
.Y(n_1080)
);

OR2x2_ASAP7_75t_L g1081 ( 
.A(n_1070),
.B(n_1053),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1060),
.Y(n_1082)
);

OR2x6_ASAP7_75t_L g1083 ( 
.A(n_1064),
.B(n_1023),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1074),
.B(n_1058),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1076),
.B(n_1071),
.Y(n_1085)
);

AOI211x1_ASAP7_75t_L g1086 ( 
.A1(n_1078),
.A2(n_1065),
.B(n_1067),
.C(n_1068),
.Y(n_1086)
);

INVxp67_ASAP7_75t_L g1087 ( 
.A(n_1073),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1079),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1077),
.Y(n_1089)
);

OA21x2_ASAP7_75t_L g1090 ( 
.A1(n_1087),
.A2(n_1075),
.B(n_1082),
.Y(n_1090)
);

NAND4xp25_ASAP7_75t_L g1091 ( 
.A(n_1086),
.B(n_1080),
.C(n_1042),
.D(n_1075),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1088),
.B(n_1084),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_1091),
.B(n_924),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1092),
.B(n_1089),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1090),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1092),
.B(n_1069),
.Y(n_1096)
);

NOR3xp33_ASAP7_75t_SL g1097 ( 
.A(n_1093),
.B(n_989),
.C(n_948),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_1095),
.B(n_1085),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1098),
.B(n_1096),
.Y(n_1099)
);

NOR2x1_ASAP7_75t_L g1100 ( 
.A(n_1097),
.B(n_948),
.Y(n_1100)
);

NOR2x1p5_ASAP7_75t_L g1101 ( 
.A(n_1099),
.B(n_1094),
.Y(n_1101)
);

XNOR2x1_ASAP7_75t_L g1102 ( 
.A(n_1101),
.B(n_1100),
.Y(n_1102)
);

BUFx2_ASAP7_75t_L g1103 ( 
.A(n_1102),
.Y(n_1103)
);

OAI22x1_ASAP7_75t_L g1104 ( 
.A1(n_1103),
.A2(n_1001),
.B1(n_929),
.B2(n_949),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1104),
.A2(n_1083),
.B(n_965),
.Y(n_1105)
);

AOI21x1_ASAP7_75t_L g1106 ( 
.A1(n_1105),
.A2(n_1076),
.B(n_1059),
.Y(n_1106)
);

AO21x2_ASAP7_75t_L g1107 ( 
.A1(n_1106),
.A2(n_1067),
.B(n_1081),
.Y(n_1107)
);

OR2x2_ASAP7_75t_L g1108 ( 
.A(n_1107),
.B(n_1071),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1108),
.A2(n_1013),
.B(n_1012),
.Y(n_1109)
);


endmodule