module fake_jpeg_30499_n_472 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_472);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_472;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_18),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_77),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_7),
.B1(n_14),
.B2(n_2),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_50),
.A2(n_28),
.B1(n_39),
.B2(n_37),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_55),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_24),
.B(n_7),
.C(n_14),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_59),
.B(n_40),
.C(n_37),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_64),
.Y(n_125)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_66),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_18),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_81),
.Y(n_107)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_73),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_20),
.B(n_8),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_74),
.B(n_84),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_20),
.B(n_8),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_83),
.Y(n_102)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_42),
.B(n_5),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_86),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_87),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_89),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_26),
.B(n_5),
.Y(n_89)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_91),
.Y(n_118)
);

BUFx8_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_93),
.Y(n_127)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_26),
.B(n_5),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_27),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_27),
.B(n_10),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_28),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_93),
.A2(n_46),
.B1(n_30),
.B2(n_22),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_101),
.A2(n_114),
.B1(n_117),
.B2(n_134),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_104),
.B(n_113),
.Y(n_156)
);

CKINVDCx12_ASAP7_75t_R g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_106),
.B(n_122),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_73),
.A2(n_46),
.B1(n_30),
.B2(n_22),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_64),
.A2(n_46),
.B1(n_30),
.B2(n_22),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_79),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_51),
.A2(n_46),
.B1(n_22),
.B2(n_30),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_124),
.A2(n_130),
.B1(n_82),
.B2(n_80),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_56),
.B(n_32),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_137),
.Y(n_150)
);

HAxp5_ASAP7_75t_SL g128 ( 
.A(n_90),
.B(n_42),
.CON(n_128),
.SN(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_139),
.B(n_149),
.C(n_41),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_147),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_60),
.A2(n_33),
.B1(n_23),
.B2(n_34),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_70),
.A2(n_45),
.B1(n_31),
.B2(n_29),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_136),
.A2(n_145),
.B(n_13),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_61),
.B(n_32),
.Y(n_137)
);

HAxp5_ASAP7_75t_SL g139 ( 
.A(n_65),
.B(n_42),
.CON(n_139),
.SN(n_139)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_52),
.A2(n_33),
.B(n_34),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_52),
.B(n_45),
.Y(n_147)
);

NOR4xp25_ASAP7_75t_SL g149 ( 
.A(n_54),
.B(n_11),
.C(n_14),
.D(n_2),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_75),
.B1(n_88),
.B2(n_63),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_153),
.A2(n_166),
.B1(n_171),
.B2(n_103),
.Y(n_243)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_154),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_155),
.B(n_168),
.Y(n_206)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_157),
.Y(n_200)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_158),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_43),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_159),
.B(n_163),
.Y(n_230)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_161),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_128),
.A2(n_58),
.B1(n_139),
.B2(n_72),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_104),
.B(n_43),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_164),
.Y(n_208)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_165),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_134),
.A2(n_78),
.B1(n_68),
.B2(n_86),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_107),
.Y(n_167)
);

INVxp67_ASAP7_75t_SL g227 ( 
.A(n_167),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_107),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_169),
.Y(n_210)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_111),
.A2(n_137),
.B1(n_108),
.B2(n_136),
.Y(n_171)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_120),
.Y(n_173)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_127),
.A2(n_31),
.B1(n_39),
.B2(n_29),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_176),
.A2(n_178),
.B1(n_197),
.B2(n_169),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_125),
.A2(n_66),
.B1(n_55),
.B2(n_35),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_177),
.A2(n_182),
.B1(n_189),
.B2(n_196),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_110),
.A2(n_35),
.B1(n_19),
.B2(n_76),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_102),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_179),
.B(n_184),
.Y(n_207)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_180),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_96),
.B(n_67),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_195),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_125),
.A2(n_67),
.B1(n_87),
.B2(n_57),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_110),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_183),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_113),
.B(n_16),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_107),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_185),
.B(n_191),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_145),
.A2(n_49),
.B(n_91),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_190),
.B(n_123),
.Y(n_204)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_188),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_115),
.A2(n_16),
.B1(n_91),
.B2(n_19),
.Y(n_189)
);

O2A1O1Ixp33_ASAP7_75t_SL g190 ( 
.A1(n_118),
.A2(n_71),
.B(n_16),
.C(n_3),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_135),
.B(n_16),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_112),
.Y(n_192)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_132),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_193),
.Y(n_232)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_135),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_194),
.Y(n_236)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_112),
.Y(n_195)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_99),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_123),
.A2(n_16),
.B1(n_10),
.B2(n_3),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_148),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_198),
.Y(n_239)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_119),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_199),
.B(n_144),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_156),
.C(n_150),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_201),
.B(n_203),
.C(n_212),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_156),
.B(n_121),
.C(n_142),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_204),
.B(n_223),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_156),
.B(n_144),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_152),
.A2(n_105),
.B1(n_99),
.B2(n_132),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_215),
.A2(n_243),
.B1(n_198),
.B2(n_161),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_216),
.A2(n_173),
.B1(n_144),
.B2(n_120),
.Y(n_282)
);

NOR2x1_ASAP7_75t_L g218 ( 
.A(n_155),
.B(n_119),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_218),
.B(n_153),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_188),
.A2(n_105),
.B1(n_142),
.B2(n_103),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_234),
.B1(n_238),
.B2(n_169),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_150),
.B(n_16),
.Y(n_223)
);

OA22x2_ASAP7_75t_L g233 ( 
.A1(n_168),
.A2(n_146),
.B1(n_143),
.B2(n_131),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_233),
.B(n_241),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_167),
.A2(n_146),
.B1(n_143),
.B2(n_131),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_163),
.B(n_100),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_235),
.B(n_237),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_167),
.A2(n_146),
.B1(n_143),
.B2(n_131),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_159),
.B(n_191),
.Y(n_241)
);

AO21x2_ASAP7_75t_L g244 ( 
.A1(n_233),
.A2(n_186),
.B(n_190),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_244),
.A2(n_210),
.B1(n_243),
.B2(n_233),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_172),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_245),
.B(n_248),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_247),
.B(n_265),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_221),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_201),
.B(n_151),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_249),
.B(n_253),
.Y(n_289)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_251),
.Y(n_294)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_208),
.Y(n_252)
);

INVx3_ASAP7_75t_SL g315 ( 
.A(n_252),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_213),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_254),
.B(n_264),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_255),
.A2(n_279),
.B(n_277),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_212),
.B(n_160),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_256),
.B(n_231),
.C(n_223),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_194),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_257),
.B(n_276),
.Y(n_288)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_258),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_259),
.A2(n_260),
.B1(n_254),
.B2(n_239),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_214),
.A2(n_158),
.B1(n_198),
.B2(n_193),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_206),
.A2(n_180),
.B1(n_196),
.B2(n_187),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_262),
.A2(n_263),
.B1(n_269),
.B2(n_282),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_206),
.A2(n_154),
.B1(n_157),
.B2(n_170),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_213),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_205),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_205),
.Y(n_266)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_266),
.Y(n_304)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_224),
.Y(n_267)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_267),
.Y(n_306)
);

INVx8_ASAP7_75t_L g268 ( 
.A(n_208),
.Y(n_268)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_268),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_206),
.A2(n_164),
.B1(n_175),
.B2(n_195),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_230),
.B(n_235),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_270),
.B(n_271),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_230),
.B(n_174),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_224),
.Y(n_272)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_272),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_232),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_273),
.B(n_275),
.Y(n_310)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_220),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_274),
.Y(n_307)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_220),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_229),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_241),
.B(n_192),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_278),
.Y(n_298)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_222),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_222),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_281),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_207),
.B(n_165),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_250),
.A2(n_204),
.B(n_218),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_283),
.A2(n_293),
.B(n_311),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_284),
.A2(n_297),
.B1(n_303),
.B2(n_298),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_203),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_286),
.B(n_253),
.C(n_238),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_259),
.A2(n_202),
.B1(n_218),
.B2(n_216),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_287),
.A2(n_244),
.B1(n_262),
.B2(n_247),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_290),
.B(n_292),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_291),
.B(n_305),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_250),
.A2(n_202),
.B(n_240),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_250),
.A2(n_210),
.B(n_236),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_300),
.A2(n_308),
.B1(n_318),
.B2(n_280),
.Y(n_327)
);

FAx1_ASAP7_75t_SL g301 ( 
.A(n_261),
.B(n_257),
.CI(n_256),
.CON(n_301),
.SN(n_301)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_302),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_233),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_279),
.A2(n_223),
.B(n_227),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_255),
.A2(n_236),
.B1(n_228),
.B2(n_239),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_244),
.A2(n_217),
.B(n_242),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_232),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_312),
.B(n_313),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_273),
.B(n_209),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_265),
.Y(n_314)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_314),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_282),
.A2(n_228),
.B1(n_226),
.B2(n_209),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_319),
.A2(n_349),
.B1(n_297),
.B2(n_339),
.Y(n_356)
);

OA22x2_ASAP7_75t_L g320 ( 
.A1(n_284),
.A2(n_244),
.B1(n_269),
.B2(n_263),
.Y(n_320)
);

O2A1O1Ixp33_ASAP7_75t_L g362 ( 
.A1(n_320),
.A2(n_298),
.B(n_288),
.C(n_302),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_283),
.A2(n_244),
.B(n_260),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_322),
.A2(n_302),
.B(n_299),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_286),
.B(n_246),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_323),
.B(n_324),
.C(n_325),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_291),
.B(n_272),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_301),
.B(n_267),
.C(n_278),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_326),
.B(n_330),
.C(n_335),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_327),
.A2(n_345),
.B1(n_297),
.B2(n_311),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_313),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_328),
.B(n_340),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_301),
.B(n_275),
.C(n_274),
.Y(n_330)
);

BUFx24_ASAP7_75t_SL g332 ( 
.A(n_285),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_343),
.Y(n_354)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_310),
.Y(n_333)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_333),
.Y(n_365)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_310),
.Y(n_334)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_334),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_317),
.B(n_226),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_301),
.B(n_242),
.C(n_221),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_336),
.B(n_337),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_289),
.B(n_217),
.C(n_200),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_289),
.B(n_268),
.Y(n_338)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_338),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_287),
.A2(n_252),
.B1(n_200),
.B2(n_276),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_339),
.B(n_296),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_304),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_285),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_314),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_344),
.B(n_347),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_300),
.A2(n_258),
.B1(n_251),
.B2(n_229),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_312),
.Y(n_347)
);

OAI32xp33_ASAP7_75t_L g348 ( 
.A1(n_303),
.A2(n_120),
.A3(n_138),
.B1(n_100),
.B2(n_4),
.Y(n_348)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_348),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_353),
.A2(n_319),
.B1(n_302),
.B2(n_318),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_333),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_355),
.B(n_362),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_356),
.A2(n_373),
.B1(n_341),
.B2(n_322),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_321),
.B(n_317),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_357),
.B(n_363),
.Y(n_394)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_334),
.Y(n_359)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_359),
.Y(n_389)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_342),
.Y(n_361)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_361),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_321),
.B(n_290),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_342),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_364),
.B(n_375),
.Y(n_379)
);

INVx13_ASAP7_75t_L g368 ( 
.A(n_348),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_368),
.B(n_308),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_326),
.B(n_293),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_370),
.B(n_371),
.C(n_325),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_336),
.B(n_288),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_337),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_372),
.B(n_374),
.Y(n_398)
);

OAI21xp33_ASAP7_75t_L g373 ( 
.A1(n_346),
.A2(n_299),
.B(n_292),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_345),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_376),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_369),
.B(n_335),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_377),
.B(n_386),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_380),
.A2(n_381),
.B1(n_383),
.B2(n_391),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_351),
.A2(n_331),
.B1(n_327),
.B2(n_296),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_384),
.B(n_390),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_350),
.B(n_323),
.C(n_330),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_385),
.B(n_388),
.C(n_393),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_367),
.B(n_354),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_365),
.B(n_324),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_387),
.B(n_396),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_350),
.B(n_329),
.C(n_341),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_366),
.B(n_331),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_372),
.B(n_329),
.C(n_320),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_358),
.B(n_320),
.C(n_305),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_395),
.B(n_397),
.C(n_399),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_351),
.A2(n_304),
.B1(n_307),
.B2(n_320),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_358),
.B(n_307),
.C(n_316),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_352),
.B(n_316),
.C(n_306),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_383),
.A2(n_376),
.B1(n_356),
.B2(n_359),
.Y(n_402)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_402),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_379),
.Y(n_403)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_403),
.Y(n_423)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_389),
.Y(n_406)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_406),
.Y(n_428)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_382),
.Y(n_407)
);

AO221x1_ASAP7_75t_L g418 ( 
.A1(n_407),
.A2(n_414),
.B1(n_417),
.B2(n_309),
.C(n_294),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_382),
.A2(n_374),
.B(n_355),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_409),
.A2(n_411),
.B(n_138),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_378),
.A2(n_375),
.B1(n_361),
.B2(n_364),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_410),
.A2(n_416),
.B1(n_315),
.B2(n_294),
.Y(n_429)
);

A2O1A1Ixp33_ASAP7_75t_SL g411 ( 
.A1(n_380),
.A2(n_362),
.B(n_368),
.C(n_363),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_392),
.A2(n_371),
.B1(n_370),
.B2(n_360),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_413),
.B(n_295),
.Y(n_427)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_398),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_388),
.B(n_352),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_415),
.B(n_315),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_393),
.A2(n_357),
.B1(n_306),
.B2(n_309),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_398),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_418),
.B(n_425),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_408),
.B(n_399),
.C(n_397),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_419),
.B(n_420),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_408),
.B(n_385),
.C(n_384),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_404),
.B(n_395),
.C(n_394),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_421),
.B(n_424),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_404),
.B(n_415),
.C(n_401),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_409),
.A2(n_394),
.B(n_295),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_426),
.B(n_427),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_429),
.B(n_431),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_406),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_430),
.B(n_414),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_401),
.B(n_315),
.Y(n_431)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_432),
.Y(n_442)
);

OA21x2_ASAP7_75t_L g433 ( 
.A1(n_432),
.A2(n_407),
.B(n_417),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_433),
.B(n_445),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_435),
.B(n_444),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_422),
.A2(n_400),
.B(n_405),
.Y(n_438)
);

AO21x1_ASAP7_75t_L g446 ( 
.A1(n_438),
.A2(n_443),
.B(n_425),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_429),
.A2(n_405),
.B1(n_411),
.B2(n_413),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_439),
.A2(n_3),
.B1(n_4),
.B2(n_11),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_431),
.B(n_411),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_423),
.B(n_412),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_420),
.B(n_411),
.Y(n_445)
);

AO21x1_ASAP7_75t_L g459 ( 
.A1(n_446),
.A2(n_455),
.B(n_441),
.Y(n_459)
);

AOI322xp5_ASAP7_75t_L g447 ( 
.A1(n_438),
.A2(n_411),
.A3(n_428),
.B1(n_427),
.B2(n_426),
.C1(n_421),
.C2(n_419),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_447),
.A2(n_450),
.B1(n_436),
.B2(n_433),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_437),
.B(n_424),
.C(n_138),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_448),
.B(n_451),
.Y(n_457)
);

AOI31xp67_ASAP7_75t_SL g450 ( 
.A1(n_433),
.A2(n_100),
.A3(n_11),
.B(n_3),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_434),
.B(n_4),
.C(n_13),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_453),
.B(n_454),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_443),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_442),
.A2(n_435),
.B(n_436),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_456),
.B(n_458),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_452),
.B(n_439),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_459),
.A2(n_440),
.B(n_447),
.Y(n_463)
);

INVx13_ASAP7_75t_L g461 ( 
.A(n_449),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_461),
.B(n_462),
.Y(n_465)
);

INVxp33_ASAP7_75t_L g462 ( 
.A(n_449),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_463),
.B(n_461),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_457),
.A2(n_15),
.B(n_0),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_466),
.B(n_460),
.C(n_459),
.Y(n_468)
);

A2O1A1O1Ixp25_ASAP7_75t_L g470 ( 
.A1(n_467),
.A2(n_468),
.B(n_469),
.C(n_465),
.D(n_0),
.Y(n_470)
);

NOR2xp67_ASAP7_75t_SL g469 ( 
.A(n_464),
.B(n_0),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_470),
.B(n_1),
.C(n_450),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_471),
.B(n_1),
.Y(n_472)
);


endmodule