module fake_jpeg_12228_n_286 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_286);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_286;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_21),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_25),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_21),
.B(n_24),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_57),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_31),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_1),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_24),
.B(n_1),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_35),
.B(n_1),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_35),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_44),
.A2(n_27),
.B1(n_22),
.B2(n_20),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_71),
.A2(n_75),
.B1(n_25),
.B2(n_40),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_27),
.B1(n_22),
.B2(n_38),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_76),
.B(n_77),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_37),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_38),
.B1(n_36),
.B2(n_20),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_80),
.A2(n_86),
.B1(n_89),
.B2(n_40),
.Y(n_116)
);

AOI21xp33_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_19),
.B(n_39),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_103),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_63),
.A2(n_36),
.B1(n_20),
.B2(n_28),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_83),
.A2(n_40),
.B(n_25),
.Y(n_121)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_36),
.B1(n_28),
.B2(n_39),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_34),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_87),
.B(n_100),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_52),
.A2(n_26),
.B1(n_34),
.B2(n_33),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_41),
.A2(n_29),
.B1(n_33),
.B2(n_26),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_96),
.A2(n_8),
.B(n_9),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_98),
.Y(n_113)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_19),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_41),
.B(n_17),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_17),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_2),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_3),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_4),
.Y(n_123)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_73),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_110),
.B(n_123),
.Y(n_158)
);

NAND2x1_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_53),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_139),
.C(n_66),
.Y(n_148)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_114),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_3),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_69),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_116),
.B(n_129),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_89),
.A2(n_83),
.B1(n_67),
.B2(n_78),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_132),
.B1(n_93),
.B2(n_97),
.Y(n_154)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_121),
.A2(n_97),
.B(n_101),
.Y(n_157)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_67),
.A2(n_40),
.B1(n_25),
.B2(n_7),
.Y(n_132)
);

AO22x2_ASAP7_75t_L g133 ( 
.A1(n_85),
.A2(n_11),
.B1(n_6),
.B2(n_7),
.Y(n_133)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_82),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_136),
.B1(n_140),
.B2(n_72),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_92),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_70),
.Y(n_138)
);

NOR4xp25_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_74),
.C(n_70),
.D(n_69),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_92),
.B(n_9),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_65),
.A2(n_10),
.B1(n_66),
.B2(n_79),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_65),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

NOR3xp33_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_161),
.C(n_167),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_147),
.B(n_166),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_149),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_72),
.C(n_79),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_124),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_155),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_117),
.A2(n_111),
.B1(n_93),
.B2(n_127),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_152),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_123),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_172),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_156),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_120),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_157),
.A2(n_118),
.B1(n_130),
.B2(n_125),
.Y(n_190)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_168),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_121),
.A2(n_102),
.B(n_70),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_165),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_112),
.B(n_101),
.Y(n_166)
);

AOI32xp33_ASAP7_75t_L g167 ( 
.A1(n_127),
.A2(n_101),
.A3(n_102),
.B1(n_107),
.B2(n_111),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_109),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_169),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_129),
.A2(n_140),
.B1(n_136),
.B2(n_133),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_170),
.A2(n_132),
.B1(n_137),
.B2(n_114),
.Y(n_195)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_171),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_113),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_133),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_133),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_153),
.B(n_134),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_176),
.B(n_186),
.Y(n_212)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_164),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_182),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_164),
.Y(n_182)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_158),
.B(n_131),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_142),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_SL g222 ( 
.A1(n_190),
.A2(n_198),
.B(n_184),
.C(n_187),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_130),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_199),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_195),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_162),
.A2(n_160),
.B1(n_156),
.B2(n_173),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_197),
.Y(n_213)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_145),
.Y(n_197)
);

AO22x1_ASAP7_75t_SL g198 ( 
.A1(n_160),
.A2(n_108),
.B1(n_162),
.B2(n_154),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_172),
.B(n_149),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_148),
.B(n_165),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_201),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_151),
.B(n_144),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_183),
.A2(n_144),
.B(n_157),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_211),
.Y(n_231)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_178),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_210),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_194),
.A2(n_161),
.B(n_162),
.Y(n_208)
);

OAI22x1_ASAP7_75t_L g240 ( 
.A1(n_208),
.A2(n_222),
.B1(n_216),
.B2(n_218),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_151),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_191),
.Y(n_211)
);

OA21x2_ASAP7_75t_L g214 ( 
.A1(n_196),
.A2(n_146),
.B(n_163),
.Y(n_214)
);

OA21x2_ASAP7_75t_L g238 ( 
.A1(n_214),
.A2(n_213),
.B(n_222),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_146),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_217),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_181),
.A2(n_166),
.B(n_188),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_192),
.Y(n_218)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_218),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_184),
.Y(n_220)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_175),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_223),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_179),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_214),
.A2(n_184),
.B1(n_188),
.B2(n_190),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_221),
.B(n_181),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_228),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_181),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_214),
.A2(n_195),
.B1(n_198),
.B2(n_185),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_229),
.A2(n_237),
.B1(n_222),
.B2(n_219),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_202),
.A2(n_174),
.B1(n_177),
.B2(n_197),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_232),
.A2(n_233),
.B1(n_238),
.B2(n_216),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_202),
.A2(n_174),
.B1(n_177),
.B2(n_182),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_209),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_239),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_211),
.A2(n_213),
.B1(n_220),
.B2(n_223),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_204),
.C(n_222),
.Y(n_239)
);

AO21x1_ASAP7_75t_L g250 ( 
.A1(n_240),
.A2(n_222),
.B(n_203),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_241),
.A2(n_238),
.B1(n_239),
.B2(n_205),
.Y(n_261)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_243),
.Y(n_256)
);

AO21x1_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_250),
.B(n_240),
.Y(n_253)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_246),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_212),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_247),
.Y(n_257)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_251),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_253),
.A2(n_261),
.B1(n_248),
.B2(n_238),
.Y(n_267)
);

XOR2x2_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_227),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_254),
.A2(n_235),
.B(n_236),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_244),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_257),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_228),
.Y(n_262)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_241),
.C(n_250),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_262),
.B(n_249),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_264),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_249),
.Y(n_264)
);

OAI221xp5_ASAP7_75t_L g271 ( 
.A1(n_265),
.A2(n_266),
.B1(n_253),
.B2(n_259),
.C(n_255),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_267),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_248),
.C(n_207),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_270),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_205),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_269),
.B(n_258),
.Y(n_272)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_271),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_264),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_263),
.B(n_268),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_276),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_278),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_266),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_280),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_279),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_281),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_277),
.B(n_274),
.Y(n_285)
);

XNOR2x2_ASAP7_75t_SL g286 ( 
.A(n_285),
.B(n_274),
.Y(n_286)
);


endmodule