module fake_aes_424_n_21 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_21);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_21;
wire n_20;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
INVx1_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_1), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_4), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_5), .Y(n_11) );
INVx3_ASAP7_75t_L g12 ( .A(n_2), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_10), .Y(n_14) );
AO21x2_ASAP7_75t_L g15 ( .A1(n_13), .A2(n_11), .B(n_9), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_15), .B(n_14), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_16), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
CKINVDCx16_ASAP7_75t_R g19 ( .A(n_18), .Y(n_19) );
OR2x6_ASAP7_75t_L g20 ( .A(n_19), .B(n_12), .Y(n_20) );
AOI22xp5_ASAP7_75t_SL g21 ( .A1(n_20), .A2(n_0), .B1(n_3), .B2(n_6), .Y(n_21) );
endmodule