module fake_netlist_6_3638_n_757 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_757);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_757;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_698;
wire n_617;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_685;
wire n_597;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_746;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_720;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_683;
wire n_420;
wire n_620;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_92),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_137),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_59),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_48),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_34),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_126),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_123),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_49),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_29),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_5),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_18),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_148),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_107),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_27),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_112),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_89),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_91),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_62),
.Y(n_169)
);

HB1xp67_ASAP7_75t_SL g170 ( 
.A(n_71),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_72),
.Y(n_171)
);

CKINVDCx11_ASAP7_75t_R g172 ( 
.A(n_26),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_60),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_101),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_11),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_4),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_76),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_149),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_1),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_73),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_35),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_0),
.Y(n_182)
);

BUFx8_ASAP7_75t_SL g183 ( 
.A(n_38),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_63),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_67),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_55),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_150),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_7),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_20),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_50),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_80),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_78),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_44),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_51),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_40),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_118),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_114),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_7),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_85),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_77),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_125),
.B(n_132),
.Y(n_203)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_154),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_161),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_158),
.B(n_0),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_1),
.Y(n_208)
);

BUFx8_ASAP7_75t_SL g209 ( 
.A(n_183),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_175),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_154),
.Y(n_211)
);

INVxp33_ASAP7_75t_SL g212 ( 
.A(n_159),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_156),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_174),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

OA21x2_ASAP7_75t_L g217 ( 
.A1(n_166),
.A2(n_2),
.B(n_3),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_5),
.Y(n_220)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_151),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_157),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_152),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_184),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_6),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_189),
.A2(n_200),
.B1(n_170),
.B2(n_182),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_167),
.B(n_6),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_153),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_155),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_160),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g236 ( 
.A(n_172),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_162),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_163),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_155),
.A2(n_164),
.B1(n_169),
.B2(n_186),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_165),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_171),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_178),
.Y(n_242)
);

OA21x2_ASAP7_75t_L g243 ( 
.A1(n_168),
.A2(n_8),
.B(n_9),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_209),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_205),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_209),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_216),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_205),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_236),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_236),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_240),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_R g252 ( 
.A(n_235),
.B(n_199),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_240),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_214),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_214),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_216),
.Y(n_256)
);

AOI21x1_ASAP7_75t_L g257 ( 
.A1(n_219),
.A2(n_192),
.B(n_201),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_240),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_211),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_240),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_240),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_211),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_221),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_221),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_221),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_239),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_223),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_216),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_214),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_223),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_214),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_218),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_226),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_223),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_235),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_R g276 ( 
.A(n_235),
.B(n_202),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_241),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_241),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_241),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_228),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_228),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_212),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_229),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_216),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_215),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_212),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_238),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_233),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_233),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_237),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_251),
.B(n_237),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_216),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_283),
.B(n_164),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_288),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_256),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_256),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_290),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_247),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_242),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_253),
.B(n_242),
.Y(n_300)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_247),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_268),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_254),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_204),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_260),
.B(n_204),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_255),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_268),
.B(n_204),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_247),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_261),
.B(n_204),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_275),
.B(n_227),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_247),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_287),
.A2(n_243),
.B1(n_217),
.B2(n_220),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_280),
.B(n_204),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_282),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_269),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_283),
.A2(n_243),
.B1(n_217),
.B2(n_208),
.Y(n_316)
);

NAND2xp33_ASAP7_75t_L g317 ( 
.A(n_277),
.B(n_207),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_278),
.B(n_215),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_252),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_276),
.B(n_231),
.Y(n_320)
);

INVx4_ASAP7_75t_SL g321 ( 
.A(n_271),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_281),
.B(n_224),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_279),
.B(n_224),
.Y(n_323)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_245),
.Y(n_324)
);

NAND3xp33_ASAP7_75t_L g325 ( 
.A(n_263),
.B(n_230),
.C(n_213),
.Y(n_325)
);

NOR3xp33_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_234),
.C(n_215),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_264),
.B(n_222),
.Y(n_327)
);

NAND2xp33_ASAP7_75t_L g328 ( 
.A(n_265),
.B(n_180),
.Y(n_328)
);

OR2x6_ASAP7_75t_L g329 ( 
.A(n_244),
.B(n_206),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_257),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_L g331 ( 
.A(n_267),
.B(n_224),
.Y(n_331)
);

NOR3xp33_ASAP7_75t_L g332 ( 
.A(n_270),
.B(n_193),
.C(n_232),
.Y(n_332)
);

OA21x2_ASAP7_75t_L g333 ( 
.A1(n_249),
.A2(n_219),
.B(n_206),
.Y(n_333)
);

NOR2xp67_ASAP7_75t_SL g334 ( 
.A(n_250),
.B(n_217),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_272),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_274),
.Y(n_336)
);

NAND2xp33_ASAP7_75t_L g337 ( 
.A(n_273),
.B(n_181),
.Y(n_337)
);

OR2x6_ASAP7_75t_L g338 ( 
.A(n_246),
.B(n_210),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_266),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_262),
.B(n_225),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_248),
.A2(n_243),
.B1(n_225),
.B2(n_210),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_259),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_247),
.Y(n_343)
);

BUFx6f_ASAP7_75t_SL g344 ( 
.A(n_254),
.Y(n_344)
);

NOR3xp33_ASAP7_75t_L g345 ( 
.A(n_285),
.B(n_203),
.C(n_187),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_288),
.B(n_225),
.Y(n_346)
);

OA21x2_ASAP7_75t_L g347 ( 
.A1(n_284),
.A2(n_197),
.B(n_194),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_254),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_285),
.B(n_169),
.Y(n_349)
);

NOR3xp33_ASAP7_75t_L g350 ( 
.A(n_285),
.B(n_188),
.C(n_190),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_254),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_256),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_285),
.B(n_225),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_285),
.B(n_186),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_295),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_293),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_296),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_298),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_302),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_316),
.B(n_17),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_292),
.Y(n_361)
);

OAI22xp33_ASAP7_75t_L g362 ( 
.A1(n_323),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_353),
.B(n_12),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_352),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_292),
.Y(n_365)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_343),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_310),
.B(n_19),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_343),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_346),
.B(n_21),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_323),
.B(n_22),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_319),
.Y(n_371)
);

AND2x6_ASAP7_75t_L g372 ( 
.A(n_330),
.B(n_23),
.Y(n_372)
);

NOR3xp33_ASAP7_75t_SL g373 ( 
.A(n_325),
.B(n_13),
.C(n_14),
.Y(n_373)
);

OR2x6_ASAP7_75t_L g374 ( 
.A(n_342),
.B(n_329),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_297),
.B(n_13),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_298),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_291),
.B(n_24),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_343),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_326),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_300),
.B(n_331),
.Y(n_380)
);

OR2x6_ASAP7_75t_L g381 ( 
.A(n_329),
.B(n_15),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_333),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_294),
.B(n_16),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_303),
.B(n_306),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_L g385 ( 
.A1(n_312),
.A2(n_25),
.B1(n_28),
.B2(n_30),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_299),
.B(n_31),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_341),
.B(n_32),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_322),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_322),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_333),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_340),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_309),
.A2(n_305),
.B(n_304),
.Y(n_392)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_329),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_315),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_318),
.B(n_33),
.Y(n_395)
);

BUFx4f_ASAP7_75t_L g396 ( 
.A(n_336),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_309),
.B(n_36),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_348),
.B(n_37),
.Y(n_398)
);

NOR3xp33_ASAP7_75t_SL g399 ( 
.A(n_349),
.B(n_39),
.C(n_41),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_351),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_350),
.B(n_42),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_327),
.B(n_43),
.Y(n_402)
);

BUFx8_ASAP7_75t_L g403 ( 
.A(n_339),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_317),
.B(n_45),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_308),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_311),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_320),
.B(n_46),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_332),
.B(n_47),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_334),
.B(n_52),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_321),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_347),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_354),
.Y(n_412)
);

NOR2xp67_ASAP7_75t_L g413 ( 
.A(n_313),
.B(n_53),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_335),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_345),
.B(n_54),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_313),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_344),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_328),
.B(n_56),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_335),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_338),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_347),
.B(n_57),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_388),
.B(n_307),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_380),
.A2(n_307),
.B(n_301),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_391),
.B(n_419),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_356),
.B(n_414),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_SL g426 ( 
.A1(n_375),
.A2(n_293),
.B1(n_337),
.B2(n_314),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_371),
.B(n_324),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_384),
.B(n_338),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_412),
.B(n_321),
.Y(n_429)
);

AOI21x1_ASAP7_75t_L g430 ( 
.A1(n_370),
.A2(n_338),
.B(n_321),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_392),
.A2(n_301),
.B(n_344),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_400),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_389),
.B(n_301),
.Y(n_433)
);

INVx2_ASAP7_75t_SL g434 ( 
.A(n_396),
.Y(n_434)
);

A2O1A1Ixp33_ASAP7_75t_L g435 ( 
.A1(n_360),
.A2(n_301),
.B(n_61),
.C(n_64),
.Y(n_435)
);

AOI22xp33_ASAP7_75t_L g436 ( 
.A1(n_360),
.A2(n_58),
.B1(n_65),
.B2(n_66),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_416),
.B(n_68),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_387),
.A2(n_69),
.B(n_70),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_361),
.B(n_74),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_382),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_355),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g442 ( 
.A(n_420),
.B(n_75),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_382),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_385),
.A2(n_387),
.B1(n_379),
.B2(n_367),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_384),
.B(n_79),
.Y(n_445)
);

NOR3xp33_ASAP7_75t_L g446 ( 
.A(n_383),
.B(n_81),
.C(n_82),
.Y(n_446)
);

O2A1O1Ixp33_ASAP7_75t_L g447 ( 
.A1(n_363),
.A2(n_83),
.B(n_84),
.C(n_86),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_403),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_407),
.A2(n_88),
.B1(n_90),
.B2(n_93),
.Y(n_449)
);

OA22x2_ASAP7_75t_L g450 ( 
.A1(n_379),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_382),
.Y(n_451)
);

OAI21x1_ASAP7_75t_L g452 ( 
.A1(n_411),
.A2(n_97),
.B(n_98),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_358),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_365),
.A2(n_99),
.B(n_100),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_358),
.Y(n_455)
);

A2O1A1Ixp33_ASAP7_75t_L g456 ( 
.A1(n_377),
.A2(n_390),
.B(n_404),
.C(n_411),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_366),
.A2(n_102),
.B(n_103),
.Y(n_457)
);

NAND2x1p5_ASAP7_75t_L g458 ( 
.A(n_410),
.B(n_104),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_374),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_366),
.A2(n_105),
.B(n_106),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_396),
.B(n_108),
.Y(n_461)
);

A2O1A1Ixp33_ASAP7_75t_L g462 ( 
.A1(n_369),
.A2(n_109),
.B(n_110),
.C(n_111),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_357),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_397),
.A2(n_421),
.B(n_409),
.Y(n_464)
);

AOI221xp5_ASAP7_75t_L g465 ( 
.A1(n_362),
.A2(n_113),
.B1(n_115),
.B2(n_116),
.C(n_117),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_418),
.A2(n_119),
.B(n_120),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_359),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_393),
.B(n_401),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_401),
.B(n_121),
.Y(n_469)
);

O2A1O1Ixp33_ASAP7_75t_L g470 ( 
.A1(n_408),
.A2(n_122),
.B(n_124),
.C(n_127),
.Y(n_470)
);

INVx3_ASAP7_75t_SL g471 ( 
.A(n_374),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_364),
.Y(n_472)
);

NAND2xp33_ASAP7_75t_L g473 ( 
.A(n_372),
.B(n_128),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_374),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_417),
.B(n_129),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_395),
.B(n_130),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_425),
.Y(n_477)
);

OAI21x1_ASAP7_75t_L g478 ( 
.A1(n_452),
.A2(n_398),
.B(n_376),
.Y(n_478)
);

AO21x2_ASAP7_75t_L g479 ( 
.A1(n_456),
.A2(n_464),
.B(n_444),
.Y(n_479)
);

CKINVDCx6p67_ASAP7_75t_R g480 ( 
.A(n_471),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_440),
.Y(n_481)
);

OAI21x1_ASAP7_75t_L g482 ( 
.A1(n_423),
.A2(n_376),
.B(n_405),
.Y(n_482)
);

BUFx2_ASAP7_75t_SL g483 ( 
.A(n_424),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_459),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_432),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_443),
.Y(n_486)
);

INVx6_ASAP7_75t_L g487 ( 
.A(n_445),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_451),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_453),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_441),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_467),
.Y(n_491)
);

OAI21x1_ASAP7_75t_L g492 ( 
.A1(n_431),
.A2(n_406),
.B(n_378),
.Y(n_492)
);

OR2x6_ASAP7_75t_L g493 ( 
.A(n_445),
.B(n_402),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_453),
.Y(n_494)
);

NAND2x1p5_ASAP7_75t_L g495 ( 
.A(n_455),
.B(n_415),
.Y(n_495)
);

AO21x2_ASAP7_75t_L g496 ( 
.A1(n_444),
.A2(n_386),
.B(n_399),
.Y(n_496)
);

INVx5_ASAP7_75t_L g497 ( 
.A(n_455),
.Y(n_497)
);

BUFx10_ASAP7_75t_L g498 ( 
.A(n_461),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_422),
.A2(n_413),
.B(n_394),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_476),
.A2(n_413),
.B(n_372),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_463),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_472),
.Y(n_502)
);

BUFx4f_ASAP7_75t_L g503 ( 
.A(n_458),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_422),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_439),
.Y(n_505)
);

INVx6_ASAP7_75t_L g506 ( 
.A(n_442),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_450),
.Y(n_507)
);

BUFx12f_ASAP7_75t_L g508 ( 
.A(n_428),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_434),
.B(n_403),
.Y(n_509)
);

NAND2x1p5_ASAP7_75t_L g510 ( 
.A(n_469),
.B(n_368),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_458),
.Y(n_511)
);

OR2x6_ASAP7_75t_L g512 ( 
.A(n_468),
.B(n_381),
.Y(n_512)
);

OA21x2_ASAP7_75t_L g513 ( 
.A1(n_438),
.A2(n_373),
.B(n_372),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_428),
.B(n_372),
.Y(n_514)
);

OA21x2_ASAP7_75t_L g515 ( 
.A1(n_438),
.A2(n_368),
.B(n_381),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_437),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_474),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g518 ( 
.A1(n_476),
.A2(n_430),
.B(n_454),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_433),
.Y(n_519)
);

AOI22x1_ASAP7_75t_L g520 ( 
.A1(n_466),
.A2(n_368),
.B1(n_381),
.B2(n_134),
.Y(n_520)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_457),
.A2(n_131),
.B(n_133),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_SL g522 ( 
.A1(n_473),
.A2(n_426),
.B1(n_475),
.B2(n_448),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_485),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_508),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_477),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_478),
.A2(n_460),
.B(n_447),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_497),
.Y(n_527)
);

BUFx6f_ASAP7_75t_SL g528 ( 
.A(n_514),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_497),
.Y(n_529)
);

BUFx12f_ASAP7_75t_L g530 ( 
.A(n_508),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_504),
.Y(n_531)
);

AO21x1_ASAP7_75t_L g532 ( 
.A1(n_516),
.A2(n_470),
.B(n_446),
.Y(n_532)
);

CKINVDCx11_ASAP7_75t_R g533 ( 
.A(n_480),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_517),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_501),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_501),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_481),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_507),
.B(n_465),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_481),
.Y(n_539)
);

OR2x2_ASAP7_75t_L g540 ( 
.A(n_515),
.B(n_427),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_488),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_490),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_491),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_488),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_502),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_494),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_494),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_484),
.Y(n_548)
);

CKINVDCx11_ASAP7_75t_R g549 ( 
.A(n_480),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_483),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_483),
.Y(n_551)
);

AO21x1_ASAP7_75t_SL g552 ( 
.A1(n_499),
.A2(n_436),
.B(n_449),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_486),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_486),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_517),
.Y(n_555)
);

NAND2x1p5_ASAP7_75t_L g556 ( 
.A(n_503),
.B(n_429),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_522),
.A2(n_513),
.B1(n_493),
.B2(n_514),
.Y(n_557)
);

INVx6_ASAP7_75t_L g558 ( 
.A(n_497),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_515),
.B(n_435),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_486),
.Y(n_560)
);

OAI21x1_ASAP7_75t_L g561 ( 
.A1(n_478),
.A2(n_462),
.B(n_136),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_515),
.B(n_135),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_513),
.B(n_138),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_R g564 ( 
.A(n_533),
.B(n_509),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_558),
.Y(n_565)
);

OR2x6_ASAP7_75t_L g566 ( 
.A(n_558),
.B(n_487),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_558),
.Y(n_567)
);

NAND2xp33_ASAP7_75t_R g568 ( 
.A(n_562),
.B(n_514),
.Y(n_568)
);

NAND2xp33_ASAP7_75t_R g569 ( 
.A(n_562),
.B(n_513),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_523),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_525),
.B(n_512),
.Y(n_571)
);

NAND3xp33_ASAP7_75t_L g572 ( 
.A(n_538),
.B(n_520),
.C(n_493),
.Y(n_572)
);

NAND2xp33_ASAP7_75t_L g573 ( 
.A(n_550),
.B(n_551),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_523),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_542),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_543),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_531),
.B(n_519),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_534),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_548),
.B(n_512),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_534),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_538),
.A2(n_493),
.B1(n_496),
.B2(n_512),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_555),
.B(n_512),
.Y(n_582)
);

CKINVDCx16_ASAP7_75t_R g583 ( 
.A(n_530),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_531),
.B(n_493),
.Y(n_584)
);

INVxp67_ASAP7_75t_L g585 ( 
.A(n_555),
.Y(n_585)
);

NOR2xp67_ASAP7_75t_R g586 ( 
.A(n_558),
.B(n_506),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_545),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_524),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_540),
.B(n_487),
.Y(n_589)
);

AND2x4_ASAP7_75t_SL g590 ( 
.A(n_527),
.B(n_498),
.Y(n_590)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_540),
.B(n_510),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_541),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_546),
.B(n_487),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_524),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_535),
.B(n_510),
.Y(n_595)
);

O2A1O1Ixp33_ASAP7_75t_SL g596 ( 
.A1(n_535),
.A2(n_519),
.B(n_511),
.C(n_505),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_549),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_547),
.B(n_487),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_L g599 ( 
.A1(n_559),
.A2(n_505),
.B(n_492),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_557),
.A2(n_506),
.B1(n_503),
.B2(n_510),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_530),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_536),
.B(n_489),
.Y(n_602)
);

OA21x2_ASAP7_75t_L g603 ( 
.A1(n_526),
.A2(n_518),
.B(n_482),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_R g604 ( 
.A(n_563),
.B(n_511),
.Y(n_604)
);

NAND2xp33_ASAP7_75t_R g605 ( 
.A(n_563),
.B(n_489),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_536),
.Y(n_606)
);

NOR2x1p5_ASAP7_75t_L g607 ( 
.A(n_547),
.B(n_489),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_532),
.A2(n_479),
.B(n_503),
.Y(n_608)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_537),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_589),
.B(n_559),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_570),
.Y(n_611)
);

NAND2x1p5_ASAP7_75t_L g612 ( 
.A(n_565),
.B(n_527),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_574),
.B(n_544),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_591),
.B(n_544),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_584),
.B(n_539),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_575),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_580),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_606),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_592),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_580),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_576),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_587),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_609),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_571),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_599),
.B(n_554),
.Y(n_625)
);

AND2x4_ASAP7_75t_SL g626 ( 
.A(n_580),
.B(n_498),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_599),
.B(n_554),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_577),
.Y(n_628)
);

AOI221xp5_ASAP7_75t_L g629 ( 
.A1(n_572),
.A2(n_496),
.B1(n_532),
.B2(n_479),
.C(n_528),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_579),
.B(n_498),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_581),
.B(n_496),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_595),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_573),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_602),
.B(n_560),
.Y(n_634)
);

INVx5_ASAP7_75t_L g635 ( 
.A(n_566),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_608),
.B(n_561),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_578),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_602),
.B(n_553),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_600),
.B(n_561),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_600),
.B(n_495),
.Y(n_640)
);

NAND3xp33_ASAP7_75t_SL g641 ( 
.A(n_564),
.B(n_495),
.C(n_556),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_596),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_598),
.B(n_529),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_641),
.A2(n_572),
.B1(n_568),
.B2(n_528),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_614),
.B(n_582),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_614),
.B(n_582),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_633),
.B(n_585),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_611),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_616),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_621),
.Y(n_650)
);

NAND3xp33_ASAP7_75t_L g651 ( 
.A(n_629),
.B(n_630),
.C(n_623),
.Y(n_651)
);

NAND2x1_ASAP7_75t_SL g652 ( 
.A(n_637),
.B(n_624),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_622),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_610),
.B(n_603),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_618),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_618),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_632),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_610),
.B(n_603),
.Y(n_658)
);

NAND2xp33_ASAP7_75t_L g659 ( 
.A(n_635),
.B(n_588),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_632),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_615),
.B(n_594),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_613),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_631),
.B(n_593),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_615),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_631),
.B(n_607),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_619),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_613),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_625),
.B(n_590),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_628),
.B(n_586),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_626),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_655),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_651),
.A2(n_552),
.B1(n_640),
.B2(n_528),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_654),
.B(n_625),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_663),
.B(n_627),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_644),
.A2(n_552),
.B1(n_640),
.B2(n_506),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_663),
.B(n_627),
.Y(n_676)
);

INVxp67_ASAP7_75t_L g677 ( 
.A(n_647),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_654),
.B(n_636),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_655),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_666),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_666),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_670),
.Y(n_682)
);

INVx1_ASAP7_75t_SL g683 ( 
.A(n_652),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_648),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_664),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_658),
.B(n_639),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_684),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_677),
.A2(n_647),
.B1(n_635),
.B2(n_646),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_679),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_674),
.B(n_657),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_684),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_685),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_672),
.A2(n_659),
.B1(n_604),
.B2(n_665),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_676),
.B(n_660),
.Y(n_694)
);

OAI21xp33_ASAP7_75t_L g695 ( 
.A1(n_675),
.A2(n_669),
.B(n_665),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_671),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_673),
.B(n_658),
.Y(n_697)
);

AOI21xp33_ASAP7_75t_SL g698 ( 
.A1(n_688),
.A2(n_583),
.B(n_597),
.Y(n_698)
);

OAI21xp33_ASAP7_75t_L g699 ( 
.A1(n_695),
.A2(n_683),
.B(n_678),
.Y(n_699)
);

AO21x1_ASAP7_75t_L g700 ( 
.A1(n_688),
.A2(n_659),
.B(n_649),
.Y(n_700)
);

NAND4xp75_ASAP7_75t_L g701 ( 
.A(n_693),
.B(n_650),
.C(n_653),
.D(n_668),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_692),
.A2(n_683),
.B1(n_682),
.B2(n_668),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_699),
.B(n_697),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_698),
.B(n_601),
.Y(n_704)
);

OAI21xp5_ASAP7_75t_L g705 ( 
.A1(n_701),
.A2(n_694),
.B(n_690),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_702),
.B(n_691),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_700),
.B(n_678),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_706),
.Y(n_708)
);

INVx1_ASAP7_75t_SL g709 ( 
.A(n_707),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_705),
.B(n_687),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_703),
.B(n_673),
.Y(n_711)
);

AOI211x1_ASAP7_75t_L g712 ( 
.A1(n_710),
.A2(n_708),
.B(n_711),
.C(n_709),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_708),
.B(n_704),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_711),
.Y(n_714)
);

OAI211xp5_ASAP7_75t_SL g715 ( 
.A1(n_713),
.A2(n_696),
.B(n_645),
.C(n_689),
.Y(n_715)
);

AOI222xp33_ASAP7_75t_SL g716 ( 
.A1(n_714),
.A2(n_679),
.B1(n_671),
.B2(n_681),
.C1(n_642),
.C2(n_667),
.Y(n_716)
);

AOI321xp33_ASAP7_75t_L g717 ( 
.A1(n_712),
.A2(n_661),
.A3(n_682),
.B1(n_638),
.B2(n_670),
.C(n_643),
.Y(n_717)
);

AOI211xp5_ASAP7_75t_L g718 ( 
.A1(n_713),
.A2(n_588),
.B(n_620),
.C(n_617),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_717),
.Y(n_719)
);

NOR2x1_ASAP7_75t_L g720 ( 
.A(n_715),
.B(n_588),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_718),
.B(n_686),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_716),
.A2(n_626),
.B1(n_620),
.B2(n_617),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_718),
.B(n_686),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_717),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_718),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_719),
.A2(n_605),
.B1(n_569),
.B2(n_638),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_721),
.Y(n_727)
);

NOR3xp33_ASAP7_75t_L g728 ( 
.A(n_725),
.B(n_565),
.C(n_567),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_723),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_720),
.Y(n_730)
);

AND3x4_ASAP7_75t_L g731 ( 
.A(n_724),
.B(n_680),
.C(n_619),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_722),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_729),
.B(n_679),
.Y(n_733)
);

NOR4xp25_ASAP7_75t_SL g734 ( 
.A(n_732),
.B(n_656),
.C(n_586),
.D(n_662),
.Y(n_734)
);

NAND4xp75_ASAP7_75t_L g735 ( 
.A(n_726),
.B(n_139),
.C(n_141),
.D(n_142),
.Y(n_735)
);

BUFx10_ASAP7_75t_L g736 ( 
.A(n_727),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_727),
.B(n_681),
.Y(n_737)
);

NAND2xp33_ASAP7_75t_L g738 ( 
.A(n_730),
.B(n_612),
.Y(n_738)
);

INVx3_ASAP7_75t_SL g739 ( 
.A(n_728),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_739),
.A2(n_731),
.B1(n_681),
.B2(n_680),
.Y(n_740)
);

INVx1_ASAP7_75t_SL g741 ( 
.A(n_736),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_733),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_737),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_738),
.A2(n_634),
.B1(n_643),
.B2(n_506),
.Y(n_744)
);

AND2x2_ASAP7_75t_SL g745 ( 
.A(n_742),
.B(n_735),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_741),
.A2(n_734),
.B1(n_735),
.B2(n_635),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_743),
.Y(n_747)
);

OA22x2_ASAP7_75t_L g748 ( 
.A1(n_744),
.A2(n_567),
.B1(n_566),
.B2(n_634),
.Y(n_748)
);

XNOR2xp5_ASAP7_75t_L g749 ( 
.A(n_745),
.B(n_740),
.Y(n_749)
);

BUFx2_ASAP7_75t_L g750 ( 
.A(n_747),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_748),
.A2(n_635),
.B1(n_612),
.B2(n_566),
.Y(n_751)
);

OAI21xp5_ASAP7_75t_L g752 ( 
.A1(n_749),
.A2(n_746),
.B(n_556),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_750),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_753),
.B(n_751),
.Y(n_754)
);

AOI222xp33_ASAP7_75t_L g755 ( 
.A1(n_754),
.A2(n_752),
.B1(n_521),
.B2(n_635),
.C1(n_497),
.C2(n_500),
.Y(n_755)
);

AOI221xp5_ASAP7_75t_SL g756 ( 
.A1(n_755),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.C(n_147),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_756),
.A2(n_556),
.B1(n_495),
.B2(n_521),
.Y(n_757)
);


endmodule