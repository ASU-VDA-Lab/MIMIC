module fake_jpeg_13810_n_429 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_429);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_429;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_2),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_7),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_56),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_57),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_58),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_16),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_59),
.B(n_63),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_60),
.Y(n_178)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_61),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_62),
.B(n_73),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_0),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_65),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx4f_ASAP7_75t_SL g169 ( 
.A(n_66),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_32),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_67),
.B(n_68),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_55),
.B(n_1),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_69),
.Y(n_153)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_71),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_32),
.B(n_3),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_72),
.B(n_88),
.Y(n_172)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_74),
.Y(n_161)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_75),
.Y(n_165)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_78),
.B(n_80),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx5_ASAP7_75t_SL g154 ( 
.A(n_79),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_19),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_81),
.B(n_86),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_20),
.B(n_3),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_82),
.B(n_5),
.Y(n_140)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_24),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_98),
.Y(n_114)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_19),
.Y(n_86)
);

BUFx16f_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_87),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_3),
.Y(n_88)
);

BUFx10_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_91),
.B(n_95),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_94),
.Y(n_171)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_49),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_99),
.B(n_100),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_49),
.Y(n_100)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_101),
.B(n_110),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

NAND2xp33_ASAP7_75t_SL g127 ( 
.A(n_102),
.B(n_103),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

NAND2xp33_ASAP7_75t_SL g166 ( 
.A(n_104),
.B(n_108),
.Y(n_166)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_26),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_105),
.B(n_107),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_46),
.B(n_4),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_106),
.B(n_109),
.Y(n_173)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_21),
.Y(n_107)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_18),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_21),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_26),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_9),
.Y(n_151)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_23),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_112),
.B(n_87),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_84),
.A2(n_36),
.B1(n_35),
.B2(n_30),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_116),
.A2(n_123),
.B1(n_124),
.B2(n_129),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_30),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_117),
.B(n_136),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_56),
.A2(n_36),
.B1(n_35),
.B2(n_50),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_56),
.A2(n_51),
.B1(n_50),
.B2(n_29),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_96),
.A2(n_51),
.B1(n_29),
.B2(n_23),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_126),
.A2(n_134),
.B1(n_138),
.B2(n_139),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_58),
.A2(n_17),
.B1(n_45),
.B2(n_42),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_17),
.B1(n_45),
.B2(n_42),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_131),
.A2(n_135),
.B1(n_176),
.B2(n_159),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_58),
.A2(n_54),
.B1(n_38),
.B2(n_33),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_133),
.A2(n_145),
.B1(n_150),
.B2(n_160),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_54),
.B1(n_38),
.B2(n_33),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_74),
.A2(n_25),
.B1(n_48),
.B2(n_6),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_70),
.B(n_25),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_75),
.B(n_4),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_137),
.B(n_141),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_102),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_57),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_140),
.B(n_144),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_85),
.B(n_8),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_60),
.A2(n_9),
.B1(n_11),
.B2(n_90),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g214 ( 
.A1(n_143),
.A2(n_174),
.B1(n_171),
.B2(n_147),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_69),
.A2(n_79),
.B1(n_103),
.B2(n_104),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_64),
.A2(n_9),
.B1(n_11),
.B2(n_77),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_148),
.A2(n_142),
.B1(n_149),
.B2(n_178),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_69),
.A2(n_9),
.B1(n_79),
.B2(n_97),
.Y(n_150)
);

INVxp33_ASAP7_75t_L g232 ( 
.A(n_151),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_92),
.B(n_94),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_157),
.B(n_164),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_61),
.A2(n_76),
.B1(n_109),
.B2(n_65),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_127),
.C(n_143),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_89),
.A2(n_93),
.B1(n_108),
.B2(n_101),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_66),
.B(n_71),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_152),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_111),
.A2(n_82),
.B1(n_105),
.B2(n_98),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_148),
.A2(n_179),
.B1(n_134),
.B2(n_143),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_180),
.A2(n_193),
.B1(n_198),
.B2(n_219),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_113),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_181),
.B(n_184),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_176),
.A2(n_87),
.B1(n_89),
.B2(n_151),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_183),
.A2(n_226),
.B1(n_235),
.B2(n_233),
.Y(n_274)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_132),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_186),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_128),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_L g271 ( 
.A1(n_187),
.A2(n_190),
.B(n_196),
.Y(n_271)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_188),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_130),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_179),
.Y(n_191)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_191),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_136),
.B(n_137),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_192),
.B(n_202),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_179),
.A2(n_143),
.B1(n_162),
.B2(n_114),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_194),
.B(n_210),
.Y(n_244)
);

OAI32xp33_ASAP7_75t_L g195 ( 
.A1(n_117),
.A2(n_140),
.A3(n_168),
.B1(n_141),
.B2(n_172),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_195),
.B(n_199),
.Y(n_265)
);

NOR4xp25_ASAP7_75t_SL g196 ( 
.A(n_173),
.B(n_125),
.C(n_154),
.D(n_127),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_132),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_197),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_162),
.A2(n_114),
.B1(n_122),
.B2(n_119),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_155),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_164),
.A2(n_139),
.B1(n_114),
.B2(n_157),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_201),
.A2(n_232),
.B(n_182),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_115),
.B(n_121),
.Y(n_202)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_115),
.Y(n_204)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_204),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_156),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_205),
.B(n_209),
.Y(n_269)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_147),
.Y(n_206)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_206),
.Y(n_260)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_119),
.Y(n_207)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_207),
.Y(n_261)
);

INVx3_ASAP7_75t_SL g208 ( 
.A(n_154),
.Y(n_208)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_208),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_158),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_122),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_121),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_211),
.Y(n_272)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_120),
.Y(n_212)
);

BUFx24_ASAP7_75t_L g257 ( 
.A(n_212),
.Y(n_257)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_163),
.Y(n_213)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

OA22x2_ASAP7_75t_L g246 ( 
.A1(n_214),
.A2(n_219),
.B1(n_215),
.B2(n_191),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_170),
.B(n_167),
.C(n_166),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_216),
.B(n_230),
.C(n_208),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_170),
.B(n_120),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_217),
.B(n_218),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_146),
.B(n_171),
.Y(n_218)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_163),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_220),
.B(n_222),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_161),
.B(n_118),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_233),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_146),
.B(n_153),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_118),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_223),
.B(n_225),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_165),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_224),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_144),
.B(n_153),
.Y(n_225)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_177),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_227),
.Y(n_251)
);

NAND3xp33_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_234),
.C(n_237),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_165),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_231),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_174),
.B(n_161),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_169),
.B(n_178),
.Y(n_231)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_142),
.Y(n_233)
);

INVx13_ASAP7_75t_L g234 ( 
.A(n_166),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_149),
.A2(n_176),
.B1(n_151),
.B2(n_143),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_169),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_236),
.A2(n_227),
.B1(n_213),
.B2(n_220),
.Y(n_278)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_169),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_201),
.B1(n_194),
.B2(n_192),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_241),
.A2(n_254),
.B1(n_276),
.B2(n_280),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_246),
.B(n_258),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_185),
.A2(n_182),
.B1(n_189),
.B2(n_203),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_195),
.B(n_200),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_255),
.B(n_266),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_263),
.B(n_274),
.Y(n_306)
);

A2O1A1Ixp33_ASAP7_75t_SL g264 ( 
.A1(n_234),
.A2(n_214),
.B(n_216),
.C(n_237),
.Y(n_264)
);

OA22x2_ASAP7_75t_L g307 ( 
.A1(n_264),
.A2(n_275),
.B1(n_279),
.B2(n_270),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_232),
.B(n_205),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_185),
.A2(n_214),
.B(n_221),
.C(n_202),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_273),
.Y(n_285)
);

NAND3xp33_ASAP7_75t_L g268 ( 
.A(n_187),
.B(n_190),
.C(n_211),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_266),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_214),
.A2(n_230),
.B(n_236),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_270),
.A2(n_264),
.B(n_240),
.Y(n_304)
);

A2O1A1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_230),
.A2(n_223),
.B(n_212),
.C(n_236),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_204),
.A2(n_210),
.B1(n_207),
.B2(n_197),
.Y(n_275)
);

OAI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_186),
.A2(n_206),
.B1(n_224),
.B2(n_229),
.Y(n_276)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_188),
.A2(n_235),
.B1(n_194),
.B2(n_226),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_180),
.A2(n_193),
.B1(n_215),
.B2(n_201),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_247),
.C(n_263),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_282),
.B(n_299),
.C(n_311),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_257),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_283),
.B(n_284),
.Y(n_318)
);

BUFx24_ASAP7_75t_SL g284 ( 
.A(n_269),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_247),
.B(n_241),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_296),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_258),
.A2(n_249),
.B(n_254),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_287),
.A2(n_291),
.B(n_300),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_289),
.B(n_310),
.Y(n_336)
);

NOR2x1_ASAP7_75t_L g291 ( 
.A(n_255),
.B(n_274),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_238),
.B(n_243),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_292),
.B(n_298),
.Y(n_319)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_262),
.Y(n_295)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_295),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_265),
.B(n_250),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_239),
.A2(n_280),
.B1(n_246),
.B2(n_244),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_297),
.A2(n_309),
.B1(n_313),
.B2(n_257),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_256),
.B(n_245),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_244),
.B(n_245),
.C(n_264),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_264),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_262),
.Y(n_301)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_301),
.Y(n_325)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_250),
.Y(n_302)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_302),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_267),
.B(n_248),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_303),
.B(n_307),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_304),
.A2(n_291),
.B(n_307),
.Y(n_341)
);

BUFx5_ASAP7_75t_L g305 ( 
.A(n_242),
.Y(n_305)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_305),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_273),
.B(n_246),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_308),
.B(n_312),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_239),
.A2(n_246),
.B1(n_264),
.B2(n_271),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_240),
.B(n_277),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_272),
.B(n_252),
.C(n_261),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_251),
.B(n_252),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_272),
.A2(n_260),
.B1(n_261),
.B2(n_251),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_275),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_314),
.A2(n_315),
.B1(n_253),
.B2(n_257),
.Y(n_320)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_260),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_282),
.B(n_257),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_316),
.B(n_338),
.C(n_307),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_317),
.A2(n_329),
.B1(n_334),
.B2(n_324),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_320),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_300),
.A2(n_281),
.B(n_259),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_321),
.B(n_322),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_306),
.A2(n_242),
.B1(n_259),
.B2(n_253),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_322),
.A2(n_333),
.B1(n_328),
.B2(n_335),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_290),
.A2(n_253),
.B1(n_259),
.B2(n_308),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_328),
.A2(n_332),
.B(n_288),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_297),
.A2(n_300),
.B1(n_288),
.B2(n_309),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_290),
.A2(n_306),
.B1(n_299),
.B2(n_294),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_306),
.A2(n_290),
.B1(n_302),
.B2(n_286),
.Y(n_333)
);

AOI211xp5_ASAP7_75t_SL g334 ( 
.A1(n_304),
.A2(n_307),
.B(n_285),
.C(n_296),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_313),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_335),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_292),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_337),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_287),
.B(n_303),
.C(n_285),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_291),
.B(n_307),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_342),
.A2(n_346),
.B(n_353),
.Y(n_371)
);

BUFx12_ASAP7_75t_L g343 ( 
.A(n_327),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_343),
.Y(n_370)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_323),
.Y(n_344)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_344),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_345),
.A2(n_329),
.B1(n_317),
.B2(n_339),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_348),
.B(n_350),
.C(n_352),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_336),
.B(n_294),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_349),
.A2(n_351),
.B1(n_356),
.B2(n_357),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_330),
.B(n_311),
.C(n_298),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_331),
.B(n_283),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_315),
.C(n_295),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_341),
.A2(n_314),
.B(n_301),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_321),
.A2(n_293),
.B(n_305),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_354),
.A2(n_320),
.B1(n_332),
.B2(n_333),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_331),
.B(n_293),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_323),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_358),
.A2(n_360),
.B1(n_362),
.B2(n_325),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_324),
.A2(n_339),
.B(n_340),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_359),
.B(n_316),
.C(n_336),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_326),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_363),
.A2(n_362),
.B1(n_357),
.B2(n_353),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_348),
.B(n_330),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_364),
.B(n_369),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_365),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_355),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_367),
.B(n_351),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_345),
.A2(n_326),
.B1(n_334),
.B2(n_338),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_368),
.A2(n_375),
.B1(n_378),
.B2(n_357),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_348),
.B(n_319),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_374),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_350),
.B(n_319),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_347),
.A2(n_337),
.B1(n_325),
.B2(n_327),
.Y(n_375)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_377),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_347),
.A2(n_318),
.B1(n_353),
.B2(n_342),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_350),
.B(n_318),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_379),
.B(n_359),
.Y(n_387)
);

NOR3xp33_ASAP7_75t_SL g381 ( 
.A(n_373),
.B(n_349),
.C(n_355),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_381),
.A2(n_385),
.B1(n_386),
.B2(n_389),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_379),
.B(n_352),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_368),
.B(n_352),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_387),
.B(n_369),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_388),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_376),
.A2(n_361),
.B1(n_342),
.B2(n_359),
.Y(n_389)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_390),
.Y(n_399)
);

CKINVDCx14_ASAP7_75t_R g391 ( 
.A(n_367),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_391),
.A2(n_383),
.B1(n_370),
.B2(n_365),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_392),
.A2(n_371),
.B(n_357),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_384),
.B(n_366),
.C(n_364),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_393),
.B(n_395),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_394),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_384),
.B(n_366),
.C(n_372),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_396),
.A2(n_380),
.B1(n_392),
.B2(n_383),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_401),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_374),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_400),
.B(n_382),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_387),
.B(n_378),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_402),
.B(n_360),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_403),
.B(n_360),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_399),
.A2(n_389),
.B(n_380),
.Y(n_404)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_404),
.Y(n_414)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_399),
.Y(n_407)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_407),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_408),
.B(n_397),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_409),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_405),
.B(n_381),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_411),
.B(n_412),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_415),
.B(n_351),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_414),
.B(n_410),
.C(n_393),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_418),
.B(n_419),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_413),
.B(n_410),
.C(n_395),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_420),
.B(n_417),
.C(n_356),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_416),
.Y(n_421)
);

AOI322xp5_ASAP7_75t_L g422 ( 
.A1(n_421),
.A2(n_370),
.A3(n_343),
.B1(n_413),
.B2(n_406),
.C1(n_373),
.C2(n_358),
.Y(n_422)
);

AOI322xp5_ASAP7_75t_L g425 ( 
.A1(n_422),
.A2(n_343),
.A3(n_406),
.B1(n_344),
.B2(n_398),
.C1(n_375),
.C2(n_346),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_424),
.B(n_409),
.C(n_398),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_425),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_427),
.B(n_423),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_428),
.B(n_426),
.Y(n_429)
);


endmodule