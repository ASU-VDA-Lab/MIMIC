module fake_jpeg_13934_n_527 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_527);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_527;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_442;
wire n_299;
wire n_300;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_18),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

AOI21xp33_ASAP7_75t_L g59 ( 
.A1(n_22),
.A2(n_50),
.B(n_57),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_59),
.B(n_84),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_22),
.B(n_17),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_64),
.B(n_73),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_65),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_23),
.B(n_16),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_67),
.B(n_74),
.Y(n_160)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_68),
.Y(n_183)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

BUFx4f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_72),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_23),
.B(n_15),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_15),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_14),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_75),
.B(n_80),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_76),
.Y(n_176)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_78),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_47),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_79),
.B(n_111),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_50),
.B(n_14),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_81),
.Y(n_155)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_83),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_13),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_85),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_53),
.B(n_0),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_86),
.B(n_92),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_87),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_89),
.Y(n_190)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_91),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_12),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_21),
.B(n_1),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_94),
.B(n_95),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_21),
.B(n_25),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_25),
.B(n_1),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_96),
.B(n_121),
.Y(n_194)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_97),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_98),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_99),
.Y(n_188)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_100),
.Y(n_153)
);

CKINVDCx9p33_ASAP7_75t_R g101 ( 
.A(n_32),
.Y(n_101)
);

CKINVDCx6p67_ASAP7_75t_R g157 ( 
.A(n_101),
.Y(n_157)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_102),
.Y(n_182)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_103),
.Y(n_166)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

INVx13_ASAP7_75t_L g204 ( 
.A(n_104),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_28),
.Y(n_105)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_29),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_110),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_28),
.Y(n_108)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_109),
.Y(n_193)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_35),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_20),
.B(n_1),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_112),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

NAND2xp33_ASAP7_75t_SL g137 ( 
.A(n_113),
.B(n_117),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_20),
.B(n_2),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_120),
.Y(n_158)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_115),
.Y(n_177)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_35),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_118),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

INVx6_ASAP7_75t_SL g142 ( 
.A(n_119),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_33),
.B(n_2),
.Y(n_120)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_35),
.Y(n_121)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_39),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_123),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_33),
.B(n_3),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_49),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_41),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_83),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_125),
.B(n_152),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_89),
.A2(n_39),
.B1(n_58),
.B2(n_56),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_128),
.A2(n_164),
.B1(n_168),
.B2(n_175),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_54),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_132),
.B(n_154),
.Y(n_216)
);

OA21x2_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_100),
.B(n_91),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_134),
.A2(n_138),
.B1(n_140),
.B2(n_173),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_121),
.A2(n_39),
.B1(n_41),
.B2(n_45),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_122),
.A2(n_41),
.B1(n_56),
.B2(n_36),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_71),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_97),
.B(n_54),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_162),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_82),
.A2(n_42),
.B1(n_24),
.B2(n_46),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_65),
.B(n_45),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_165),
.B(n_174),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_104),
.A2(n_40),
.B(n_19),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_167),
.B(n_197),
.C(n_185),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_85),
.A2(n_118),
.B1(n_42),
.B2(n_40),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_98),
.A2(n_51),
.B1(n_44),
.B2(n_36),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_65),
.B(n_51),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_102),
.A2(n_19),
.B1(n_46),
.B2(n_24),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_78),
.B(n_44),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_179),
.B(n_186),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_107),
.A2(n_30),
.B1(n_52),
.B2(n_27),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_185),
.A2(n_197),
.B1(n_149),
.B2(n_143),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_78),
.B(n_30),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_124),
.B(n_30),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_189),
.B(n_191),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_124),
.B(n_4),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_115),
.A2(n_52),
.B1(n_27),
.B2(n_47),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_195),
.A2(n_201),
.B1(n_113),
.B2(n_11),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_63),
.B(n_5),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_196),
.B(n_198),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_109),
.A2(n_52),
.B1(n_27),
.B2(n_47),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_88),
.B(n_6),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_105),
.B(n_6),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_205),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_119),
.A2(n_47),
.B1(n_8),
.B2(n_10),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_117),
.A2(n_47),
.B1(n_8),
.B2(n_11),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_202),
.A2(n_157),
.B1(n_166),
.B2(n_192),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_108),
.B(n_7),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_133),
.A2(n_93),
.B1(n_66),
.B2(n_87),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_206),
.A2(n_214),
.B(n_252),
.Y(n_313)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_139),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_207),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_208),
.Y(n_282)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_7),
.B(n_8),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_209),
.B(n_264),
.Y(n_279)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_129),
.Y(n_211)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_211),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_132),
.B(n_60),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_212),
.B(n_233),
.C(n_234),
.Y(n_301)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_129),
.Y(n_213)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_213),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_167),
.A2(n_72),
.B(n_76),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_215),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_154),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_217),
.B(n_222),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_204),
.Y(n_218)
);

BUFx24_ASAP7_75t_L g284 ( 
.A(n_218),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_153),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_220),
.Y(n_289)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_130),
.Y(n_221)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_221),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_142),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_130),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_223),
.Y(n_300)
);

AO22x1_ASAP7_75t_L g224 ( 
.A1(n_137),
.A2(n_7),
.B1(n_12),
.B2(n_142),
.Y(n_224)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_224),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_131),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_226),
.B(n_229),
.Y(n_286)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_146),
.Y(n_227)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_227),
.Y(n_302)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_228),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_131),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_131),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_230),
.B(n_259),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_178),
.A2(n_159),
.B1(n_170),
.B2(n_160),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_231),
.A2(n_236),
.B1(n_248),
.B2(n_249),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_126),
.B(n_158),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_232),
.B(n_235),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_144),
.B(n_183),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_144),
.B(n_183),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_146),
.B(n_140),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_137),
.A2(n_202),
.B1(n_138),
.B2(n_134),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_144),
.B(n_145),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_237),
.B(n_238),
.C(n_240),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_136),
.B(n_156),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_163),
.A2(n_199),
.B(n_155),
.C(n_147),
.Y(n_239)
);

A2O1A1Ixp33_ASAP7_75t_L g293 ( 
.A1(n_239),
.A2(n_232),
.B(n_273),
.C(n_219),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_134),
.B(n_181),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_135),
.Y(n_241)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_241),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_171),
.B(n_150),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_243),
.B(n_246),
.Y(n_287)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_184),
.Y(n_244)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_244),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_135),
.B(n_169),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_245),
.B(n_253),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_171),
.B(n_150),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_141),
.Y(n_247)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_247),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_127),
.A2(n_193),
.B1(n_192),
.B2(n_190),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_169),
.Y(n_250)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_250),
.Y(n_311)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_184),
.Y(n_251)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_251),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_181),
.B(n_153),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_L g254 ( 
.A1(n_127),
.A2(n_193),
.B1(n_177),
.B2(n_203),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_254),
.A2(n_255),
.B1(n_270),
.B2(n_272),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_157),
.A2(n_177),
.B1(n_203),
.B2(n_143),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_180),
.Y(n_256)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_256),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_180),
.B(n_151),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_257),
.B(n_267),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_151),
.B(n_149),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_258),
.B(n_233),
.C(n_234),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_157),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_157),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_261),
.B(n_263),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_141),
.Y(n_263)
);

BUFx5_ASAP7_75t_L g266 ( 
.A(n_148),
.Y(n_266)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_266),
.Y(n_324)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_182),
.Y(n_267)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_148),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_269),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_176),
.A2(n_187),
.B1(n_182),
.B2(n_172),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_176),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_271),
.B(n_259),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_187),
.A2(n_172),
.B1(n_161),
.B2(n_139),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_260),
.A2(n_139),
.B1(n_161),
.B2(n_188),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_278),
.A2(n_280),
.B1(n_285),
.B2(n_249),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_260),
.A2(n_161),
.B1(n_188),
.B2(n_216),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_216),
.A2(n_188),
.B1(n_252),
.B2(n_235),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_206),
.A2(n_264),
.B1(n_240),
.B2(n_273),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_288),
.A2(n_222),
.B1(n_258),
.B2(n_267),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_218),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_290),
.B(n_298),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_293),
.B(n_305),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_253),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_245),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_303),
.B(n_227),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_265),
.B(n_237),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_306),
.B(n_309),
.C(n_211),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_237),
.B(n_212),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_212),
.B(n_268),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_312),
.B(n_323),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_242),
.B(n_262),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_316),
.B(n_319),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_239),
.B(n_225),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_320),
.Y(n_338)
);

AOI22x1_ASAP7_75t_L g321 ( 
.A1(n_210),
.A2(n_248),
.B1(n_214),
.B2(n_224),
.Y(n_321)
);

OA22x2_ASAP7_75t_L g349 ( 
.A1(n_321),
.A2(n_221),
.B1(n_223),
.B2(n_207),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_238),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_233),
.B(n_234),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_257),
.B(n_238),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_325),
.B(n_277),
.Y(n_355)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_275),
.Y(n_327)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_327),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_317),
.A2(n_224),
.B1(n_272),
.B2(n_263),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_328),
.A2(n_341),
.B1(n_342),
.B2(n_358),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_329),
.B(n_354),
.C(n_297),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_330),
.A2(n_331),
.B(n_352),
.Y(n_388)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_275),
.Y(n_332)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_332),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_334),
.B(n_346),
.Y(n_373)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_291),
.Y(n_335)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_335),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_336),
.B(n_309),
.Y(n_368)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_291),
.Y(n_337)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_337),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_280),
.A2(n_254),
.B1(n_271),
.B2(n_213),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_339),
.A2(n_356),
.B1(n_307),
.B2(n_310),
.Y(n_371)
);

BUFx12f_ASAP7_75t_L g340 ( 
.A(n_284),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_340),
.B(n_345),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_317),
.A2(n_208),
.B1(n_269),
.B2(n_250),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_313),
.A2(n_241),
.B1(n_247),
.B2(n_244),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_302),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_343),
.Y(n_375)
);

INVx6_ASAP7_75t_L g345 ( 
.A(n_282),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_302),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_287),
.B(n_251),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_347),
.Y(n_380)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_304),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_348),
.B(n_351),
.Y(n_374)
);

AND2x2_ASAP7_75t_SL g377 ( 
.A(n_349),
.B(n_364),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_279),
.A2(n_258),
.B(n_256),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_350),
.A2(n_360),
.B(n_361),
.Y(n_366)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_282),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_313),
.A2(n_228),
.B(n_266),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_283),
.B(n_312),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_353),
.B(n_365),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_277),
.B(n_306),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_355),
.B(n_357),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_285),
.A2(n_281),
.B1(n_278),
.B2(n_279),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_304),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_281),
.A2(n_321),
.B1(n_294),
.B2(n_296),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_284),
.B(n_286),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_359),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_294),
.A2(n_296),
.B(n_279),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_305),
.A2(n_321),
.B1(n_301),
.B2(n_322),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_292),
.B(n_297),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_362),
.B(n_289),
.Y(n_387)
);

MAJx2_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_274),
.C(n_318),
.Y(n_379)
);

FAx1_ASAP7_75t_L g364 ( 
.A(n_301),
.B(n_284),
.CI(n_293),
.CON(n_364),
.SN(n_364)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_325),
.B(n_323),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_368),
.B(n_370),
.C(n_378),
.Y(n_420)
);

OA21x2_ASAP7_75t_L g369 ( 
.A1(n_358),
.A2(n_284),
.B(n_274),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_369),
.B(n_391),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_371),
.A2(n_384),
.B1(n_396),
.B2(n_365),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_354),
.B(n_310),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_379),
.B(n_366),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_328),
.A2(n_324),
.B1(n_314),
.B2(n_276),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_383),
.A2(n_352),
.B(n_342),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_356),
.A2(n_314),
.B1(n_318),
.B2(n_299),
.Y(n_384)
);

AND2x6_ASAP7_75t_L g385 ( 
.A(n_364),
.B(n_308),
.Y(n_385)
);

AOI21xp33_ASAP7_75t_L g424 ( 
.A1(n_385),
.A2(n_395),
.B(n_350),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_387),
.B(n_338),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_341),
.A2(n_315),
.B1(n_299),
.B2(n_324),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_389),
.A2(n_348),
.B1(n_357),
.B2(n_343),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_344),
.B(n_295),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_344),
.B(n_295),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_392),
.B(n_337),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_333),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_393),
.B(n_380),
.Y(n_410)
);

AND2x6_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_308),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_330),
.A2(n_361),
.B1(n_331),
.B2(n_360),
.Y(n_396)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_394),
.Y(n_398)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_398),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_399),
.B(n_421),
.Y(n_425)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_394),
.Y(n_400)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_400),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_374),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_401),
.B(n_407),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_402),
.A2(n_424),
.B(n_375),
.Y(n_445)
);

XOR2x2_ASAP7_75t_L g442 ( 
.A(n_403),
.B(n_378),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_367),
.A2(n_339),
.B1(n_363),
.B2(n_349),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_404),
.A2(n_405),
.B1(n_369),
.B2(n_384),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_368),
.B(n_336),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_406),
.B(n_370),
.C(n_366),
.Y(n_428)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_372),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_409),
.A2(n_423),
.B1(n_367),
.B2(n_383),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_410),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_374),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_411),
.B(n_412),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_390),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_413),
.B(n_414),
.Y(n_430)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_372),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_381),
.B(n_338),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_415),
.B(n_416),
.Y(n_439)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_376),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_377),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_417),
.B(n_419),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_377),
.A2(n_353),
.B1(n_349),
.B2(n_329),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_418),
.A2(n_388),
.B(n_377),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_373),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_391),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_393),
.B(n_326),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_422),
.B(n_387),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_369),
.A2(n_349),
.B1(n_329),
.B2(n_335),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_426),
.A2(n_431),
.B1(n_434),
.B2(n_446),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_427),
.A2(n_445),
.B1(n_402),
.B2(n_433),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_428),
.B(n_415),
.C(n_404),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_429),
.B(n_433),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_409),
.A2(n_397),
.B1(n_379),
.B2(n_396),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_417),
.A2(n_388),
.B(n_395),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_423),
.A2(n_392),
.B1(n_381),
.B2(n_397),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_437),
.B(n_444),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_418),
.A2(n_385),
.B(n_386),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_440),
.B(n_443),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_448),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_408),
.A2(n_386),
.B(n_380),
.Y(n_443)
);

OA21x2_ASAP7_75t_L g444 ( 
.A1(n_408),
.A2(n_389),
.B(n_375),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_421),
.A2(n_382),
.B1(n_376),
.B2(n_346),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_406),
.B(n_382),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_448),
.B(n_420),
.Y(n_452)
);

MAJx2_ASAP7_75t_L g450 ( 
.A(n_428),
.B(n_403),
.C(n_420),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_450),
.B(n_457),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_452),
.B(n_456),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_453),
.A2(n_426),
.B(n_440),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_419),
.Y(n_455)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_455),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_442),
.B(n_413),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_458),
.B(n_462),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_412),
.C(n_411),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_459),
.B(n_460),
.C(n_463),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_431),
.B(n_401),
.C(n_398),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_438),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_461),
.B(n_464),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_443),
.B(n_405),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_441),
.B(n_416),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_437),
.B(n_340),
.Y(n_464)
);

XNOR2x1_ASAP7_75t_L g465 ( 
.A(n_434),
.B(n_340),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_465),
.B(n_466),
.C(n_467),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_445),
.B(n_400),
.C(n_407),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_441),
.B(n_414),
.C(n_332),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_469),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_454),
.A2(n_429),
.B(n_439),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_473),
.B(n_478),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_449),
.A2(n_447),
.B(n_425),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_474),
.B(n_483),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_467),
.B(n_438),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_475),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_457),
.B(n_447),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_459),
.B(n_425),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_479),
.B(n_482),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_460),
.B(n_340),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_452),
.B(n_439),
.C(n_430),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_471),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_484),
.B(n_495),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_470),
.B(n_466),
.C(n_450),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_485),
.B(n_488),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_472),
.A2(n_451),
.B(n_444),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_472),
.B(n_465),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_490),
.B(n_491),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_470),
.B(n_456),
.C(n_462),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_480),
.B(n_458),
.C(n_468),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_494),
.B(n_481),
.C(n_480),
.Y(n_500)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_477),
.Y(n_495)
);

XNOR2x1_ASAP7_75t_L g496 ( 
.A(n_490),
.B(n_481),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_496),
.B(n_502),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_493),
.A2(n_469),
.B1(n_473),
.B2(n_475),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_498),
.B(n_500),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_489),
.A2(n_475),
.B(n_483),
.Y(n_499)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_499),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_485),
.B(n_494),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_501),
.B(n_505),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_493),
.A2(n_427),
.B1(n_444),
.B2(n_446),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_487),
.A2(n_486),
.B1(n_444),
.B2(n_432),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_503),
.A2(n_492),
.B(n_491),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_507),
.B(n_510),
.Y(n_515)
);

CKINVDCx14_ASAP7_75t_R g508 ( 
.A(n_497),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_508),
.B(n_476),
.Y(n_514)
);

AOI322xp5_ASAP7_75t_L g510 ( 
.A1(n_502),
.A2(n_488),
.A3(n_432),
.B1(n_435),
.B2(n_430),
.C1(n_463),
.C2(n_476),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_501),
.B(n_500),
.C(n_504),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_512),
.B(n_496),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_514),
.B(n_518),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_516),
.B(n_517),
.Y(n_520)
);

A2O1A1Ixp33_ASAP7_75t_SL g517 ( 
.A1(n_509),
.A2(n_435),
.B(n_327),
.C(n_345),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_512),
.B(n_351),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_513),
.B(n_276),
.C(n_311),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_519),
.A2(n_511),
.B(n_507),
.Y(n_521)
);

NAND3xp33_ASAP7_75t_L g524 ( 
.A(n_521),
.B(n_506),
.C(n_300),
.Y(n_524)
);

AOI21x1_ASAP7_75t_L g523 ( 
.A1(n_522),
.A2(n_515),
.B(n_517),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_523),
.A2(n_524),
.B1(n_520),
.B2(n_506),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_525),
.A2(n_300),
.B(n_311),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_526),
.B(n_315),
.Y(n_527)
);


endmodule