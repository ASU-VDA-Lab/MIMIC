module fake_jpeg_23327_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_37),
.Y(n_45)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_40),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_22),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_41),
.B(n_30),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_56),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_27),
.B1(n_18),
.B2(n_17),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_38),
.B(n_37),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_27),
.B1(n_18),
.B2(n_20),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_54),
.B1(n_26),
.B2(n_28),
.Y(n_69)
);

CKINVDCx12_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_50),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_33),
.C(n_39),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_58),
.C(n_36),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_27),
.B1(n_22),
.B2(n_29),
.Y(n_54)
);

NAND3xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_0),
.C(n_1),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_0),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_20),
.C(n_29),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_78),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_65),
.Y(n_89)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_67),
.Y(n_90)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_70),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_69),
.A2(n_12),
.B1(n_11),
.B2(n_4),
.Y(n_111)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_71),
.A2(n_73),
.B(n_78),
.Y(n_101)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_76),
.Y(n_104)
);

AND2x4_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

FAx1_ASAP7_75t_SL g75 ( 
.A(n_54),
.B(n_39),
.CI(n_35),
.CON(n_75),
.SN(n_75)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_75),
.B(n_77),
.Y(n_94)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_40),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_38),
.C(n_16),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_80),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_37),
.B1(n_42),
.B2(n_47),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_24),
.B1(n_23),
.B2(n_32),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_82),
.B(n_83),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_19),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_85),
.Y(n_110)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_26),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_44),
.B(n_28),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_24),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

NAND2xp33_ASAP7_75t_SL g93 ( 
.A(n_88),
.B(n_52),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_69),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_42),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_81),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_71),
.B(n_88),
.Y(n_118)
);

OA22x2_ASAP7_75t_SL g97 ( 
.A1(n_73),
.A2(n_42),
.B1(n_32),
.B2(n_31),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_99),
.B1(n_100),
.B2(n_107),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_65),
.A2(n_24),
.B1(n_23),
.B2(n_32),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_80),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_73),
.A2(n_31),
.B1(n_15),
.B2(n_13),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_73),
.A2(n_31),
.B1(n_2),
.B2(n_3),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_109),
.A2(n_111),
.B1(n_12),
.B2(n_4),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_97),
.A2(n_66),
.B1(n_70),
.B2(n_76),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_114),
.Y(n_144)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_124),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_104),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_116),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_101),
.C(n_108),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_118),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_59),
.C(n_62),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_94),
.A2(n_75),
.B(n_82),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_127),
.B(n_130),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_123),
.Y(n_145)
);

AOI32xp33_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_75),
.A3(n_82),
.B1(n_67),
.B2(n_59),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_63),
.Y(n_125)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_126),
.B(n_132),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_1),
.Y(n_127)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_129),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_3),
.Y(n_131)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_95),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_133),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_113),
.Y(n_139)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_141),
.B(n_147),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_105),
.B(n_109),
.C(n_106),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_122),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_122),
.A2(n_102),
.B1(n_100),
.B2(n_106),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_151),
.A2(n_129),
.B1(n_127),
.B2(n_131),
.Y(n_163)
);

AOI221xp5_ASAP7_75t_L g152 ( 
.A1(n_145),
.A2(n_130),
.B1(n_107),
.B2(n_127),
.C(n_117),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_154),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_134),
.B(n_96),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_144),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_161),
.Y(n_176)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_128),
.Y(n_158)
);

AOI21x1_ASAP7_75t_L g169 ( 
.A1(n_158),
.A2(n_147),
.B(n_136),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_119),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_160),
.C(n_141),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_143),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_165),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_164),
.B1(n_151),
.B2(n_137),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_124),
.B1(n_96),
.B2(n_126),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_142),
.A2(n_111),
.B(n_103),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_150),
.B(n_148),
.Y(n_167)
);

OA21x2_ASAP7_75t_L g178 ( 
.A1(n_167),
.A2(n_169),
.B(n_153),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_162),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_172),
.C(n_160),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_143),
.C(n_136),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_174),
.B(n_135),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_178),
.A2(n_186),
.B(n_139),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_179),
.A2(n_185),
.B1(n_175),
.B2(n_169),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_177),
.A2(n_166),
.B(n_161),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_182),
.C(n_172),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_137),
.C(n_103),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_184),
.A2(n_171),
.B1(n_114),
.B2(n_139),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_173),
.B(n_91),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_176),
.B(n_158),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_187),
.B(n_183),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_188),
.A2(n_192),
.B1(n_193),
.B2(n_190),
.Y(n_198)
);

FAx1_ASAP7_75t_SL g190 ( 
.A(n_178),
.B(n_167),
.CI(n_168),
.CON(n_190),
.SN(n_190)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_191),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_158),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_193),
.A2(n_189),
.B(n_190),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_198),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_195),
.B(n_197),
.Y(n_201)
);

AOI322xp5_ASAP7_75t_L g197 ( 
.A1(n_188),
.A2(n_99),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_196),
.A2(n_191),
.B1(n_187),
.B2(n_7),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_199),
.B(n_194),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_202),
.A2(n_203),
.B(n_201),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_200),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_203)
);

NOR3xp33_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_199),
.C(n_5),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_9),
.Y(n_206)
);


endmodule