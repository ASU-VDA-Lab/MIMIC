module fake_netlist_5_1912_n_191 (n_29, n_16, n_43, n_0, n_12, n_9, n_47, n_36, n_25, n_18, n_27, n_42, n_22, n_1, n_8, n_45, n_10, n_24, n_28, n_46, n_21, n_44, n_40, n_34, n_38, n_4, n_32, n_35, n_41, n_51, n_11, n_17, n_19, n_7, n_37, n_15, n_26, n_30, n_20, n_5, n_33, n_14, n_48, n_2, n_31, n_23, n_13, n_50, n_3, n_49, n_52, n_6, n_39, n_191);

input n_29;
input n_16;
input n_43;
input n_0;
input n_12;
input n_9;
input n_47;
input n_36;
input n_25;
input n_18;
input n_27;
input n_42;
input n_22;
input n_1;
input n_8;
input n_45;
input n_10;
input n_24;
input n_28;
input n_46;
input n_21;
input n_44;
input n_40;
input n_34;
input n_38;
input n_4;
input n_32;
input n_35;
input n_41;
input n_51;
input n_11;
input n_17;
input n_19;
input n_7;
input n_37;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_33;
input n_14;
input n_48;
input n_2;
input n_31;
input n_23;
input n_13;
input n_50;
input n_3;
input n_49;
input n_52;
input n_6;
input n_39;

output n_191;

wire n_137;
wire n_168;
wire n_164;
wire n_91;
wire n_82;
wire n_122;
wire n_142;
wire n_176;
wire n_140;
wire n_124;
wire n_86;
wire n_136;
wire n_146;
wire n_182;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_101;
wire n_75;
wire n_180;
wire n_184;
wire n_65;
wire n_78;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_189;
wire n_165;
wire n_111;
wire n_108;
wire n_129;
wire n_66;
wire n_98;
wire n_177;
wire n_60;
wire n_155;
wire n_152;
wire n_107;
wire n_58;
wire n_69;
wire n_116;
wire n_117;
wire n_94;
wire n_113;
wire n_123;
wire n_139;
wire n_105;
wire n_80;
wire n_179;
wire n_125;
wire n_167;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_156;
wire n_126;
wire n_84;
wire n_130;
wire n_157;
wire n_79;
wire n_131;
wire n_151;
wire n_173;
wire n_53;
wire n_160;
wire n_188;
wire n_190;
wire n_158;
wire n_154;
wire n_100;
wire n_62;
wire n_138;
wire n_148;
wire n_71;
wire n_109;
wire n_112;
wire n_85;
wire n_159;
wire n_163;
wire n_95;
wire n_119;
wire n_183;
wire n_185;
wire n_175;
wire n_169;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_181;
wire n_54;
wire n_147;
wire n_178;
wire n_67;
wire n_121;
wire n_76;
wire n_87;
wire n_150;
wire n_170;
wire n_162;
wire n_64;
wire n_106;
wire n_77;
wire n_102;
wire n_161;
wire n_81;
wire n_118;
wire n_89;
wire n_115;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_174;
wire n_186;
wire n_134;
wire n_187;
wire n_104;
wire n_172;
wire n_103;
wire n_56;
wire n_63;
wire n_97;
wire n_141;
wire n_166;
wire n_171;
wire n_153;
wire n_145;
wire n_88;
wire n_110;

INVx2_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

BUFx2_ASAP7_75t_SL g64 ( 
.A(n_35),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

INVxp67_ASAP7_75t_SL g69 ( 
.A(n_15),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_13),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_38),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_0),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_2),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_88),
.Y(n_98)
);

AND2x6_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_53),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_69),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

AND2x4_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_54),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_64),
.B1(n_73),
.B2(n_76),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_55),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

AND2x4_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_83),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_84),
.B(n_78),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_90),
.Y(n_114)
);

AND2x4_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_78),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_67),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_77),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_99),
.Y(n_126)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_102),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_114),
.A2(n_97),
.B(n_96),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_99),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_72),
.B1(n_75),
.B2(n_74),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_70),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

OAI21x1_ASAP7_75t_L g138 ( 
.A1(n_126),
.A2(n_131),
.B(n_130),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

AND2x4_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_4),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

OAI21x1_ASAP7_75t_L g143 ( 
.A1(n_136),
.A2(n_52),
.B(n_7),
.Y(n_143)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_9),
.B(n_10),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_12),
.Y(n_146)
);

OAI21x1_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_125),
.B(n_134),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_127),
.Y(n_148)
);

OAI221xp5_ASAP7_75t_L g149 ( 
.A1(n_146),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.C(n_24),
.Y(n_149)
);

OAI21x1_ASAP7_75t_L g150 ( 
.A1(n_143),
.A2(n_25),
.B(n_27),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_29),
.Y(n_152)
);

OR2x6_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_30),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_152),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_154),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_157),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_160),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_164),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_158),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_144),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_165),
.Y(n_174)
);

AND2x4_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_162),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_31),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_171),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_168),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_172),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_180),
.Y(n_181)
);

NAND2xp33_ASAP7_75t_SL g182 ( 
.A(n_181),
.B(n_178),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_181),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_175),
.Y(n_184)
);

OA22x2_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_176),
.B1(n_173),
.B2(n_177),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_185),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_186),
.Y(n_187)
);

OR3x1_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_33),
.C(n_34),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_R g189 ( 
.A1(n_188),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_191)
);


endmodule