module fake_jpeg_3423_n_190 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_190);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_26),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx8_ASAP7_75t_SL g59 ( 
.A(n_31),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_5),
.B(n_6),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_67),
.Y(n_74)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx5_ASAP7_75t_SL g72 ( 
.A(n_65),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_61),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_46),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_71),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_55),
.B1(n_45),
.B2(n_54),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_47),
.B1(n_46),
.B2(n_66),
.Y(n_87)
);

AO22x1_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_46),
.B1(n_45),
.B2(n_59),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_68),
.B1(n_63),
.B2(n_66),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_65),
.B(n_51),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_78),
.B(n_60),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_52),
.B1(n_58),
.B2(n_62),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_58),
.C(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_52),
.Y(n_92)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_17),
.B1(n_42),
.B2(n_40),
.Y(n_112)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_53),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_1),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_92),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_93),
.B(n_94),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_72),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_96),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_50),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_62),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_98),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_50),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_44),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_71),
.B1(n_77),
.B2(n_79),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_100),
.A2(n_101),
.B1(n_112),
.B2(n_6),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_90),
.A2(n_77),
.B1(n_73),
.B2(n_3),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_4),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_18),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_110),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_97),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_34),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_2),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_115),
.B(n_116),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_3),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_91),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_9),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_91),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_119),
.B(n_16),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_91),
.C(n_85),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_121),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_100),
.A2(n_88),
.B1(n_21),
.B2(n_22),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_107),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_126),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_4),
.B(n_5),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_128),
.Y(n_153)
);

OA21x2_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_39),
.B(n_38),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_114),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_129),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_37),
.C(n_36),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_132),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_7),
.B(n_8),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_10),
.B(n_11),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_30),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_SL g139 ( 
.A(n_133),
.B(n_101),
.C(n_108),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_142),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_123),
.B(n_111),
.Y(n_142)
);

NOR3xp33_ASAP7_75t_SL g143 ( 
.A(n_126),
.B(n_112),
.C(n_32),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_144),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_126),
.B(n_103),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_146),
.B(n_151),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_150),
.Y(n_162)
);

OAI22x1_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_28),
.B1(n_25),
.B2(n_24),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_128),
.Y(n_161)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_119),
.C(n_122),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_166),
.C(n_167),
.Y(n_172)
);

NOR2xp67_ASAP7_75t_R g159 ( 
.A(n_152),
.B(n_130),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_161),
.Y(n_176)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_163),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_131),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_12),
.C(n_13),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_140),
.A2(n_13),
.B(n_14),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_168),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_157),
.A2(n_145),
.B1(n_164),
.B2(n_165),
.Y(n_169)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_158),
.B(n_151),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_138),
.C(n_14),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_166),
.C(n_162),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_145),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_178),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_176),
.B(n_139),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_170),
.A2(n_143),
.B1(n_138),
.B2(n_16),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_181),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_180),
.A2(n_175),
.B(n_170),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_173),
.B(n_172),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_182),
.C(n_181),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_183),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_171),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_15),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_15),
.Y(n_190)
);


endmodule