module fake_netlist_5_1854_n_1160 (n_91, n_82, n_122, n_10, n_24, n_124, n_86, n_83, n_61, n_90, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_105, n_80, n_4, n_125, n_35, n_73, n_17, n_92, n_19, n_120, n_30, n_5, n_33, n_14, n_84, n_23, n_29, n_79, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_1160);

input n_91;
input n_82;
input n_122;
input n_10;
input n_24;
input n_124;
input n_86;
input n_83;
input n_61;
input n_90;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_30;
input n_5;
input n_33;
input n_14;
input n_84;
input n_23;
input n_29;
input n_79;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1160;

wire n_137;
wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_1141;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_136;
wire n_146;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_127;
wire n_1150;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_1139;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_1055;
wire n_351;
wire n_643;
wire n_620;
wire n_367;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_525;
wire n_493;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_155;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_1157;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_823;
wire n_983;
wire n_725;
wire n_501;
wire n_1128;
wire n_139;
wire n_280;
wire n_744;
wire n_1021;
wire n_629;
wire n_590;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_864;
wire n_443;
wire n_173;
wire n_859;
wire n_1110;
wire n_951;
wire n_1121;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_314;
wire n_247;
wire n_433;
wire n_368;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_946;
wire n_1048;
wire n_417;
wire n_612;
wire n_1001;
wire n_212;
wire n_385;
wire n_516;
wire n_933;
wire n_498;
wire n_788;
wire n_507;
wire n_1152;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_133;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_147;
wire n_936;
wire n_757;
wire n_1090;
wire n_307;
wire n_633;
wire n_530;
wire n_439;
wire n_150;
wire n_1024;
wire n_1063;
wire n_556;
wire n_1107;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1143;
wire n_804;
wire n_867;
wire n_186;
wire n_1124;
wire n_537;
wire n_1158;
wire n_134;
wire n_902;
wire n_191;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_171;
wire n_153;
wire n_756;
wire n_1145;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_1049;
wire n_1153;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_1154;
wire n_286;
wire n_883;
wire n_1135;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_519;
wire n_406;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_1108;
wire n_325;
wire n_449;
wire n_1100;
wire n_132;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_1147;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_167;
wire n_607;
wire n_976;
wire n_1096;
wire n_234;
wire n_343;
wire n_1095;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_156;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_157;
wire n_814;
wire n_131;
wire n_192;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_1142;
wire n_660;
wire n_223;
wire n_1114;
wire n_1129;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_138;
wire n_1148;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_163;
wire n_339;
wire n_1146;
wire n_1149;
wire n_882;
wire n_185;
wire n_243;
wire n_183;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_169;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_1073;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_181;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_141;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_922;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_145;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_837;
wire n_673;
wire n_528;
wire n_479;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_974;
wire n_432;
wire n_395;
wire n_164;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_1159;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_142;
wire n_743;
wire n_214;
wire n_328;
wire n_140;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_829;
wire n_749;
wire n_928;
wire n_144;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_1151;
wire n_1134;
wire n_881;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_129;
wire n_342;
wire n_517;
wire n_482;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_1069;
wire n_236;
wire n_1075;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_338;
wire n_149;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_130;
wire n_322;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_1122;
wire n_151;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_770;
wire n_288;
wire n_188;
wire n_190;
wire n_844;
wire n_201;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_1041;
wire n_989;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1015;
wire n_1000;
wire n_891;
wire n_1140;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_846;
wire n_586;
wire n_1058;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_170;
wire n_332;
wire n_1053;
wire n_1101;
wire n_161;
wire n_273;
wire n_585;
wire n_349;
wire n_1106;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_917;
wire n_1014;
wire n_279;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_174;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1116;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_993;
wire n_440;
wire n_425;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1131;
wire n_1059;
wire n_1084;
wire n_176;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_182;
wire n_143;
wire n_1005;
wire n_354;
wire n_575;
wire n_647;
wire n_480;
wire n_679;
wire n_237;
wire n_513;
wire n_710;
wire n_407;
wire n_527;
wire n_707;
wire n_795;
wire n_832;
wire n_857;
wire n_695;
wire n_1072;
wire n_180;
wire n_1094;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_1027;
wire n_805;
wire n_490;
wire n_1156;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_1136;
wire n_815;
wire n_246;
wire n_596;
wire n_179;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_128;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_135;
wire n_1109;
wire n_657;
wire n_126;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_202;
wire n_1080;
wire n_266;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_154;
wire n_148;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_159;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_1138;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_200;
wire n_1032;
wire n_1056;
wire n_162;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_1155;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_1123;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_187;
wire n_401;
wire n_348;
wire n_1029;
wire n_166;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_1144;
wire n_1137;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

INVx1_ASAP7_75t_L g126 ( 
.A(n_30),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_120),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_49),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

BUFx2_ASAP7_75t_SL g133 ( 
.A(n_104),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_100),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_113),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_80),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_24),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_5),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_122),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_24),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_66),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_101),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_4),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_7),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_53),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_41),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_14),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_111),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_4),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_14),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_102),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_116),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_38),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_51),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_64),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_32),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_123),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_78),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_37),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_117),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_88),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_1),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_94),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_125),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g171 ( 
.A(n_29),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_86),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_106),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_43),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_11),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_114),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_52),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_74),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_6),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_46),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_118),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_139),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_141),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_148),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_138),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_134),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_135),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_140),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_130),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_149),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_142),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_145),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_127),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_127),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_151),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_153),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_158),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_161),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_165),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_166),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_167),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_152),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_170),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_156),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_154),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_172),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_203),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_189),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_191),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_192),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_184),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_184),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_195),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_185),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_186),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_211),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_193),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_196),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_198),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_200),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_201),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_202),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_204),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_205),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_206),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_210),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_207),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_208),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_189),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_203),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_187),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_184),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_198),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_187),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_187),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_193),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_194),
.B(n_168),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_187),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_187),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_203),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_203),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_187),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_222),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_215),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_226),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_223),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_224),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_227),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_260),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_214),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_225),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_215),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_244),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_218),
.Y(n_278)
);

INVxp67_ASAP7_75t_SL g279 ( 
.A(n_253),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

INVxp67_ASAP7_75t_SL g281 ( 
.A(n_253),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_214),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_228),
.Y(n_283)
);

INVxp33_ASAP7_75t_L g284 ( 
.A(n_242),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_264),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_221),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_238),
.Y(n_287)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_253),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_217),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_231),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_219),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_220),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_244),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_254),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_265),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_229),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_262),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_257),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_261),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_238),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_258),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_253),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_250),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_230),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_256),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_232),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_240),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_233),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_234),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_236),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_239),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_237),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_237),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_240),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_278),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_292),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_287),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_272),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_307),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_300),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_268),
.Y(n_321)
);

INVxp33_ASAP7_75t_SL g322 ( 
.A(n_283),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_273),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_314),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_292),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_290),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_314),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_271),
.B(n_216),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_276),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_312),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_276),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_293),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_294),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_293),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_312),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_294),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_305),
.Y(n_337)
);

NAND2xp33_ASAP7_75t_R g338 ( 
.A(n_304),
.B(n_216),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_273),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_295),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_295),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_297),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_267),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_297),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_298),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_313),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_282),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_267),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_310),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_313),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_298),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_282),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_299),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_284),
.B(n_235),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_289),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_303),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_304),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_275),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_303),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_301),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_316),
.B(n_306),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_343),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_358),
.Y(n_363)
);

BUFx12f_ASAP7_75t_L g364 ( 
.A(n_315),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_331),
.A2(n_249),
.B1(n_251),
.B2(n_246),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_358),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_323),
.Y(n_367)
);

NOR2x1_ASAP7_75t_L g368 ( 
.A(n_328),
.B(n_248),
.Y(n_368)
);

OAI22x1_ASAP7_75t_L g369 ( 
.A1(n_346),
.A2(n_296),
.B1(n_308),
.B2(n_306),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_323),
.B(n_289),
.Y(n_370)
);

OAI21x1_ASAP7_75t_L g371 ( 
.A1(n_348),
.A2(n_302),
.B(n_269),
.Y(n_371)
);

BUFx8_ASAP7_75t_L g372 ( 
.A(n_354),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_325),
.Y(n_373)
);

AND2x4_ASAP7_75t_L g374 ( 
.A(n_339),
.B(n_291),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_355),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_333),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_360),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_336),
.B(n_308),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_355),
.B(n_291),
.Y(n_379)
);

CKINVDCx6p67_ASAP7_75t_R g380 ( 
.A(n_319),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_326),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_340),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_341),
.B(n_309),
.Y(n_383)
);

OAI21x1_ASAP7_75t_L g384 ( 
.A1(n_342),
.A2(n_302),
.B(n_269),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_344),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_355),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_345),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_351),
.Y(n_388)
);

INVx5_ASAP7_75t_L g389 ( 
.A(n_355),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_347),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_353),
.B(n_309),
.Y(n_391)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_356),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_357),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_359),
.A2(n_296),
.B1(n_311),
.B2(n_301),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_349),
.B(n_311),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_321),
.B(n_330),
.Y(n_396)
);

NAND2xp33_ASAP7_75t_L g397 ( 
.A(n_350),
.B(n_156),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_335),
.B(n_286),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_352),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_319),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_352),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_318),
.Y(n_402)
);

INVx2_ASAP7_75t_SL g403 ( 
.A(n_320),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_337),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_329),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_327),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_332),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_334),
.Y(n_408)
);

INVx6_ASAP7_75t_L g409 ( 
.A(n_324),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_331),
.Y(n_410)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_322),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_317),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_338),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_338),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_356),
.B(n_241),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_357),
.B(n_255),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_323),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_358),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_316),
.B(n_286),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_358),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_357),
.B(n_243),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_331),
.A2(n_249),
.B1(n_251),
.B2(n_246),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_324),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_315),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_323),
.Y(n_425)
);

OA21x2_ASAP7_75t_L g426 ( 
.A1(n_358),
.A2(n_270),
.B(n_266),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_332),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_315),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_358),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_323),
.B(n_245),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_356),
.A2(n_241),
.B1(n_252),
.B2(n_247),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_358),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_319),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_323),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_315),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_358),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_358),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_358),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_323),
.B(n_266),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_347),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_357),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_323),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_323),
.Y(n_443)
);

OAI21x1_ASAP7_75t_L g444 ( 
.A1(n_343),
.A2(n_274),
.B(n_270),
.Y(n_444)
);

AND2x6_ASAP7_75t_L g445 ( 
.A(n_316),
.B(n_160),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_357),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_358),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_389),
.Y(n_448)
);

AND3x1_ASAP7_75t_L g449 ( 
.A(n_410),
.B(n_157),
.C(n_129),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_396),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_447),
.Y(n_451)
);

CKINVDCx8_ASAP7_75t_R g452 ( 
.A(n_381),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_381),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_366),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_366),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_377),
.B(n_252),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_379),
.B(n_274),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_361),
.B(n_378),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_424),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_436),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_436),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_363),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_441),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_426),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_426),
.Y(n_465)
);

AND3x1_ASAP7_75t_L g466 ( 
.A(n_399),
.B(n_157),
.C(n_132),
.Y(n_466)
);

INVx6_ASAP7_75t_L g467 ( 
.A(n_364),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_424),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_361),
.B(n_275),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_418),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_365),
.A2(n_259),
.B1(n_137),
.B2(n_182),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_377),
.B(n_277),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_420),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_378),
.B(n_277),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_429),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_432),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_362),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_437),
.Y(n_478)
);

AND2x6_ASAP7_75t_L g479 ( 
.A(n_375),
.B(n_160),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_414),
.B(n_259),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_400),
.B(n_183),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_438),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_385),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_441),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_387),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_387),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_388),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_446),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_376),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_375),
.Y(n_490)
);

OA21x2_ASAP7_75t_L g491 ( 
.A1(n_371),
.A2(n_285),
.B(n_280),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_421),
.A2(n_159),
.B1(n_150),
.B2(n_182),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_375),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_382),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_386),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_386),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_383),
.B(n_391),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_386),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_383),
.B(n_280),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_403),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_379),
.B(n_285),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_489),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_500),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_464),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_494),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_453),
.Y(n_506)
);

NAND2xp33_ASAP7_75t_SL g507 ( 
.A(n_458),
.B(n_413),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_453),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_459),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_459),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_463),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_483),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_497),
.B(n_395),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_452),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_464),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_452),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_468),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_485),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_468),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_500),
.Y(n_520)
);

BUFx10_ASAP7_75t_L g521 ( 
.A(n_480),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_484),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_450),
.B(n_413),
.Y(n_523)
);

NOR2xp67_ASAP7_75t_L g524 ( 
.A(n_456),
.B(n_411),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_467),
.Y(n_525)
);

AND3x2_ASAP7_75t_L g526 ( 
.A(n_456),
.B(n_421),
.C(n_446),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_486),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_499),
.B(n_395),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_487),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_R g530 ( 
.A(n_467),
.B(n_428),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_465),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_462),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_488),
.B(n_416),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_467),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_465),
.Y(n_535)
);

OAI21x1_ASAP7_75t_L g536 ( 
.A1(n_491),
.A2(n_444),
.B(n_384),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_481),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_R g538 ( 
.A(n_448),
.B(n_428),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_471),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_448),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_502),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_504),
.Y(n_542)
);

OR2x6_ASAP7_75t_L g543 ( 
.A(n_524),
.B(n_409),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_540),
.Y(n_544)
);

NAND2xp33_ASAP7_75t_L g545 ( 
.A(n_538),
.B(n_513),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_504),
.Y(n_546)
);

NAND2xp33_ASAP7_75t_L g547 ( 
.A(n_530),
.B(n_448),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_540),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_515),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_528),
.B(n_392),
.Y(n_550)
);

BUFx10_ASAP7_75t_L g551 ( 
.A(n_508),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_505),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_520),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_533),
.B(n_393),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_540),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_540),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_515),
.Y(n_557)
);

AND3x2_ASAP7_75t_L g558 ( 
.A(n_511),
.B(n_480),
.C(n_503),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_523),
.B(n_431),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_532),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_512),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_517),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_507),
.B(n_369),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_517),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_518),
.Y(n_565)
);

BUFx4f_ASAP7_75t_L g566 ( 
.A(n_527),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_531),
.Y(n_567)
);

BUFx10_ASAP7_75t_L g568 ( 
.A(n_509),
.Y(n_568)
);

CKINVDCx16_ASAP7_75t_R g569 ( 
.A(n_506),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_531),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_522),
.B(n_407),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_507),
.B(n_391),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_521),
.B(n_399),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_529),
.B(n_412),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_535),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_519),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_535),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_536),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_521),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_536),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_521),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_526),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_539),
.A2(n_397),
.B1(n_419),
.B2(n_373),
.Y(n_583)
);

INVxp33_ASAP7_75t_SL g584 ( 
.A(n_510),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_514),
.B(n_423),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_516),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_525),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_534),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_539),
.B(n_394),
.Y(n_589)
);

INVx4_ASAP7_75t_L g590 ( 
.A(n_537),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_506),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_502),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_507),
.B(n_499),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_533),
.B(n_398),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_520),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_540),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_513),
.B(n_415),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_513),
.A2(n_397),
.B1(n_419),
.B2(n_492),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_530),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_504),
.Y(n_600)
);

CKINVDCx6p67_ASAP7_75t_R g601 ( 
.A(n_506),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_520),
.Y(n_602)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_540),
.Y(n_603)
);

OR2x6_ASAP7_75t_L g604 ( 
.A(n_524),
.B(n_409),
.Y(n_604)
);

NAND2xp33_ASAP7_75t_SL g605 ( 
.A(n_538),
.B(n_448),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_520),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_540),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_503),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_504),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_528),
.B(n_408),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_504),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_504),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_504),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_504),
.Y(n_614)
);

AO21x2_ASAP7_75t_L g615 ( 
.A1(n_536),
.A2(n_474),
.B(n_469),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_520),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_504),
.Y(n_617)
);

OA22x2_ASAP7_75t_L g618 ( 
.A1(n_526),
.A2(n_422),
.B1(n_415),
.B2(n_405),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_503),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_540),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_524),
.A2(n_435),
.B1(n_404),
.B2(n_433),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_520),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_524),
.A2(n_435),
.B1(n_400),
.B2(n_433),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_559),
.B(n_427),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_560),
.Y(n_625)
);

INVx4_ASAP7_75t_SL g626 ( 
.A(n_543),
.Y(n_626)
);

INVx4_ASAP7_75t_L g627 ( 
.A(n_599),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_544),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_541),
.Y(n_629)
);

BUFx10_ASAP7_75t_L g630 ( 
.A(n_576),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_544),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_552),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_544),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_566),
.B(n_368),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_569),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_566),
.B(n_411),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_601),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_573),
.B(n_466),
.Y(n_638)
);

INVx5_ASAP7_75t_L g639 ( 
.A(n_543),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_544),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_586),
.B(n_390),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_598),
.B(n_406),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_592),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_555),
.Y(n_644)
);

NAND3xp33_ASAP7_75t_L g645 ( 
.A(n_598),
.B(n_583),
.C(n_589),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_560),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_610),
.B(n_398),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_610),
.B(n_401),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_555),
.Y(n_649)
);

NOR2x1p5_ASAP7_75t_L g650 ( 
.A(n_597),
.B(n_380),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_561),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_565),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_595),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_562),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_575),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_542),
.Y(n_656)
);

AO21x2_ASAP7_75t_L g657 ( 
.A1(n_572),
.A2(n_473),
.B(n_470),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_621),
.B(n_406),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_577),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_546),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_546),
.Y(n_661)
);

BUFx4f_ASAP7_75t_L g662 ( 
.A(n_543),
.Y(n_662)
);

AND3x4_ASAP7_75t_L g663 ( 
.A(n_591),
.B(n_440),
.C(n_390),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_549),
.Y(n_664)
);

AND2x6_ASAP7_75t_L g665 ( 
.A(n_581),
.B(n_472),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_594),
.B(n_405),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_557),
.B(n_460),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_608),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_557),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_581),
.B(n_493),
.Y(n_670)
);

XNOR2x2_ASAP7_75t_L g671 ( 
.A(n_618),
.B(n_449),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_578),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_567),
.B(n_461),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_608),
.Y(n_674)
);

BUFx4f_ASAP7_75t_L g675 ( 
.A(n_604),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_567),
.B(n_461),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_584),
.B(n_440),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_585),
.B(n_409),
.Y(n_678)
);

AOI22x1_ASAP7_75t_L g679 ( 
.A1(n_582),
.A2(n_406),
.B1(n_430),
.B2(n_457),
.Y(n_679)
);

INVx6_ASAP7_75t_L g680 ( 
.A(n_551),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_589),
.B(n_402),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_619),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_570),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_570),
.B(n_451),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_600),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_600),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_583),
.A2(n_171),
.B1(n_178),
.B2(n_164),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_609),
.Y(n_688)
);

AND2x6_ASAP7_75t_L g689 ( 
.A(n_579),
.B(n_472),
.Y(n_689)
);

BUFx2_ASAP7_75t_L g690 ( 
.A(n_619),
.Y(n_690)
);

AO21x2_ASAP7_75t_L g691 ( 
.A1(n_572),
.A2(n_476),
.B(n_475),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_553),
.B(n_430),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_579),
.B(n_493),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_568),
.Y(n_694)
);

AO21x2_ASAP7_75t_L g695 ( 
.A1(n_593),
.A2(n_482),
.B(n_478),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_609),
.B(n_454),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_611),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_554),
.B(n_477),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_580),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_611),
.B(n_455),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_587),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_582),
.B(n_372),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_695),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_629),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_626),
.B(n_558),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_652),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_628),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_632),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_645),
.B(n_623),
.Y(n_709)
);

AO22x2_ASAP7_75t_L g710 ( 
.A1(n_645),
.A2(n_563),
.B1(n_593),
.B2(n_580),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_643),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_638),
.B(n_591),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_625),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_701),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_687),
.A2(n_663),
.B1(n_618),
.B2(n_681),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_651),
.Y(n_716)
);

INVx1_ASAP7_75t_SL g717 ( 
.A(n_690),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_655),
.B(n_558),
.Y(n_718)
);

NOR2x1p5_ASAP7_75t_L g719 ( 
.A(n_627),
.B(n_590),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_646),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_644),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_666),
.B(n_587),
.Y(n_722)
);

HB1xp67_ASAP7_75t_L g723 ( 
.A(n_695),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_628),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_626),
.B(n_588),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_662),
.B(n_588),
.Y(n_726)
);

NAND3xp33_ASAP7_75t_L g727 ( 
.A(n_687),
.B(n_563),
.C(n_545),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_656),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_630),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_672),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_672),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_659),
.Y(n_732)
);

AND2x6_ASAP7_75t_L g733 ( 
.A(n_693),
.B(n_555),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_628),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_639),
.B(n_548),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_664),
.Y(n_736)
);

A2O1A1Ixp33_ASAP7_75t_L g737 ( 
.A1(n_642),
.A2(n_545),
.B(n_605),
.C(n_547),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_680),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_631),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_669),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_683),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_680),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_653),
.Y(n_743)
);

CKINVDCx16_ASAP7_75t_R g744 ( 
.A(n_635),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_631),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_657),
.Y(n_746)
);

AOI22x1_ASAP7_75t_L g747 ( 
.A1(n_650),
.A2(n_564),
.B1(n_606),
.B2(n_602),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_660),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_685),
.Y(n_749)
);

INVx4_ASAP7_75t_L g750 ( 
.A(n_639),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_637),
.Y(n_751)
);

NAND3xp33_ASAP7_75t_L g752 ( 
.A(n_679),
.B(n_550),
.C(n_571),
.Y(n_752)
);

INVx4_ASAP7_75t_L g753 ( 
.A(n_639),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_688),
.B(n_612),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_661),
.Y(n_755)
);

INVx8_ASAP7_75t_L g756 ( 
.A(n_631),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_624),
.B(n_616),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_657),
.B(n_612),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_662),
.B(n_605),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_647),
.B(n_622),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_654),
.Y(n_761)
);

OAI22xp33_ASAP7_75t_L g762 ( 
.A1(n_675),
.A2(n_604),
.B1(n_574),
.B2(n_590),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_686),
.Y(n_763)
);

AO22x2_ASAP7_75t_L g764 ( 
.A1(n_658),
.A2(n_614),
.B1(n_617),
.B2(n_613),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_697),
.Y(n_765)
);

NAND3xp33_ASAP7_75t_L g766 ( 
.A(n_648),
.B(n_571),
.C(n_547),
.Y(n_766)
);

AND2x6_ASAP7_75t_L g767 ( 
.A(n_693),
.B(n_555),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_668),
.B(n_548),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_699),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_674),
.B(n_556),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_675),
.B(n_568),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_682),
.B(n_556),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_704),
.Y(n_773)
);

NAND3xp33_ASAP7_75t_SL g774 ( 
.A(n_709),
.B(n_634),
.C(n_641),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_737),
.A2(n_636),
.B(n_691),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_708),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_713),
.B(n_698),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_752),
.B(n_694),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_717),
.B(n_678),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_744),
.B(n_702),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_727),
.A2(n_715),
.B1(n_762),
.B2(n_759),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_743),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_738),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_706),
.B(n_665),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_712),
.B(n_677),
.Y(n_785)
);

O2A1O1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_715),
.A2(n_671),
.B(n_604),
.C(n_178),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_711),
.B(n_665),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_744),
.B(n_627),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_727),
.A2(n_692),
.B1(n_665),
.B2(n_689),
.Y(n_789)
);

O2A1O1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_752),
.A2(n_164),
.B(n_131),
.C(n_136),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_716),
.Y(n_791)
);

BUFx8_ASAP7_75t_L g792 ( 
.A(n_742),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_732),
.B(n_720),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_705),
.B(n_670),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_718),
.B(n_736),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_718),
.B(n_740),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_730),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_741),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_749),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_757),
.B(n_372),
.Y(n_800)
);

BUFx5_ASAP7_75t_L g801 ( 
.A(n_733),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_707),
.Y(n_802)
);

NAND2xp33_ASAP7_75t_L g803 ( 
.A(n_719),
.B(n_689),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_705),
.B(n_670),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_714),
.B(n_665),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_728),
.Y(n_806)
);

BUFx8_ASAP7_75t_L g807 ( 
.A(n_729),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_726),
.B(n_644),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_771),
.B(n_633),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_748),
.Y(n_810)
);

AND2x6_ASAP7_75t_L g811 ( 
.A(n_725),
.B(n_633),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_766),
.A2(n_689),
.B1(n_445),
.B2(n_479),
.Y(n_812)
);

NOR3xp33_ASAP7_75t_L g813 ( 
.A(n_766),
.B(n_603),
.C(n_596),
.Y(n_813)
);

AND2x6_ASAP7_75t_SL g814 ( 
.A(n_725),
.B(n_126),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_710),
.A2(n_596),
.B1(n_603),
.B2(n_649),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_731),
.B(n_649),
.Y(n_816)
);

OAI221xp5_ASAP7_75t_L g817 ( 
.A1(n_747),
.A2(n_174),
.B1(n_173),
.B2(n_143),
.C(n_144),
.Y(n_817)
);

OR2x6_ASAP7_75t_L g818 ( 
.A(n_750),
.B(n_640),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_714),
.B(n_689),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_755),
.B(n_615),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_769),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_710),
.A2(n_445),
.B1(n_479),
.B2(n_457),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_763),
.B(n_684),
.Y(n_823)
);

INVx4_ASAP7_75t_L g824 ( 
.A(n_707),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_750),
.B(n_640),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_753),
.B(n_640),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_765),
.B(n_684),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_753),
.B(n_607),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_761),
.B(n_607),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_707),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_764),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_754),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_760),
.B(n_146),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_735),
.B(n_607),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_735),
.B(n_607),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_751),
.B(n_722),
.Y(n_836)
);

INVxp33_ASAP7_75t_L g837 ( 
.A(n_770),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_768),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_768),
.A2(n_133),
.B1(n_445),
.B2(n_171),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_SL g840 ( 
.A(n_772),
.B(n_756),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_754),
.B(n_696),
.Y(n_841)
);

OR2x2_ASAP7_75t_L g842 ( 
.A(n_758),
.B(n_696),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_721),
.B(n_620),
.Y(n_843)
);

BUFx6f_ASAP7_75t_SL g844 ( 
.A(n_724),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_758),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_SL g846 ( 
.A(n_756),
.B(n_367),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_756),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_773),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_845),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_831),
.B(n_703),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_795),
.B(n_723),
.Y(n_851)
);

CKINVDCx8_ASAP7_75t_R g852 ( 
.A(n_814),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_837),
.B(n_746),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_796),
.B(n_777),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_816),
.B(n_703),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_778),
.A2(n_721),
.B(n_162),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_783),
.Y(n_857)
);

INVx4_ASAP7_75t_L g858 ( 
.A(n_783),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_816),
.B(n_724),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_832),
.B(n_724),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_791),
.Y(n_861)
);

INVxp67_ASAP7_75t_L g862 ( 
.A(n_785),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_781),
.B(n_734),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_821),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_797),
.B(n_734),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_779),
.B(n_739),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_776),
.B(n_739),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_783),
.Y(n_868)
);

AND2x4_ASAP7_75t_SL g869 ( 
.A(n_813),
.B(n_739),
.Y(n_869)
);

NAND2xp33_ASAP7_75t_SL g870 ( 
.A(n_844),
.B(n_745),
.Y(n_870)
);

NOR2x1p5_ASAP7_75t_L g871 ( 
.A(n_774),
.B(n_782),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_793),
.B(n_745),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_792),
.Y(n_873)
);

AND2x2_ASAP7_75t_SL g874 ( 
.A(n_803),
.B(n_745),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_798),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_799),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_806),
.Y(n_877)
);

INVx4_ASAP7_75t_L g878 ( 
.A(n_802),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_842),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_810),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_788),
.B(n_620),
.Y(n_881)
);

AND2x2_ASAP7_75t_SL g882 ( 
.A(n_822),
.B(n_177),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_820),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_823),
.Y(n_884)
);

INVx1_ASAP7_75t_SL g885 ( 
.A(n_838),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_787),
.B(n_733),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_805),
.B(n_733),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_800),
.B(n_147),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_784),
.B(n_733),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_802),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_827),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_825),
.B(n_767),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_836),
.B(n_819),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_826),
.B(n_767),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_802),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_815),
.B(n_767),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_841),
.B(n_767),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_790),
.A2(n_169),
.B(n_163),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_792),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_882),
.A2(n_789),
.B1(n_812),
.B2(n_786),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_874),
.B(n_775),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_882),
.A2(n_804),
.B1(n_794),
.B2(n_780),
.Y(n_902)
);

AOI21xp33_ASAP7_75t_L g903 ( 
.A1(n_888),
.A2(n_833),
.B(n_808),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_887),
.B(n_834),
.Y(n_904)
);

A2O1A1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_871),
.A2(n_817),
.B(n_809),
.C(n_840),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_870),
.A2(n_828),
.B(n_843),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_889),
.B(n_887),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_870),
.A2(n_835),
.B(n_829),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_852),
.A2(n_847),
.B1(n_818),
.B2(n_824),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_884),
.B(n_891),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_884),
.B(n_811),
.Y(n_911)
);

INVx4_ASAP7_75t_L g912 ( 
.A(n_873),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_856),
.A2(n_874),
.B(n_863),
.Y(n_913)
);

NOR2xp67_ASAP7_75t_L g914 ( 
.A(n_858),
.B(n_830),
.Y(n_914)
);

NOR2x1_ASAP7_75t_R g915 ( 
.A(n_873),
.B(n_801),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_889),
.B(n_801),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_858),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_898),
.A2(n_176),
.B(n_818),
.C(n_839),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_864),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_852),
.A2(n_899),
.B(n_869),
.C(n_881),
.Y(n_920)
);

OAI21xp33_ASAP7_75t_L g921 ( 
.A1(n_854),
.A2(n_846),
.B(n_179),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_879),
.B(n_811),
.Y(n_922)
);

NAND2xp33_ASAP7_75t_L g923 ( 
.A(n_857),
.B(n_801),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_857),
.B(n_801),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_899),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_851),
.A2(n_700),
.B(n_667),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_897),
.B(n_807),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_857),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_855),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_858),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_869),
.A2(n_894),
.B(n_892),
.Y(n_931)
);

INVxp67_ASAP7_75t_L g932 ( 
.A(n_865),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_892),
.A2(n_676),
.B(n_673),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_886),
.A2(n_479),
.B1(n_617),
.B2(n_614),
.Y(n_934)
);

INVx1_ASAP7_75t_SL g935 ( 
.A(n_885),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_892),
.A2(n_894),
.B(n_886),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_859),
.B(n_855),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_872),
.A2(n_177),
.B(n_370),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_862),
.B(n_479),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_857),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_853),
.B(n_479),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_893),
.A2(n_896),
.B(n_853),
.C(n_857),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_848),
.B(n_0),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_883),
.B(n_0),
.Y(n_944)
);

INVx2_ASAP7_75t_SL g945 ( 
.A(n_868),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_883),
.A2(n_370),
.B(n_179),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_867),
.B(n_1),
.Y(n_947)
);

NAND3xp33_ASAP7_75t_L g948 ( 
.A(n_850),
.B(n_180),
.C(n_128),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_867),
.B(n_877),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_877),
.B(n_2),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_932),
.B(n_866),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_901),
.A2(n_850),
.B(n_896),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_912),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_944),
.B(n_866),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_907),
.B(n_850),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_925),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_902),
.A2(n_868),
.B1(n_859),
.B2(n_878),
.Y(n_957)
);

OR2x6_ASAP7_75t_L g958 ( 
.A(n_925),
.B(n_868),
.Y(n_958)
);

INVx4_ASAP7_75t_L g959 ( 
.A(n_925),
.Y(n_959)
);

NOR2xp67_ASAP7_75t_L g960 ( 
.A(n_931),
.B(n_849),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_L g961 ( 
.A1(n_905),
.A2(n_880),
.B(n_860),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_933),
.B(n_860),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_900),
.A2(n_909),
.B1(n_913),
.B2(n_916),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_903),
.A2(n_868),
.B1(n_878),
.B2(n_890),
.Y(n_964)
);

NOR3xp33_ASAP7_75t_L g965 ( 
.A(n_948),
.B(n_878),
.C(n_880),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_946),
.A2(n_868),
.B(n_861),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_928),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_942),
.A2(n_876),
.B(n_875),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_923),
.A2(n_876),
.B(n_875),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_920),
.B(n_890),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_954),
.B(n_965),
.Y(n_971)
);

AO22x1_ASAP7_75t_L g972 ( 
.A1(n_953),
.A2(n_935),
.B1(n_917),
.B2(n_930),
.Y(n_972)
);

O2A1O1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_970),
.A2(n_943),
.B(n_950),
.C(n_938),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_963),
.A2(n_915),
.B(n_924),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_961),
.A2(n_906),
.B(n_918),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_955),
.B(n_949),
.Y(n_976)
);

INVx4_ASAP7_75t_L g977 ( 
.A(n_956),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_951),
.Y(n_978)
);

INVxp67_ASAP7_75t_L g979 ( 
.A(n_956),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_967),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_959),
.Y(n_981)
);

NOR3xp33_ASAP7_75t_L g982 ( 
.A(n_957),
.B(n_921),
.C(n_947),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_958),
.A2(n_936),
.B1(n_934),
.B2(n_904),
.Y(n_983)
);

INVxp67_ASAP7_75t_L g984 ( 
.A(n_967),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_962),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_960),
.B(n_968),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_952),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_966),
.B(n_937),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_964),
.A2(n_939),
.B(n_941),
.C(n_945),
.Y(n_989)
);

AND2x6_ASAP7_75t_L g990 ( 
.A(n_969),
.B(n_928),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_954),
.B(n_929),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_954),
.B(n_910),
.Y(n_992)
);

OAI22xp33_ASAP7_75t_L g993 ( 
.A1(n_963),
.A2(n_908),
.B1(n_922),
.B2(n_911),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_963),
.A2(n_914),
.B(n_927),
.C(n_926),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_959),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_991),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_995),
.B(n_977),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_978),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_992),
.B(n_919),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_975),
.A2(n_986),
.B1(n_993),
.B2(n_985),
.Y(n_1000)
);

INVx4_ASAP7_75t_L g1001 ( 
.A(n_981),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_979),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_980),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_SL g1004 ( 
.A(n_997),
.B(n_987),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_1001),
.B(n_984),
.Y(n_1005)
);

INVxp67_ASAP7_75t_SL g1006 ( 
.A(n_1000),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_1006),
.A2(n_994),
.B(n_971),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_1005),
.Y(n_1008)
);

AO31x2_ASAP7_75t_L g1009 ( 
.A1(n_1007),
.A2(n_1001),
.A3(n_1003),
.B(n_998),
.Y(n_1009)
);

AO31x2_ASAP7_75t_L g1010 ( 
.A1(n_1008),
.A2(n_1004),
.A3(n_996),
.B(n_974),
.Y(n_1010)
);

OR2x2_ASAP7_75t_L g1011 ( 
.A(n_1009),
.B(n_999),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_1009),
.Y(n_1012)
);

OR2x2_ASAP7_75t_L g1013 ( 
.A(n_1011),
.B(n_1010),
.Y(n_1013)
);

NAND3xp33_ASAP7_75t_SL g1014 ( 
.A(n_1012),
.B(n_1002),
.C(n_982),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1013),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_1014),
.Y(n_1016)
);

INVxp67_ASAP7_75t_L g1017 ( 
.A(n_1015),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_1016),
.B(n_986),
.Y(n_1018)
);

OR2x2_ASAP7_75t_L g1019 ( 
.A(n_1017),
.B(n_999),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_1018),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_1017),
.B(n_976),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1021),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_1020),
.B(n_988),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_1019),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_1023),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_1024),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_1026),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_1025),
.B(n_1022),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1028),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_1027),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_1030),
.Y(n_1031)
);

INVx1_ASAP7_75t_SL g1032 ( 
.A(n_1029),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1031),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_1032),
.Y(n_1034)
);

BUFx2_ASAP7_75t_L g1035 ( 
.A(n_1034),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_1033),
.B(n_972),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1036),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_1035),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_1035),
.Y(n_1039)
);

INVx4_ASAP7_75t_L g1040 ( 
.A(n_1038),
.Y(n_1040)
);

INVx2_ASAP7_75t_SL g1041 ( 
.A(n_1039),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1037),
.B(n_990),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_1041),
.A2(n_990),
.B1(n_983),
.B2(n_928),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_1042),
.B(n_990),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_1044),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1043),
.B(n_1040),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_1045),
.B(n_940),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1046),
.B(n_2),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_1047),
.B(n_973),
.Y(n_1049)
);

INVx1_ASAP7_75t_SL g1050 ( 
.A(n_1048),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1050),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1049),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_1051),
.A2(n_180),
.B(n_128),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_1052),
.B(n_3),
.Y(n_1054)
);

OAI222xp33_ASAP7_75t_L g1055 ( 
.A1(n_1054),
.A2(n_374),
.B1(n_989),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1053),
.Y(n_1056)
);

AO21x1_ASAP7_75t_L g1057 ( 
.A1(n_1053),
.A2(n_3),
.B(n_5),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1057),
.Y(n_1058)
);

AOI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_1056),
.A2(n_367),
.B1(n_417),
.B2(n_425),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_1055),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1058),
.B(n_1060),
.Y(n_1061)
);

INVx2_ASAP7_75t_SL g1062 ( 
.A(n_1059),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1062),
.B(n_8),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_1061),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1064),
.Y(n_1065)
);

AOI211xp5_ASAP7_75t_L g1066 ( 
.A1(n_1063),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1065),
.Y(n_1067)
);

NOR2x1_ASAP7_75t_L g1068 ( 
.A(n_1066),
.B(n_374),
.Y(n_1068)
);

INVxp67_ASAP7_75t_SL g1069 ( 
.A(n_1067),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1068),
.Y(n_1070)
);

NAND3xp33_ASAP7_75t_SL g1071 ( 
.A(n_1070),
.B(n_9),
.C(n_10),
.Y(n_1071)
);

OAI21xp33_ASAP7_75t_L g1072 ( 
.A1(n_1069),
.A2(n_281),
.B(n_279),
.Y(n_1072)
);

NOR3xp33_ASAP7_75t_L g1073 ( 
.A(n_1072),
.B(n_12),
.C(n_13),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1071),
.B(n_12),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_1072),
.A2(n_443),
.B1(n_442),
.B2(n_434),
.Y(n_1075)
);

NAND4xp25_ASAP7_75t_L g1076 ( 
.A(n_1074),
.B(n_13),
.C(n_15),
.D(n_16),
.Y(n_1076)
);

NAND4xp25_ASAP7_75t_L g1077 ( 
.A(n_1073),
.B(n_15),
.C(n_16),
.D(n_17),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1075),
.B(n_17),
.Y(n_1078)
);

NOR2x1_ASAP7_75t_L g1079 ( 
.A(n_1077),
.B(n_367),
.Y(n_1079)
);

NOR2x1_ASAP7_75t_L g1080 ( 
.A(n_1078),
.B(n_417),
.Y(n_1080)
);

NAND3xp33_ASAP7_75t_SL g1081 ( 
.A(n_1079),
.B(n_1076),
.C(n_18),
.Y(n_1081)
);

NOR5xp2_ASAP7_75t_L g1082 ( 
.A(n_1080),
.B(n_18),
.C(n_19),
.D(n_20),
.E(n_21),
.Y(n_1082)
);

NOR2x1_ASAP7_75t_L g1083 ( 
.A(n_1081),
.B(n_417),
.Y(n_1083)
);

NAND4xp75_ASAP7_75t_L g1084 ( 
.A(n_1082),
.B(n_19),
.C(n_20),
.D(n_21),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1083),
.Y(n_1085)
);

AOI31xp33_ASAP7_75t_L g1086 ( 
.A1(n_1084),
.A2(n_22),
.A3(n_23),
.B(n_25),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1085),
.Y(n_1087)
);

NAND4xp25_ASAP7_75t_SL g1088 ( 
.A(n_1086),
.B(n_22),
.C(n_23),
.D(n_25),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1087),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1088),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_1089),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_1090),
.Y(n_1092)
);

XNOR2x1_ASAP7_75t_L g1093 ( 
.A(n_1089),
.B(n_26),
.Y(n_1093)
);

XOR2xp5_ASAP7_75t_L g1094 ( 
.A(n_1092),
.B(n_27),
.Y(n_1094)
);

AO211x2_ASAP7_75t_L g1095 ( 
.A1(n_1091),
.A2(n_28),
.B(n_31),
.C(n_33),
.Y(n_1095)
);

CKINVDCx20_ASAP7_75t_R g1096 ( 
.A(n_1093),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1096),
.Y(n_1097)
);

INVxp67_ASAP7_75t_L g1098 ( 
.A(n_1094),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1097),
.B(n_1095),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_1098),
.A2(n_425),
.B1(n_434),
.B2(n_442),
.Y(n_1100)
);

NOR3xp33_ASAP7_75t_SL g1101 ( 
.A(n_1099),
.B(n_34),
.C(n_35),
.Y(n_1101)
);

XNOR2xp5_ASAP7_75t_L g1102 ( 
.A(n_1100),
.B(n_36),
.Y(n_1102)
);

NOR3xp33_ASAP7_75t_L g1103 ( 
.A(n_1101),
.B(n_1102),
.C(n_288),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_1101),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1104),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1103),
.Y(n_1106)
);

NOR2x1p5_ASAP7_75t_L g1107 ( 
.A(n_1106),
.B(n_425),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_1105),
.A2(n_434),
.B1(n_442),
.B2(n_443),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1107),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1108),
.A2(n_940),
.B1(n_443),
.B2(n_439),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_1107),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1109),
.A2(n_940),
.B1(n_895),
.B2(n_890),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1111),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1110),
.Y(n_1114)
);

AOI31xp33_ASAP7_75t_L g1115 ( 
.A1(n_1109),
.A2(n_439),
.A3(n_40),
.B(n_42),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1113),
.B(n_39),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1114),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1115),
.A2(n_895),
.B1(n_890),
.B2(n_498),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1117),
.A2(n_1112),
.B1(n_895),
.B2(n_890),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1118),
.A2(n_895),
.B(n_501),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1116),
.B(n_44),
.Y(n_1121)
);

NAND3xp33_ASAP7_75t_L g1122 ( 
.A(n_1120),
.B(n_895),
.C(n_495),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1121),
.A2(n_45),
.B(n_47),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1119),
.A2(n_48),
.B(n_50),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1120),
.B(n_54),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1120),
.A2(n_55),
.B(n_56),
.Y(n_1126)
);

AOI221xp5_ASAP7_75t_L g1127 ( 
.A1(n_1120),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.C(n_60),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1120),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1120),
.Y(n_1129)
);

AO221x1_ASAP7_75t_L g1130 ( 
.A1(n_1120),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.C(n_65),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1120),
.A2(n_501),
.B1(n_498),
.B2(n_496),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1120),
.B(n_67),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1120),
.A2(n_68),
.B(n_69),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1128),
.Y(n_1134)
);

INVxp67_ASAP7_75t_L g1135 ( 
.A(n_1129),
.Y(n_1135)
);

INVxp67_ASAP7_75t_SL g1136 ( 
.A(n_1122),
.Y(n_1136)
);

NOR2x1_ASAP7_75t_L g1137 ( 
.A(n_1125),
.B(n_501),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1132),
.Y(n_1138)
);

INVxp67_ASAP7_75t_SL g1139 ( 
.A(n_1131),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1130),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_1126),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1133),
.B(n_1124),
.Y(n_1142)
);

INVx4_ASAP7_75t_L g1143 ( 
.A(n_1134),
.Y(n_1143)
);

OA21x2_ASAP7_75t_L g1144 ( 
.A1(n_1135),
.A2(n_1123),
.B(n_1127),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1140),
.A2(n_498),
.B1(n_496),
.B2(n_495),
.Y(n_1145)
);

AOI32xp33_ASAP7_75t_L g1146 ( 
.A1(n_1141),
.A2(n_70),
.A3(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_SL g1147 ( 
.A1(n_1138),
.A2(n_1142),
.B1(n_1139),
.B2(n_1136),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_1137),
.A2(n_498),
.B1(n_496),
.B2(n_495),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_SL g1149 ( 
.A1(n_1143),
.A2(n_496),
.B1(n_495),
.B2(n_490),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1147),
.B(n_75),
.Y(n_1150)
);

AOI21xp33_ASAP7_75t_L g1151 ( 
.A1(n_1144),
.A2(n_76),
.B(n_77),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1148),
.B(n_79),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_SL g1153 ( 
.A1(n_1152),
.A2(n_1146),
.B1(n_1145),
.B2(n_83),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1153),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_1154),
.B(n_1150),
.Y(n_1155)
);

OAI221xp5_ASAP7_75t_R g1156 ( 
.A1(n_1155),
.A2(n_1151),
.B1(n_1149),
.B2(n_84),
.C(n_85),
.Y(n_1156)
);

AOI221xp5_ASAP7_75t_L g1157 ( 
.A1(n_1156),
.A2(n_81),
.B1(n_82),
.B2(n_87),
.C(n_89),
.Y(n_1157)
);

AOI21xp33_ASAP7_75t_L g1158 ( 
.A1(n_1157),
.A2(n_91),
.B(n_92),
.Y(n_1158)
);

AOI211xp5_ASAP7_75t_L g1159 ( 
.A1(n_1158),
.A2(n_93),
.B(n_95),
.C(n_96),
.Y(n_1159)
);

AOI211xp5_ASAP7_75t_L g1160 ( 
.A1(n_1159),
.A2(n_97),
.B(n_98),
.C(n_99),
.Y(n_1160)
);


endmodule