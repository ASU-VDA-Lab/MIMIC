module fake_ariane_3338_n_1252 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1252);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1252;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_423;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_187;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_232;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_200;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_868;
wire n_884;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_238;
wire n_365;
wire n_1013;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_440;
wire n_273;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_461;
wire n_1121;
wire n_490;
wire n_209;
wire n_225;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_555;
wire n_804;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_513;
wire n_288;
wire n_179;
wire n_1178;
wire n_1026;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_746;
wire n_292;
wire n_1079;
wire n_615;
wire n_1139;
wire n_517;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_299;
wire n_836;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_776;
wire n_424;
wire n_466;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_553;
wire n_814;
wire n_578;
wire n_405;
wire n_320;
wire n_1134;
wire n_647;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_218;
wire n_247;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_233;
wire n_957;
wire n_388;
wire n_1242;
wire n_1218;
wire n_321;
wire n_221;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_845;
wire n_888;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_769;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_999;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1243;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_317;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_687;
wire n_797;
wire n_480;
wire n_642;
wire n_211;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_516;
wire n_1137;
wire n_197;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_752;
wire n_985;
wire n_421;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_649;
wire n_374;
wire n_643;
wire n_226;
wire n_682;
wire n_819;
wire n_586;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_272;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_224;
wire n_894;
wire n_420;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_168;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_181;
wire n_617;
wire n_543;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_613;
wire n_1022;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_213;
wire n_1014;
wire n_724;
wire n_493;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_981;
wire n_1110;
wire n_243;
wire n_185;
wire n_1204;
wire n_994;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_828;
wire n_322;
wire n_558;
wire n_653;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1167;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_244;
wire n_679;
wire n_220;
wire n_663;
wire n_443;
wire n_528;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_385;
wire n_917;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1064;
wire n_633;
wire n_900;
wire n_1093;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_835;
wire n_446;
wire n_1076;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_188;
wire n_323;
wire n_550;
wire n_997;
wire n_635;
wire n_694;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1236;
wire n_228;
wire n_671;
wire n_1148;
wire n_654;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_196;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1229;
wire n_415;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_895;
wire n_304;
wire n_583;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_265;
wire n_208;
wire n_174;
wire n_275;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_963;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1001;
wire n_1115;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_250;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_573;
wire n_796;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_15),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_147),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_9),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_6),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_157),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_139),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_115),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_110),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_3),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_39),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_109),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_145),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

CKINVDCx12_ASAP7_75t_R g184 ( 
.A(n_158),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_166),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_48),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_26),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_150),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_123),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_20),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_132),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_106),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_54),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_131),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_36),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_129),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_72),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_11),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_124),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_13),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_66),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_15),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_45),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_62),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_85),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_128),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_103),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_2),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_120),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_100),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_138),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_10),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_149),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_96),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_95),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_1),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_46),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_36),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_125),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_33),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_156),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_140),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_59),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_40),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_7),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_38),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_154),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_46),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_70),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_113),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_19),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_114),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_101),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_33),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_8),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_13),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_164),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_84),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_43),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_82),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_81),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_83),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_146),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_151),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_104),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_68),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_99),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_116),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_122),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_64),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_148),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_163),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_0),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_67),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_71),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_39),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_141),
.Y(n_260)
);

BUFx2_ASAP7_75t_SL g261 ( 
.A(n_19),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_86),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_60),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_88),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_102),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_126),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_165),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_42),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_43),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_142),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_77),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_162),
.Y(n_272)
);

BUFx5_ASAP7_75t_L g273 ( 
.A(n_34),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_152),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_161),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_35),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_135),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_45),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_31),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_137),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_136),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_61),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_14),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_50),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_143),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_94),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_105),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

INVxp67_ASAP7_75t_SL g290 ( 
.A(n_210),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_205),
.Y(n_291)
);

INVxp33_ASAP7_75t_L g292 ( 
.A(n_200),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_266),
.B(n_0),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_273),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_168),
.Y(n_296)
);

INVxp33_ASAP7_75t_SL g297 ( 
.A(n_173),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_273),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_273),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_262),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_208),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_208),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_227),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_178),
.B(n_1),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_254),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_268),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_236),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_233),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_233),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_282),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_279),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_236),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_261),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_202),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_174),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_182),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_175),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_259),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_176),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_178),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_180),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_183),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_185),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_167),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_194),
.B(n_2),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_182),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_197),
.B(n_3),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_199),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_201),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_285),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_L g332 ( 
.A(n_167),
.B(n_4),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_186),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_186),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_213),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_254),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_179),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_196),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_219),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_196),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_225),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_187),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_230),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_240),
.B(n_4),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_241),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_247),
.B(n_5),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_187),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_270),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_257),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_287),
.B(n_5),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_238),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_258),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_267),
.Y(n_353)
);

INVxp33_ASAP7_75t_L g354 ( 
.A(n_248),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_238),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_256),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_284),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_271),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_256),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_278),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_270),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_275),
.B(n_6),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_274),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_274),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_277),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_284),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_278),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_280),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_277),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_281),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_184),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_169),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_170),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_179),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_204),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_204),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_239),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_177),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_288),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_289),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_293),
.Y(n_381)
);

CKINVDCx14_ASAP7_75t_R g382 ( 
.A(n_371),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_295),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_298),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_357),
.B(n_177),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_315),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_299),
.Y(n_387)
);

INVx6_ASAP7_75t_L g388 ( 
.A(n_306),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_301),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_309),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_309),
.Y(n_391)
);

BUFx8_ASAP7_75t_L g392 ( 
.A(n_325),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_310),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_310),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_370),
.Y(n_395)
);

BUFx8_ASAP7_75t_L g396 ( 
.A(n_325),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_370),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_357),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_354),
.B(n_239),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_326),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_316),
.Y(n_401)
);

AND2x4_ASAP7_75t_L g402 ( 
.A(n_306),
.B(n_272),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_318),
.B(n_272),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_320),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_331),
.B(n_297),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_322),
.Y(n_406)
);

OR2x6_ASAP7_75t_L g407 ( 
.A(n_332),
.B(n_248),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_323),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_324),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_329),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_328),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_330),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_335),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_339),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_341),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_343),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_345),
.Y(n_417)
);

AND2x6_ASAP7_75t_L g418 ( 
.A(n_349),
.B(n_250),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_352),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_353),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_358),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_368),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_377),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_378),
.B(n_242),
.Y(n_424)
);

BUFx12f_ASAP7_75t_L g425 ( 
.A(n_291),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_304),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_307),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_344),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_290),
.B(n_242),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_346),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_312),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_350),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_314),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_337),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_362),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_336),
.B(n_276),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_294),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_366),
.Y(n_438)
);

AND2x6_ASAP7_75t_L g439 ( 
.A(n_374),
.B(n_250),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_375),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_376),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_317),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_317),
.Y(n_443)
);

OA21x2_ASAP7_75t_L g444 ( 
.A1(n_311),
.A2(n_251),
.B(n_191),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_327),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_327),
.B(n_181),
.Y(n_446)
);

OA21x2_ASAP7_75t_L g447 ( 
.A1(n_311),
.A2(n_251),
.B(n_214),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_333),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_380),
.Y(n_449)
);

OR2x6_ASAP7_75t_L g450 ( 
.A(n_407),
.B(n_305),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_386),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_380),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_379),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_379),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_381),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_441),
.B(n_333),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_428),
.A2(n_297),
.B1(n_347),
.B2(n_369),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_388),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_381),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_442),
.B(n_334),
.Y(n_460)
);

INVx5_ASAP7_75t_L g461 ( 
.A(n_379),
.Y(n_461)
);

INVxp33_ASAP7_75t_L g462 ( 
.A(n_431),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_441),
.B(n_430),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_442),
.B(n_334),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_379),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_388),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_383),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_398),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_428),
.A2(n_292),
.B1(n_373),
.B2(n_372),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_379),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_431),
.B(n_319),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_398),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_441),
.B(n_342),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_L g474 ( 
.A1(n_432),
.A2(n_435),
.B1(n_447),
.B2(n_444),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_398),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_442),
.B(n_342),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_388),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_446),
.B(n_291),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_441),
.B(n_347),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_446),
.B(n_296),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_383),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_443),
.B(n_296),
.Y(n_482)
);

OR2x6_ASAP7_75t_L g483 ( 
.A(n_407),
.B(n_305),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_399),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_399),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_379),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_384),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_388),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_388),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_384),
.Y(n_490)
);

NAND3xp33_ASAP7_75t_L g491 ( 
.A(n_430),
.B(n_361),
.C(n_348),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_432),
.A2(n_276),
.B1(n_237),
.B2(n_220),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_384),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_440),
.Y(n_494)
);

AO22x2_ASAP7_75t_L g495 ( 
.A1(n_435),
.A2(n_216),
.B1(n_244),
.B2(n_264),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_384),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_384),
.Y(n_497)
);

CKINVDCx6p67_ASAP7_75t_R g498 ( 
.A(n_425),
.Y(n_498)
);

NAND3xp33_ASAP7_75t_L g499 ( 
.A(n_430),
.B(n_389),
.C(n_387),
.Y(n_499)
);

INVx6_ASAP7_75t_L g500 ( 
.A(n_440),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_443),
.B(n_300),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_442),
.B(n_348),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_430),
.B(n_400),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_384),
.Y(n_504)
);

AND2x6_ASAP7_75t_L g505 ( 
.A(n_442),
.B(n_198),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_391),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_391),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_398),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_398),
.Y(n_509)
);

BUFx8_ASAP7_75t_SL g510 ( 
.A(n_425),
.Y(n_510)
);

OR2x6_ASAP7_75t_L g511 ( 
.A(n_407),
.B(n_198),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_436),
.Y(n_512)
);

BUFx6f_ASAP7_75t_SL g513 ( 
.A(n_442),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_387),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_445),
.B(n_300),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_389),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_395),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_445),
.B(n_361),
.Y(n_518)
);

INVx1_ASAP7_75t_SL g519 ( 
.A(n_423),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_480),
.B(n_478),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_458),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_512),
.A2(n_437),
.B1(n_448),
.B2(n_430),
.Y(n_522)
);

INVx4_ASAP7_75t_L g523 ( 
.A(n_513),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_491),
.B(n_448),
.Y(n_524)
);

AO221x1_ASAP7_75t_L g525 ( 
.A1(n_495),
.A2(n_448),
.B1(n_437),
.B2(n_434),
.C(n_430),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_449),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_495),
.A2(n_439),
.B1(n_447),
.B2(n_444),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_517),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_512),
.A2(n_518),
.B1(n_484),
.B2(n_485),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_517),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_484),
.A2(n_437),
.B1(n_448),
.B2(n_411),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_491),
.B(n_448),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_456),
.B(n_448),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_485),
.A2(n_437),
.B1(n_411),
.B2(n_400),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_519),
.B(n_313),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_513),
.Y(n_536)
);

NAND3xp33_ASAP7_75t_L g537 ( 
.A(n_469),
.B(n_457),
.C(n_482),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_495),
.A2(n_439),
.B1(n_447),
.B2(n_444),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_458),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_473),
.B(n_437),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_479),
.B(n_437),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_460),
.B(n_438),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_449),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_452),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_462),
.B(n_424),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_519),
.B(n_313),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_452),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_451),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_474),
.B(n_438),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_463),
.B(n_400),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_501),
.B(n_400),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_SL g552 ( 
.A(n_498),
.B(n_392),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_466),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_451),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_515),
.B(n_400),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_466),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_455),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_455),
.B(n_400),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_459),
.B(n_411),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_459),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_467),
.B(n_411),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_467),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_481),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_481),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_514),
.B(n_411),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_514),
.B(n_411),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_516),
.Y(n_567)
);

NAND2x1_ASAP7_75t_L g568 ( 
.A(n_500),
.B(n_494),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_503),
.B(n_440),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_516),
.B(n_440),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_464),
.B(n_436),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_495),
.A2(n_439),
.B1(n_447),
.B2(n_444),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_506),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_476),
.B(n_440),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_502),
.B(n_440),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_471),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_499),
.B(n_405),
.Y(n_577)
);

NOR2x1p5_ASAP7_75t_L g578 ( 
.A(n_498),
.B(n_425),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_506),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_507),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_471),
.B(n_424),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_511),
.B(n_429),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_511),
.B(n_405),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_511),
.B(n_429),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_511),
.B(n_434),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_507),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_513),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_499),
.B(n_407),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_494),
.B(n_453),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_492),
.B(n_402),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_492),
.B(n_402),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_453),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_453),
.B(n_402),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_450),
.B(n_372),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_494),
.B(n_404),
.Y(n_595)
);

NAND3xp33_ASAP7_75t_L g596 ( 
.A(n_470),
.B(n_364),
.C(n_363),
.Y(n_596)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_450),
.B(n_373),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_450),
.B(n_363),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_450),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_454),
.B(n_402),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_510),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_483),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_454),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_483),
.B(n_364),
.Y(n_604)
);

OR2x2_ASAP7_75t_L g605 ( 
.A(n_483),
.B(n_365),
.Y(n_605)
);

O2A1O1Ixp5_ASAP7_75t_L g606 ( 
.A1(n_454),
.A2(n_415),
.B(n_404),
.C(n_413),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_465),
.B(n_404),
.Y(n_607)
);

BUFx6f_ASAP7_75t_SL g608 ( 
.A(n_483),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_465),
.B(n_404),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_465),
.B(n_413),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_470),
.Y(n_611)
);

OAI221xp5_ASAP7_75t_L g612 ( 
.A1(n_497),
.A2(n_403),
.B1(n_407),
.B2(n_433),
.C(n_408),
.Y(n_612)
);

NAND3xp33_ASAP7_75t_L g613 ( 
.A(n_486),
.B(n_369),
.C(n_365),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_497),
.B(n_413),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_497),
.B(n_413),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_486),
.B(n_382),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_487),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_487),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_520),
.B(n_408),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_528),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_542),
.B(n_408),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_537),
.B(n_392),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_583),
.B(n_392),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_540),
.A2(n_493),
.B(n_490),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_533),
.A2(n_493),
.B(n_490),
.Y(n_625)
);

OR2x2_ASAP7_75t_L g626 ( 
.A(n_535),
.B(n_415),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_550),
.A2(n_504),
.B(n_496),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_523),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_601),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_528),
.Y(n_630)
);

NOR2x2_ASAP7_75t_L g631 ( 
.A(n_554),
.B(n_392),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_541),
.A2(n_555),
.B(n_551),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_521),
.Y(n_633)
);

A2O1A1Ixp33_ASAP7_75t_L g634 ( 
.A1(n_542),
.A2(n_415),
.B(n_504),
.C(n_496),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_541),
.A2(n_488),
.B(n_477),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_583),
.B(n_396),
.Y(n_636)
);

AOI21xp33_ASAP7_75t_L g637 ( 
.A1(n_588),
.A2(n_396),
.B(n_303),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_L g638 ( 
.A(n_544),
.B(n_505),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_522),
.B(n_531),
.Y(n_639)
);

NAND2xp33_ASAP7_75t_L g640 ( 
.A(n_544),
.B(n_505),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_529),
.B(n_415),
.Y(n_641)
);

NOR2xp67_ASAP7_75t_L g642 ( 
.A(n_546),
.B(n_433),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_560),
.B(n_461),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_585),
.B(n_396),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_590),
.B(n_433),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_558),
.A2(n_488),
.B(n_477),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_559),
.A2(n_489),
.B(n_461),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_591),
.B(n_396),
.Y(n_648)
);

NOR2xp67_ASAP7_75t_L g649 ( 
.A(n_596),
.B(n_426),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_523),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_585),
.B(n_500),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_560),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_548),
.Y(n_653)
);

OAI21xp5_ASAP7_75t_L g654 ( 
.A1(n_606),
.A2(n_461),
.B(n_505),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_526),
.B(n_409),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_576),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_543),
.B(n_409),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_561),
.A2(n_489),
.B(n_461),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_565),
.A2(n_461),
.B(n_509),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_547),
.B(n_412),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_566),
.A2(n_461),
.B(n_509),
.Y(n_661)
);

A2O1A1Ixp33_ASAP7_75t_L g662 ( 
.A1(n_588),
.A2(n_403),
.B(n_416),
.C(n_417),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_607),
.A2(n_614),
.B(n_610),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_589),
.A2(n_595),
.B(n_532),
.Y(n_664)
);

INVx11_ASAP7_75t_L g665 ( 
.A(n_578),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_581),
.B(n_302),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_530),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_571),
.B(n_500),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_589),
.A2(n_472),
.B(n_468),
.Y(n_669)
);

AOI21x1_ASAP7_75t_L g670 ( 
.A1(n_570),
.A2(n_385),
.B(n_390),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_523),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_582),
.B(n_500),
.Y(n_672)
);

AO21x1_ASAP7_75t_L g673 ( 
.A1(n_524),
.A2(n_393),
.B(n_390),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_595),
.A2(n_472),
.B(n_468),
.Y(n_674)
);

AO21x2_ASAP7_75t_L g675 ( 
.A1(n_524),
.A2(n_393),
.B(n_385),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_532),
.A2(n_472),
.B(n_468),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_557),
.B(n_412),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_530),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_609),
.A2(n_615),
.B(n_569),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_L g680 ( 
.A(n_562),
.B(n_567),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_609),
.A2(n_472),
.B(n_468),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_615),
.A2(n_472),
.B(n_468),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_L g683 ( 
.A(n_562),
.B(n_567),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_611),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_545),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_577),
.A2(n_584),
.B1(n_604),
.B2(n_598),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_536),
.B(n_421),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_569),
.A2(n_508),
.B(n_475),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_563),
.B(n_416),
.Y(n_689)
);

OAI21xp5_ASAP7_75t_L g690 ( 
.A1(n_534),
.A2(n_505),
.B(n_439),
.Y(n_690)
);

BUFx8_ASAP7_75t_L g691 ( 
.A(n_608),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_536),
.B(n_421),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_570),
.A2(n_508),
.B(n_475),
.Y(n_693)
);

AO21x1_ASAP7_75t_L g694 ( 
.A1(n_577),
.A2(n_419),
.B(n_417),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_574),
.A2(n_508),
.B(n_475),
.Y(n_695)
);

AO21x1_ASAP7_75t_L g696 ( 
.A1(n_575),
.A2(n_420),
.B(n_419),
.Y(n_696)
);

OAI21xp33_ASAP7_75t_L g697 ( 
.A1(n_564),
.A2(n_218),
.B(n_188),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_593),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_616),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_597),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_594),
.B(n_308),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_521),
.Y(n_702)
);

O2A1O1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_600),
.A2(n_426),
.B(n_420),
.C(n_422),
.Y(n_703)
);

O2A1O1Ixp33_ASAP7_75t_L g704 ( 
.A1(n_592),
.A2(n_401),
.B(n_406),
.C(n_410),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_611),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_525),
.B(n_401),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_527),
.B(n_401),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_617),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_568),
.A2(n_508),
.B(n_475),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_527),
.B(n_406),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_536),
.B(n_475),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_538),
.B(n_572),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_539),
.Y(n_713)
);

AOI33xp33_ASAP7_75t_L g714 ( 
.A1(n_538),
.A2(n_427),
.A3(n_406),
.B1(n_410),
.B2(n_414),
.B3(n_422),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_605),
.B(n_421),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_603),
.A2(n_508),
.B(n_414),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_572),
.B(n_410),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_652),
.Y(n_718)
);

A2O1A1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_622),
.A2(n_636),
.B(n_623),
.C(n_715),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_666),
.B(n_599),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_644),
.B(n_321),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_656),
.B(n_552),
.Y(n_722)
);

OR2x6_ASAP7_75t_L g723 ( 
.A(n_629),
.B(n_602),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_632),
.A2(n_612),
.B(n_587),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_620),
.Y(n_725)
);

INVx5_ASAP7_75t_L g726 ( 
.A(n_628),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_623),
.B(n_636),
.Y(n_727)
);

OR2x6_ASAP7_75t_L g728 ( 
.A(n_700),
.B(n_587),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_619),
.A2(n_613),
.B1(n_539),
.B2(n_521),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_680),
.A2(n_580),
.B(n_573),
.Y(n_730)
);

INVx6_ASAP7_75t_L g731 ( 
.A(n_691),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_644),
.B(n_549),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_656),
.B(n_521),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_622),
.B(n_553),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_653),
.B(n_338),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_630),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_667),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_678),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_655),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_657),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_685),
.B(n_414),
.Y(n_741)
);

O2A1O1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_653),
.A2(n_422),
.B(n_427),
.C(n_586),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_701),
.B(n_340),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_633),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_699),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_660),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_686),
.B(n_351),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_SL g748 ( 
.A(n_691),
.B(n_355),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_713),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_637),
.A2(n_359),
.B1(n_360),
.B2(n_356),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_677),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_642),
.B(n_427),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_648),
.A2(n_367),
.B1(n_608),
.B2(n_698),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_651),
.B(n_553),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_713),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_651),
.B(n_553),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_683),
.A2(n_580),
.B(n_573),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_689),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_633),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_665),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_663),
.A2(n_617),
.B(n_579),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_628),
.B(n_553),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_626),
.B(n_618),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_715),
.B(n_421),
.Y(n_764)
);

INVx4_ASAP7_75t_L g765 ( 
.A(n_650),
.Y(n_765)
);

CKINVDCx16_ASAP7_75t_R g766 ( 
.A(n_631),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_704),
.Y(n_767)
);

NOR2x1_ASAP7_75t_SL g768 ( 
.A(n_633),
.B(n_702),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_633),
.Y(n_769)
);

O2A1O1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_662),
.A2(n_395),
.B(n_223),
.C(n_228),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_639),
.A2(n_439),
.B1(n_231),
.B2(n_234),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_702),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_639),
.A2(n_556),
.B(n_505),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_621),
.A2(n_439),
.B1(n_269),
.B2(n_229),
.Y(n_774)
);

BUFx8_ASAP7_75t_L g775 ( 
.A(n_702),
.Y(n_775)
);

A2O1A1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_668),
.A2(n_421),
.B(n_395),
.C(n_556),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_684),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_705),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_702),
.B(n_556),
.Y(n_779)
);

OAI21xp33_ASAP7_75t_L g780 ( 
.A1(n_697),
.A2(n_283),
.B(n_221),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_664),
.A2(n_635),
.B(n_674),
.Y(n_781)
);

O2A1O1Ixp5_ASAP7_75t_L g782 ( 
.A1(n_696),
.A2(n_505),
.B(n_556),
.C(n_439),
.Y(n_782)
);

INVx4_ASAP7_75t_L g783 ( 
.A(n_650),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_R g784 ( 
.A(n_671),
.B(n_505),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_708),
.Y(n_785)
);

OA22x2_ASAP7_75t_L g786 ( 
.A1(n_641),
.A2(n_232),
.B1(n_172),
.B2(n_189),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_671),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_760),
.Y(n_788)
);

AO31x2_ASAP7_75t_L g789 ( 
.A1(n_781),
.A2(n_694),
.A3(n_673),
.B(n_712),
.Y(n_789)
);

OAI21x1_ASAP7_75t_L g790 ( 
.A1(n_761),
.A2(n_676),
.B(n_625),
.Y(n_790)
);

A2O1A1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_727),
.A2(n_649),
.B(n_703),
.C(n_668),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_718),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_719),
.A2(n_640),
.B(n_638),
.Y(n_793)
);

OAI21x1_ASAP7_75t_L g794 ( 
.A1(n_773),
.A2(n_624),
.B(n_627),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_739),
.A2(n_645),
.B1(n_634),
.B2(n_706),
.Y(n_795)
);

CKINVDCx20_ASAP7_75t_R g796 ( 
.A(n_731),
.Y(n_796)
);

OAI21x1_ASAP7_75t_L g797 ( 
.A1(n_782),
.A2(n_688),
.B(n_695),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_721),
.B(n_421),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_724),
.A2(n_654),
.B(n_679),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_732),
.A2(n_709),
.B(n_669),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_764),
.A2(n_661),
.B(n_659),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_743),
.B(n_747),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_735),
.B(n_749),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_776),
.A2(n_693),
.B(n_643),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_725),
.Y(n_805)
);

OAI21x1_ASAP7_75t_L g806 ( 
.A1(n_730),
.A2(n_670),
.B(n_716),
.Y(n_806)
);

AOI221xp5_ASAP7_75t_L g807 ( 
.A1(n_753),
.A2(n_672),
.B1(n_397),
.B2(n_391),
.C(n_394),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_757),
.A2(n_643),
.B(n_647),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_740),
.A2(n_672),
.B1(n_717),
.B2(n_710),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_755),
.B(n_720),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_736),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_745),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_737),
.Y(n_813)
);

OAI22xp33_ASAP7_75t_L g814 ( 
.A1(n_748),
.A2(n_690),
.B1(n_707),
.B2(n_711),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_746),
.B(n_714),
.Y(n_815)
);

A2O1A1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_770),
.A2(n_646),
.B(n_711),
.C(n_658),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_751),
.A2(n_682),
.B(n_681),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_767),
.A2(n_692),
.B(n_687),
.Y(n_818)
);

OAI21x1_ASAP7_75t_L g819 ( 
.A1(n_734),
.A2(n_675),
.B(n_397),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_777),
.Y(n_820)
);

NOR4xp25_ASAP7_75t_L g821 ( 
.A(n_742),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_821)
);

OAI21x1_ASAP7_75t_L g822 ( 
.A1(n_754),
.A2(n_675),
.B(n_397),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_758),
.A2(n_756),
.B(n_729),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_763),
.A2(n_779),
.B(n_765),
.Y(n_824)
);

CKINVDCx11_ASAP7_75t_R g825 ( 
.A(n_723),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_765),
.A2(n_394),
.B(n_391),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_738),
.B(n_391),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_766),
.B(n_391),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_783),
.A2(n_394),
.B(n_397),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_783),
.A2(n_394),
.B(n_397),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_778),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_750),
.B(n_394),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_752),
.A2(n_394),
.B(n_397),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_741),
.B(n_723),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_744),
.Y(n_835)
);

O2A1O1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_780),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_836)
);

OAI21x1_ASAP7_75t_L g837 ( 
.A1(n_733),
.A2(n_398),
.B(n_439),
.Y(n_837)
);

AO31x2_ASAP7_75t_L g838 ( 
.A1(n_785),
.A2(n_418),
.A3(n_217),
.B(n_198),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_771),
.A2(n_222),
.B(n_286),
.C(n_265),
.Y(n_839)
);

AO31x2_ASAP7_75t_L g840 ( 
.A1(n_768),
.A2(n_418),
.A3(n_217),
.B(n_198),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_L g841 ( 
.A1(n_771),
.A2(n_418),
.B(n_263),
.Y(n_841)
);

AO31x2_ASAP7_75t_L g842 ( 
.A1(n_774),
.A2(n_418),
.A3(n_217),
.B(n_198),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_772),
.Y(n_843)
);

OAI21x1_ASAP7_75t_L g844 ( 
.A1(n_722),
.A2(n_418),
.B(n_112),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_726),
.A2(n_762),
.B(n_774),
.Y(n_845)
);

OAI21xp33_ASAP7_75t_SL g846 ( 
.A1(n_786),
.A2(n_12),
.B(n_14),
.Y(n_846)
);

AOI221x1_ASAP7_75t_L g847 ( 
.A1(n_762),
.A2(n_217),
.B1(n_418),
.B2(n_18),
.C(n_20),
.Y(n_847)
);

OAI21xp5_ASAP7_75t_SL g848 ( 
.A1(n_836),
.A2(n_787),
.B(n_731),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_802),
.A2(n_418),
.B1(n_728),
.B2(n_775),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_832),
.A2(n_418),
.B1(n_728),
.B2(n_775),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_803),
.B(n_744),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_807),
.A2(n_787),
.B1(n_784),
.B2(n_769),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_831),
.A2(n_787),
.B1(n_769),
.B2(n_759),
.Y(n_853)
);

CKINVDCx11_ASAP7_75t_R g854 ( 
.A(n_788),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_789),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_792),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_810),
.B(n_744),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_SL g858 ( 
.A1(n_846),
.A2(n_726),
.B1(n_759),
.B2(n_769),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_789),
.Y(n_859)
);

BUFx12f_ASAP7_75t_L g860 ( 
.A(n_825),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_839),
.A2(n_726),
.B1(n_759),
.B2(n_260),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_798),
.A2(n_255),
.B1(n_253),
.B2(n_252),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_805),
.Y(n_863)
);

CKINVDCx20_ASAP7_75t_R g864 ( 
.A(n_796),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_821),
.B(n_16),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_841),
.A2(n_217),
.B1(n_246),
.B2(n_245),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_843),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_811),
.Y(n_868)
);

NAND2x1p5_ASAP7_75t_L g869 ( 
.A(n_834),
.B(n_49),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_812),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_813),
.Y(n_871)
);

CKINVDCx20_ASAP7_75t_R g872 ( 
.A(n_828),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_820),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_835),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_835),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_835),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_815),
.B(n_16),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_827),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_841),
.A2(n_249),
.B1(n_243),
.B2(n_235),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_814),
.A2(n_226),
.B1(n_224),
.B2(n_215),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_827),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_SL g882 ( 
.A1(n_793),
.A2(n_795),
.B1(n_809),
.B2(n_845),
.Y(n_882)
);

CKINVDCx11_ASAP7_75t_R g883 ( 
.A(n_795),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_818),
.Y(n_884)
);

BUFx10_ASAP7_75t_L g885 ( 
.A(n_847),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_809),
.A2(n_212),
.B1(n_211),
.B2(n_209),
.Y(n_886)
);

BUFx4f_ASAP7_75t_SL g887 ( 
.A(n_824),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_SL g888 ( 
.A1(n_821),
.A2(n_823),
.B1(n_844),
.B2(n_818),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_789),
.Y(n_889)
);

OAI22xp33_ASAP7_75t_L g890 ( 
.A1(n_799),
.A2(n_207),
.B1(n_206),
.B2(n_203),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_SL g891 ( 
.A1(n_842),
.A2(n_195),
.B1(n_193),
.B2(n_192),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_837),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_819),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_838),
.Y(n_894)
);

INVx2_ASAP7_75t_R g895 ( 
.A(n_842),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_822),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_794),
.Y(n_897)
);

INVx6_ASAP7_75t_L g898 ( 
.A(n_791),
.Y(n_898)
);

INVx4_ASAP7_75t_L g899 ( 
.A(n_826),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_829),
.Y(n_900)
);

INVx3_ASAP7_75t_L g901 ( 
.A(n_797),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_838),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_842),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_SL g904 ( 
.A1(n_804),
.A2(n_190),
.B1(n_171),
.B2(n_21),
.Y(n_904)
);

INVx4_ASAP7_75t_L g905 ( 
.A(n_830),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_816),
.A2(n_17),
.B1(n_18),
.B2(n_21),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_SL g907 ( 
.A1(n_833),
.A2(n_17),
.B1(n_22),
.B2(n_23),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_838),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_855),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_855),
.B(n_840),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_883),
.A2(n_865),
.B1(n_898),
.B2(n_906),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_859),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_898),
.B(n_22),
.Y(n_913)
);

AO21x2_ASAP7_75t_L g914 ( 
.A1(n_894),
.A2(n_801),
.B(n_800),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_859),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_889),
.B(n_817),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_898),
.A2(n_808),
.B1(n_24),
.B2(n_25),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_889),
.Y(n_918)
);

BUFx2_ASAP7_75t_SL g919 ( 
.A(n_905),
.Y(n_919)
);

BUFx12f_ASAP7_75t_L g920 ( 
.A(n_854),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_901),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_884),
.B(n_840),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_878),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_881),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_901),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_901),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_902),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_893),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_893),
.Y(n_929)
);

OAI21x1_ASAP7_75t_L g930 ( 
.A1(n_897),
.A2(n_790),
.B(n_806),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_896),
.Y(n_931)
);

INVxp67_ASAP7_75t_SL g932 ( 
.A(n_896),
.Y(n_932)
);

INVx6_ASAP7_75t_L g933 ( 
.A(n_898),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_897),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_908),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_905),
.Y(n_936)
);

OA21x2_ASAP7_75t_L g937 ( 
.A1(n_903),
.A2(n_840),
.B(n_24),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_903),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_882),
.B(n_23),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_863),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_892),
.Y(n_941)
);

OA21x2_ASAP7_75t_L g942 ( 
.A1(n_868),
.A2(n_25),
.B(n_26),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_883),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_892),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_892),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_856),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_871),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_873),
.Y(n_948)
);

O2A1O1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_917),
.A2(n_865),
.B(n_877),
.C(n_848),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_917),
.A2(n_888),
.B(n_900),
.Y(n_950)
);

AO32x2_ASAP7_75t_L g951 ( 
.A1(n_946),
.A2(n_905),
.A3(n_899),
.B1(n_895),
.B2(n_861),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_948),
.B(n_876),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_946),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_948),
.B(n_876),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_911),
.A2(n_880),
.B1(n_886),
.B2(n_904),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_948),
.Y(n_956)
);

INVx5_ASAP7_75t_L g957 ( 
.A(n_933),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_913),
.A2(n_870),
.B(n_890),
.C(n_857),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_948),
.Y(n_959)
);

AO21x1_ASAP7_75t_SL g960 ( 
.A1(n_911),
.A2(n_851),
.B(n_887),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_925),
.Y(n_961)
);

OR2x2_ASAP7_75t_L g962 ( 
.A(n_947),
.B(n_895),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_911),
.A2(n_872),
.B1(n_867),
.B2(n_850),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_940),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_940),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_940),
.B(n_900),
.Y(n_966)
);

INVxp67_ASAP7_75t_L g967 ( 
.A(n_913),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_938),
.B(n_875),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_947),
.B(n_885),
.Y(n_969)
);

AO21x2_ASAP7_75t_L g970 ( 
.A1(n_922),
.A2(n_862),
.B(n_885),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_947),
.B(n_885),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_920),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_923),
.B(n_872),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_939),
.A2(n_866),
.B(n_879),
.C(n_858),
.Y(n_974)
);

OA21x2_ASAP7_75t_L g975 ( 
.A1(n_930),
.A2(n_853),
.B(n_852),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_923),
.B(n_874),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_939),
.A2(n_891),
.B(n_907),
.C(n_849),
.Y(n_977)
);

OA21x2_ASAP7_75t_L g978 ( 
.A1(n_930),
.A2(n_899),
.B(n_869),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_923),
.B(n_899),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_938),
.B(n_875),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_924),
.B(n_875),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_939),
.A2(n_943),
.B(n_938),
.C(n_922),
.Y(n_982)
);

AO32x2_ASAP7_75t_L g983 ( 
.A1(n_938),
.A2(n_867),
.A3(n_869),
.B1(n_875),
.B2(n_874),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_924),
.B(n_875),
.Y(n_984)
);

OA21x2_ASAP7_75t_L g985 ( 
.A1(n_930),
.A2(n_874),
.B(n_28),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_924),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_936),
.B(n_27),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_927),
.B(n_27),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_936),
.B(n_28),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_936),
.B(n_29),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_956),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_961),
.B(n_925),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_953),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_959),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_966),
.B(n_921),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_966),
.B(n_921),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_963),
.A2(n_943),
.B1(n_933),
.B2(n_942),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_956),
.B(n_927),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_972),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_979),
.B(n_921),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_979),
.B(n_921),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_981),
.B(n_941),
.Y(n_1002)
);

NAND2x1p5_ASAP7_75t_L g1003 ( 
.A(n_957),
.B(n_943),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_962),
.Y(n_1004)
);

INVxp67_ASAP7_75t_L g1005 ( 
.A(n_970),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_964),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_965),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_972),
.B(n_920),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_962),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_986),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_976),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_970),
.B(n_982),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_961),
.B(n_925),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_981),
.B(n_941),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_984),
.B(n_941),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_985),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_984),
.B(n_961),
.Y(n_1017)
);

AO22x1_ASAP7_75t_L g1018 ( 
.A1(n_1012),
.A2(n_943),
.B1(n_957),
.B2(n_967),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_1017),
.B(n_982),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_1017),
.B(n_983),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_1003),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_997),
.A2(n_950),
.B1(n_949),
.B2(n_974),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_1003),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_1011),
.B(n_969),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_992),
.Y(n_1025)
);

NOR2xp67_ASAP7_75t_L g1026 ( 
.A(n_991),
.B(n_920),
.Y(n_1026)
);

INVx2_ASAP7_75t_SL g1027 ( 
.A(n_1017),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_994),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_995),
.B(n_983),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_994),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_992),
.B(n_952),
.Y(n_1031)
);

INVx4_ASAP7_75t_L g1032 ( 
.A(n_999),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_993),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_998),
.Y(n_1034)
);

OAI33xp33_ASAP7_75t_L g1035 ( 
.A1(n_1012),
.A2(n_955),
.A3(n_973),
.B1(n_988),
.B2(n_958),
.B3(n_927),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_1011),
.B(n_969),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_998),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1006),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_1019),
.B(n_1003),
.Y(n_1039)
);

BUFx12f_ASAP7_75t_L g1040 ( 
.A(n_1032),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_1019),
.B(n_1003),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1020),
.B(n_995),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_1020),
.B(n_1029),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1038),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_1025),
.B(n_1016),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_1022),
.A2(n_997),
.B1(n_970),
.B2(n_933),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_1034),
.B(n_1006),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_1029),
.B(n_995),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_1034),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_1031),
.B(n_996),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_1040),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_1039),
.B(n_1031),
.Y(n_1052)
);

NAND2x1p5_ASAP7_75t_L g1053 ( 
.A(n_1039),
.B(n_987),
.Y(n_1053)
);

NAND2x1p5_ASAP7_75t_L g1054 ( 
.A(n_1041),
.B(n_987),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_1041),
.B(n_1031),
.Y(n_1055)
);

INVx2_ASAP7_75t_SL g1056 ( 
.A(n_1040),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1044),
.Y(n_1057)
);

OR2x2_ASAP7_75t_L g1058 ( 
.A(n_1043),
.B(n_1033),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1053),
.B(n_1049),
.Y(n_1059)
);

INVxp67_ASAP7_75t_L g1060 ( 
.A(n_1051),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_1055),
.B(n_1043),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1053),
.B(n_1049),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_1055),
.B(n_1050),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1061),
.B(n_1051),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1060),
.Y(n_1065)
);

NAND2xp33_ASAP7_75t_SL g1066 ( 
.A(n_1059),
.B(n_1056),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1060),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_1063),
.A2(n_1046),
.B1(n_1054),
.B2(n_1058),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_1062),
.A2(n_1046),
.B1(n_1054),
.B2(n_1052),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1061),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1061),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1061),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1061),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1061),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_SL g1075 ( 
.A1(n_1065),
.A2(n_1056),
.B(n_860),
.Y(n_1075)
);

AOI221xp5_ASAP7_75t_L g1076 ( 
.A1(n_1068),
.A2(n_1035),
.B1(n_1018),
.B2(n_1005),
.C(n_1057),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1074),
.B(n_1042),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1067),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_1074),
.B(n_1040),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1070),
.Y(n_1080)
);

OAI221xp5_ASAP7_75t_L g1081 ( 
.A1(n_1069),
.A2(n_974),
.B1(n_977),
.B2(n_1005),
.C(n_1016),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_1064),
.B(n_1032),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1071),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1066),
.A2(n_1018),
.B(n_1032),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1072),
.Y(n_1085)
);

INVxp67_ASAP7_75t_L g1086 ( 
.A(n_1066),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1073),
.Y(n_1087)
);

OAI322xp33_ASAP7_75t_L g1088 ( 
.A1(n_1065),
.A2(n_988),
.A3(n_1016),
.B1(n_1044),
.B2(n_1047),
.C1(n_1037),
.C2(n_1008),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_1066),
.B(n_920),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1065),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1078),
.Y(n_1091)
);

AOI222xp33_ASAP7_75t_L g1092 ( 
.A1(n_1076),
.A2(n_977),
.B1(n_860),
.B2(n_1045),
.C1(n_1048),
.C2(n_990),
.Y(n_1092)
);

OAI221xp5_ASAP7_75t_L g1093 ( 
.A1(n_1081),
.A2(n_1026),
.B1(n_942),
.B2(n_985),
.C(n_1047),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1090),
.B(n_1042),
.Y(n_1094)
);

INVx1_ASAP7_75t_SL g1095 ( 
.A(n_1082),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1079),
.B(n_1086),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1080),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1086),
.Y(n_1098)
);

NAND2xp33_ASAP7_75t_L g1099 ( 
.A(n_1084),
.B(n_864),
.Y(n_1099)
);

NAND3xp33_ASAP7_75t_L g1100 ( 
.A(n_1083),
.B(n_990),
.C(n_989),
.Y(n_1100)
);

INVxp67_ASAP7_75t_L g1101 ( 
.A(n_1085),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_1087),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1077),
.Y(n_1103)
);

OAI221xp5_ASAP7_75t_L g1104 ( 
.A1(n_1089),
.A2(n_942),
.B1(n_985),
.B2(n_1023),
.C(n_1021),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1089),
.B(n_1048),
.Y(n_1105)
);

OR2x2_ASAP7_75t_L g1106 ( 
.A(n_1075),
.B(n_1037),
.Y(n_1106)
);

OAI222xp33_ASAP7_75t_L g1107 ( 
.A1(n_1088),
.A2(n_1045),
.B1(n_1023),
.B2(n_1021),
.C1(n_864),
.C2(n_989),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1086),
.A2(n_1045),
.B(n_942),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1078),
.Y(n_1109)
);

NOR3x1_ASAP7_75t_L g1110 ( 
.A(n_1103),
.B(n_854),
.C(n_1027),
.Y(n_1110)
);

NAND4xp25_ASAP7_75t_L g1111 ( 
.A(n_1095),
.B(n_1025),
.C(n_1050),
.D(n_1045),
.Y(n_1111)
);

NOR3xp33_ASAP7_75t_L g1112 ( 
.A(n_1098),
.B(n_1036),
.C(n_1024),
.Y(n_1112)
);

NOR3xp33_ASAP7_75t_L g1113 ( 
.A(n_1098),
.B(n_1030),
.C(n_1028),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1102),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_1096),
.B(n_1025),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_1100),
.B(n_1038),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1094),
.B(n_1027),
.Y(n_1117)
);

AOI221xp5_ASAP7_75t_L g1118 ( 
.A1(n_1093),
.A2(n_1030),
.B1(n_1028),
.B2(n_971),
.C(n_1007),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1099),
.A2(n_942),
.B(n_991),
.Y(n_1119)
);

NOR2x1_ASAP7_75t_L g1120 ( 
.A(n_1091),
.B(n_942),
.Y(n_1120)
);

NOR2xp67_ASAP7_75t_L g1121 ( 
.A(n_1102),
.B(n_1101),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1097),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1101),
.B(n_991),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1109),
.B(n_1007),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_1106),
.B(n_1105),
.Y(n_1125)
);

NAND3xp33_ASAP7_75t_L g1126 ( 
.A(n_1092),
.B(n_1108),
.C(n_1104),
.Y(n_1126)
);

INVxp67_ASAP7_75t_L g1127 ( 
.A(n_1121),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1114),
.A2(n_1107),
.B(n_942),
.Y(n_1128)
);

AOI222xp33_ASAP7_75t_L g1129 ( 
.A1(n_1126),
.A2(n_971),
.B1(n_1004),
.B2(n_1009),
.C1(n_933),
.C2(n_983),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1124),
.Y(n_1130)
);

XNOR2xp5_ASAP7_75t_L g1131 ( 
.A(n_1115),
.B(n_29),
.Y(n_1131)
);

OAI21xp33_ASAP7_75t_L g1132 ( 
.A1(n_1125),
.A2(n_996),
.B(n_1014),
.Y(n_1132)
);

AOI211xp5_ASAP7_75t_L g1133 ( 
.A1(n_1122),
.A2(n_996),
.B(n_1010),
.C(n_1001),
.Y(n_1133)
);

OAI31xp33_ASAP7_75t_L g1134 ( 
.A1(n_1119),
.A2(n_983),
.A3(n_1009),
.B(n_1004),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1110),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_1120),
.A2(n_1010),
.B(n_1004),
.C(n_1009),
.Y(n_1136)
);

AOI222xp33_ASAP7_75t_L g1137 ( 
.A1(n_1118),
.A2(n_933),
.B1(n_935),
.B2(n_951),
.C1(n_952),
.C2(n_954),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1117),
.Y(n_1138)
);

NOR2x1_ASAP7_75t_L g1139 ( 
.A(n_1111),
.B(n_30),
.Y(n_1139)
);

NAND3xp33_ASAP7_75t_SL g1140 ( 
.A(n_1112),
.B(n_30),
.C(n_31),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_1123),
.A2(n_937),
.B(n_34),
.C(n_35),
.Y(n_1141)
);

OAI211xp5_ASAP7_75t_L g1142 ( 
.A1(n_1116),
.A2(n_1113),
.B(n_37),
.C(n_38),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1120),
.A2(n_960),
.B1(n_933),
.B2(n_957),
.Y(n_1143)
);

AOI221xp5_ASAP7_75t_L g1144 ( 
.A1(n_1126),
.A2(n_1015),
.B1(n_1014),
.B2(n_1002),
.C(n_952),
.Y(n_1144)
);

AOI221xp5_ASAP7_75t_SL g1145 ( 
.A1(n_1114),
.A2(n_1001),
.B1(n_1000),
.B2(n_1002),
.C(n_1015),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_1114),
.Y(n_1146)
);

NAND4xp25_ASAP7_75t_L g1147 ( 
.A(n_1121),
.B(n_32),
.C(n_37),
.D(n_40),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_1126),
.A2(n_954),
.B(n_1014),
.C(n_1015),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1121),
.A2(n_1013),
.B(n_992),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1121),
.A2(n_933),
.B1(n_1002),
.B2(n_1001),
.Y(n_1150)
);

NAND4xp25_ASAP7_75t_L g1151 ( 
.A(n_1135),
.B(n_1013),
.C(n_992),
.D(n_1000),
.Y(n_1151)
);

AO22x2_ASAP7_75t_L g1152 ( 
.A1(n_1127),
.A2(n_1138),
.B1(n_1130),
.B2(n_1142),
.Y(n_1152)
);

AOI32xp33_ASAP7_75t_L g1153 ( 
.A1(n_1139),
.A2(n_1000),
.A3(n_954),
.B1(n_980),
.B2(n_968),
.Y(n_1153)
);

OAI222xp33_ASAP7_75t_L g1154 ( 
.A1(n_1146),
.A2(n_957),
.B1(n_951),
.B2(n_935),
.C1(n_968),
.C2(n_980),
.Y(n_1154)
);

NOR3xp33_ASAP7_75t_L g1155 ( 
.A(n_1147),
.B(n_1140),
.C(n_1141),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_SL g1156 ( 
.A1(n_1128),
.A2(n_32),
.B(n_41),
.C(n_42),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1131),
.A2(n_1148),
.B1(n_1133),
.B2(n_1150),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1147),
.A2(n_968),
.B(n_980),
.C(n_47),
.Y(n_1158)
);

AO221x1_ASAP7_75t_L g1159 ( 
.A1(n_1149),
.A2(n_925),
.B1(n_926),
.B2(n_47),
.C(n_41),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1129),
.A2(n_937),
.B1(n_978),
.B2(n_957),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_1136),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1132),
.Y(n_1162)
);

A2O1A1Ixp33_ASAP7_75t_SL g1163 ( 
.A1(n_1134),
.A2(n_44),
.B(n_925),
.C(n_926),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1145),
.B(n_44),
.Y(n_1164)
);

NOR4xp25_ASAP7_75t_SL g1165 ( 
.A(n_1144),
.B(n_951),
.C(n_935),
.D(n_919),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1143),
.Y(n_1166)
);

OAI211xp5_ASAP7_75t_L g1167 ( 
.A1(n_1137),
.A2(n_926),
.B(n_925),
.C(n_937),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1139),
.A2(n_937),
.B1(n_978),
.B2(n_975),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1147),
.B(n_978),
.Y(n_1169)
);

AOI31xp33_ASAP7_75t_L g1170 ( 
.A1(n_1127),
.A2(n_1013),
.A3(n_992),
.B(n_944),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_R g1171 ( 
.A(n_1146),
.B(n_51),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1127),
.A2(n_1013),
.B1(n_919),
.B2(n_926),
.Y(n_1172)
);

AOI221xp5_ASAP7_75t_L g1173 ( 
.A1(n_1127),
.A2(n_914),
.B1(n_951),
.B2(n_944),
.C(n_945),
.Y(n_1173)
);

AOI221xp5_ASAP7_75t_SL g1174 ( 
.A1(n_1127),
.A2(n_919),
.B1(n_926),
.B2(n_944),
.C(n_945),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1152),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1159),
.B(n_1013),
.Y(n_1176)
);

NOR3xp33_ASAP7_75t_L g1177 ( 
.A(n_1164),
.B(n_932),
.C(n_916),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1152),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1161),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1166),
.Y(n_1180)
);

OR2x2_ASAP7_75t_L g1181 ( 
.A(n_1162),
.B(n_1156),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1155),
.A2(n_937),
.B1(n_975),
.B2(n_914),
.Y(n_1182)
);

NOR2x1_ASAP7_75t_L g1183 ( 
.A(n_1158),
.B(n_926),
.Y(n_1183)
);

XNOR2xp5_ASAP7_75t_L g1184 ( 
.A(n_1157),
.B(n_937),
.Y(n_1184)
);

XNOR2xp5_ASAP7_75t_L g1185 ( 
.A(n_1151),
.B(n_937),
.Y(n_1185)
);

INVxp33_ASAP7_75t_L g1186 ( 
.A(n_1171),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1169),
.Y(n_1187)
);

NOR2x1p5_ASAP7_75t_L g1188 ( 
.A(n_1163),
.B(n_941),
.Y(n_1188)
);

NAND2x1p5_ASAP7_75t_L g1189 ( 
.A(n_1168),
.B(n_975),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1160),
.B(n_944),
.Y(n_1190)
);

INVxp67_ASAP7_75t_L g1191 ( 
.A(n_1170),
.Y(n_1191)
);

NAND4xp75_ASAP7_75t_L g1192 ( 
.A(n_1174),
.B(n_910),
.C(n_951),
.D(n_945),
.Y(n_1192)
);

NOR2x1_ASAP7_75t_L g1193 ( 
.A(n_1167),
.B(n_914),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1172),
.Y(n_1194)
);

XOR2x2_ASAP7_75t_L g1195 ( 
.A(n_1153),
.B(n_52),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1173),
.Y(n_1196)
);

NAND3xp33_ASAP7_75t_SL g1197 ( 
.A(n_1175),
.B(n_1165),
.C(n_1154),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1175),
.A2(n_945),
.B(n_914),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1178),
.A2(n_1181),
.B(n_1191),
.Y(n_1199)
);

NAND3xp33_ASAP7_75t_L g1200 ( 
.A(n_1179),
.B(n_931),
.C(n_916),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1176),
.B(n_914),
.Y(n_1201)
);

AOI221xp5_ASAP7_75t_L g1202 ( 
.A1(n_1187),
.A2(n_914),
.B1(n_932),
.B2(n_931),
.C(n_934),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_1194),
.B(n_930),
.Y(n_1203)
);

NOR2x1p5_ASAP7_75t_L g1204 ( 
.A(n_1180),
.B(n_916),
.Y(n_1204)
);

NAND3xp33_ASAP7_75t_L g1205 ( 
.A(n_1186),
.B(n_934),
.C(n_910),
.Y(n_1205)
);

OAI322xp33_ASAP7_75t_L g1206 ( 
.A1(n_1196),
.A2(n_934),
.A3(n_929),
.B1(n_928),
.B2(n_918),
.C1(n_915),
.C2(n_912),
.Y(n_1206)
);

AOI31xp33_ASAP7_75t_L g1207 ( 
.A1(n_1183),
.A2(n_53),
.A3(n_55),
.B(n_56),
.Y(n_1207)
);

XNOR2xp5_ASAP7_75t_L g1208 ( 
.A(n_1195),
.B(n_57),
.Y(n_1208)
);

AOI21xp33_ASAP7_75t_L g1209 ( 
.A1(n_1184),
.A2(n_58),
.B(n_63),
.Y(n_1209)
);

O2A1O1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1177),
.A2(n_934),
.B(n_929),
.C(n_928),
.Y(n_1210)
);

NOR3xp33_ASAP7_75t_L g1211 ( 
.A(n_1193),
.B(n_65),
.C(n_69),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1199),
.A2(n_1188),
.B(n_1190),
.C(n_1182),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1208),
.Y(n_1213)
);

XOR2x1_ASAP7_75t_L g1214 ( 
.A(n_1203),
.B(n_1190),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1204),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1203),
.B(n_1185),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1201),
.B(n_1192),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1197),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1207),
.Y(n_1219)
);

OA22x2_ASAP7_75t_L g1220 ( 
.A1(n_1209),
.A2(n_1189),
.B1(n_929),
.B2(n_928),
.Y(n_1220)
);

XOR2xp5_ASAP7_75t_L g1221 ( 
.A(n_1200),
.B(n_1205),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1211),
.Y(n_1222)
);

NAND4xp75_ASAP7_75t_L g1223 ( 
.A(n_1198),
.B(n_73),
.C(n_74),
.D(n_75),
.Y(n_1223)
);

OAI22x1_ASAP7_75t_L g1224 ( 
.A1(n_1210),
.A2(n_929),
.B1(n_928),
.B2(n_910),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1206),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1202),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1218),
.Y(n_1227)
);

OAI22x1_ASAP7_75t_L g1228 ( 
.A1(n_1219),
.A2(n_909),
.B1(n_78),
.B2(n_79),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1215),
.Y(n_1229)
);

BUFx4f_ASAP7_75t_SL g1230 ( 
.A(n_1213),
.Y(n_1230)
);

AO22x2_ASAP7_75t_L g1231 ( 
.A1(n_1222),
.A2(n_76),
.B1(n_80),
.B2(n_87),
.Y(n_1231)
);

AO22x2_ASAP7_75t_L g1232 ( 
.A1(n_1225),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_1232)
);

AOI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1217),
.A2(n_918),
.B1(n_915),
.B2(n_912),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1216),
.A2(n_1221),
.B1(n_1226),
.B2(n_1212),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1220),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1223),
.A2(n_918),
.B1(n_915),
.B2(n_912),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1227),
.A2(n_1223),
.B1(n_1214),
.B2(n_1224),
.Y(n_1237)
);

HB1xp67_ASAP7_75t_L g1238 ( 
.A(n_1228),
.Y(n_1238)
);

INVx1_ASAP7_75t_SL g1239 ( 
.A(n_1230),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1229),
.B(n_92),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1235),
.A2(n_918),
.B1(n_915),
.B2(n_912),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1232),
.Y(n_1242)
);

AOI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1242),
.A2(n_1238),
.B1(n_1234),
.B2(n_1239),
.Y(n_1243)
);

XNOR2xp5_ASAP7_75t_L g1244 ( 
.A(n_1237),
.B(n_1231),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1240),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1241),
.A2(n_1233),
.B(n_1236),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1243),
.A2(n_93),
.B(n_97),
.Y(n_1247)
);

NAND3xp33_ASAP7_75t_L g1248 ( 
.A(n_1247),
.B(n_1244),
.C(n_1245),
.Y(n_1248)
);

AOI211xp5_ASAP7_75t_L g1249 ( 
.A1(n_1248),
.A2(n_1246),
.B(n_107),
.C(n_108),
.Y(n_1249)
);

XOR2xp5_ASAP7_75t_L g1250 ( 
.A(n_1249),
.B(n_98),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1250),
.A2(n_111),
.B1(n_117),
.B2(n_118),
.Y(n_1251)
);

AOI211xp5_ASAP7_75t_L g1252 ( 
.A1(n_1251),
.A2(n_119),
.B(n_121),
.C(n_127),
.Y(n_1252)
);


endmodule