module fake_jpeg_7350_n_81 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_81);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_81;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx2_ASAP7_75t_SL g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_9),
.B(n_25),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_28),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_30),
.B1(n_29),
.B2(n_5),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_2),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_42),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_44),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_3),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_3),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_46),
.Y(n_61)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_29),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_44),
.B(n_33),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_54),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_5),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_56),
.B1(n_60),
.B2(n_62),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_32),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_11),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_12),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_13),
.B1(n_14),
.B2(n_18),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_27),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_68),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_19),
.C(n_20),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_63),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_52),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_74),
.Y(n_75)
);

FAx1_ASAP7_75t_SL g74 ( 
.A(n_71),
.B(n_70),
.CI(n_67),
.CON(n_74),
.SN(n_74)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_74),
.C(n_66),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_67),
.C(n_74),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_50),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_69),
.C(n_51),
.Y(n_79)
);

AOI322xp5_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_64),
.A3(n_62),
.B1(n_56),
.B2(n_22),
.C1(n_23),
.C2(n_26),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_21),
.Y(n_81)
);


endmodule