module fake_jpeg_12450_n_141 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_141);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_0),
.B(n_5),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_15),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_19),
.B(n_1),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_4),
.Y(n_45)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_34),
.Y(n_54)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_3),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_17),
.A2(n_4),
.B(n_6),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_14),
.C(n_4),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_38),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_35),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_26),
.B1(n_17),
.B2(n_29),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_51),
.B1(n_37),
.B2(n_32),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_45),
.B(n_52),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_46),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_27),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_50),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_27),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_31),
.A2(n_26),
.B1(n_19),
.B2(n_24),
.Y(n_51)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_27),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_56),
.B(n_61),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_63),
.C(n_52),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_73),
.Y(n_83)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx24_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_30),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_28),
.B1(n_16),
.B2(n_24),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_21),
.B1(n_20),
.B2(n_28),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_18),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_18),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_20),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_79),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_77),
.B(n_21),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_57),
.A2(n_50),
.B(n_47),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_59),
.A2(n_54),
.B(n_50),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_85),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_47),
.B1(n_35),
.B2(n_34),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_84),
.A2(n_89),
.B1(n_35),
.B2(n_58),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_54),
.B(n_44),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_66),
.B1(n_63),
.B2(n_68),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_66),
.B1(n_70),
.B2(n_69),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_94),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_62),
.B1(n_71),
.B2(n_58),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_81),
.B(n_62),
.Y(n_98)
);

BUFx12f_ASAP7_75t_SL g99 ( 
.A(n_86),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_101),
.B1(n_102),
.B2(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_79),
.C(n_89),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_109),
.C(n_86),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_82),
.B(n_85),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_111),
.B(n_94),
.Y(n_117)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_83),
.C(n_80),
.Y(n_109)
);

A2O1A1O1Ixp25_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_76),
.B(n_81),
.C(n_84),
.D(n_77),
.Y(n_111)
);

AOI322xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_22),
.A3(n_16),
.B1(n_14),
.B2(n_86),
.C1(n_44),
.C2(n_11),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_99),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_117),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_109),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_119),
.C(n_108),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_91),
.B(n_86),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_105),
.Y(n_124)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_106),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_126),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

NOR2xp67_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_111),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_117),
.C(n_108),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_116),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_131),
.C(n_23),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_123),
.B(n_113),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_122),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_133),
.A2(n_134),
.B1(n_136),
.B2(n_6),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_115),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_128),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_13),
.Y(n_136)
);

NAND4xp25_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_7),
.C(n_10),
.D(n_11),
.Y(n_139)
);

NOR3xp33_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_13),
.C(n_137),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_140),
.Y(n_141)
);


endmodule