module fake_jpeg_1356_n_227 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_227);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_50),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx4f_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx16f_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_10),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_8),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_7),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_22),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_82),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_85),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_72),
.B(n_0),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_56),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_94),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_81),
.A2(n_64),
.B1(n_58),
.B2(n_54),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_74),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_59),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_87),
.A2(n_54),
.B1(n_65),
.B2(n_79),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_70),
.C(n_77),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_68),
.B1(n_76),
.B2(n_62),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_62),
.B1(n_70),
.B2(n_86),
.Y(n_113)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_94),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_105),
.B(n_110),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_107),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_78),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_100),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_114),
.Y(n_129)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_115),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_113),
.A2(n_59),
.B1(n_97),
.B2(n_68),
.Y(n_121)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_88),
.B(n_73),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_119),
.Y(n_137)
);

BUFx4f_ASAP7_75t_SL g117 ( 
.A(n_95),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_117),
.Y(n_133)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_99),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_61),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_96),
.C(n_90),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_139),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_109),
.A2(n_103),
.B1(n_113),
.B2(n_118),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_122),
.A2(n_131),
.B1(n_132),
.B2(n_138),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_109),
.A2(n_92),
.B(n_99),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_123),
.A2(n_53),
.B(n_52),
.Y(n_152)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_60),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_0),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_55),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_128),
.B(n_136),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_83),
.B1(n_69),
.B2(n_71),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_99),
.B1(n_68),
.B2(n_76),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_134),
.B(n_51),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_57),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_76),
.B1(n_77),
.B2(n_57),
.Y(n_138)
);

BUFx24_ASAP7_75t_SL g139 ( 
.A(n_117),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_126),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_147),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_125),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_150),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_130),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_71),
.B1(n_69),
.B2(n_75),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_151),
.A2(n_161),
.B1(n_35),
.B2(n_33),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_38),
.B(n_37),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_154),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_133),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_158),
.Y(n_175)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

NOR3xp33_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_1),
.C(n_2),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_123),
.A2(n_129),
.B1(n_120),
.B2(n_131),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_129),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_163),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_140),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_49),
.Y(n_164)
);

A2O1A1O1Ixp25_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_3),
.B(n_4),
.C(n_6),
.D(n_7),
.Y(n_169)
);

NAND2x1p5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_3),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_165),
.A2(n_4),
.B(n_8),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_165),
.B(n_46),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_152),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_174),
.B(n_153),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_43),
.C(n_42),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_173),
.C(n_176),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_41),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_40),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_146),
.Y(n_179)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_181),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_143),
.A2(n_148),
.B1(n_144),
.B2(n_142),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_184),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_165),
.C(n_156),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_16),
.C(n_17),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_186),
.B(n_189),
.Y(n_208)
);

FAx1_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_144),
.CI(n_151),
.CON(n_187),
.SN(n_187)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_187),
.A2(n_180),
.B(n_169),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_166),
.Y(n_202)
);

OAI322xp33_ASAP7_75t_L g189 ( 
.A1(n_182),
.A2(n_157),
.A3(n_32),
.B1(n_30),
.B2(n_29),
.C1(n_27),
.C2(n_25),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_190),
.A2(n_174),
.B1(n_181),
.B2(n_167),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_11),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_196),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_172),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_168),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_170),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_197),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_199),
.B(n_202),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_200),
.A2(n_204),
.B1(n_198),
.B2(n_175),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_201),
.A2(n_206),
.B1(n_207),
.B2(n_173),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_187),
.A2(n_183),
.B1(n_171),
.B2(n_178),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_205),
.A2(n_186),
.B(n_198),
.Y(n_212)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_200),
.Y(n_210)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_210),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_211),
.A2(n_214),
.B(n_215),
.Y(n_218)
);

NAND4xp25_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_208),
.C(n_203),
.D(n_20),
.Y(n_216)
);

XNOR2x1_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_203),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_207),
.A2(n_176),
.B(n_191),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_205),
.A2(n_191),
.B1(n_19),
.B2(n_20),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_217),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_209),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_215),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_220),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_214),
.C(n_219),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_224),
.A2(n_18),
.B(n_19),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_18),
.B(n_21),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_23),
.Y(n_227)
);


endmodule